TASK_RSTEN;
TASK_RST;
TASK_INIT_WRITE_SPI;
// write data into LB and array
TASK_LBWR(16'h0000);
TASK_LBWR(16'h0001);
TASK_LBWR(16'h0002);
TASK_LBWR(16'h0003);
TASK_LBWR(16'h0004);
TASK_LBWR(16'h0005);
TASK_LBWR(16'h0006);
TASK_LBWR(16'h0007);
TASK_LBWR(16'h0008);
TASK_LBWR(16'h0009);
TASK_PP(16'h0000,4);
TASK_PP(16'h0001,4);
TASK_PP(16'h0002,4);
TASK_PP(16'h0003,4);
TASK_PP(16'h0004,4);
TASK_PP(16'h0005,4);
TASK_PP(16'h0006,4);
TASK_PP(16'h0007,4);
TASK_PP(16'h0008,4);
TASK_PP(16'h0009,4);
TASK_PP(16'h000A,4);
TASK_PP(16'h000B,4);
TASK_PP(16'h000C,4);
TASK_PP(16'h000D,4);
TASK_PP(16'h000E,4);
TASK_PP(16'h000F,4);
TASK_PP(16'h0010,4);
TASK_PP(16'h0011,4);
TASK_PP(16'h0012,4);
TASK_PP(16'h0013,4);
TASK_PP(16'h0014,4);
TASK_PP(16'h0015,4);
TASK_PP(16'h0016,4);
TASK_PP(16'h0017,4);
TASK_PP(16'h0018,4);
TASK_PP(16'h0019,4);
TASK_PP(16'h001A,4);
TASK_PP(16'h001B,4);
TASK_PP(16'h001C,4);
TASK_PP(16'h001D,4);
TASK_PP(16'h001E,4);
TASK_PP(16'h001F,4);
TASK_PP(16'h0020,4);
TASK_PP(16'h0021,4);
TASK_PP(16'h0022,4);
TASK_PP(16'h0023,4);
TASK_PP(16'h0024,4);
TASK_PP(16'h0025,4);
TASK_PP(16'h0026,4);
TASK_PP(16'h0027,4);
TASK_PP(16'h0028,4);
TASK_PP(16'h0029,4);
TASK_PP(16'h002A,4);
TASK_PP(16'h002B,4);
TASK_PP(16'h002C,4);
TASK_PP(16'h002D,4);
TASK_PP(16'h002E,4);
TASK_PP(16'h002F,4);
TASK_PP(16'h0030,4);
TASK_PP(16'h0031,4);
TASK_PP(16'h0032,4);
TASK_PP(16'h0033,4);
TASK_PP(16'h0034,4);
TASK_PP(16'h0035,4);
TASK_PP(16'h0036,4);
TASK_PP(16'h0037,4);
TASK_PP(16'h0038,4);
TASK_PP(16'h0039,4);
TASK_PP(16'h003A,4);
TASK_PP(16'h003B,4);
TASK_PP(16'h003C,4);
TASK_PP(16'h003D,4);
TASK_PP(16'h003E,4);
TASK_PP(16'h003F,4);
TASK_PP(16'h0040,4);
TASK_PP(16'h0041,4);
TASK_PP(16'h0042,4);
TASK_PP(16'h0043,4);
TASK_PP(16'h0044,4);
TASK_PP(16'h0045,4);
TASK_PP(16'h0046,4);
TASK_PP(16'h0047,4);
TASK_PP(16'h0048,4);
TASK_PP(16'h0049,4);
TASK_PP(16'h004A,4);
TASK_PP(16'h004B,4);
TASK_PP(16'h004C,4);
TASK_PP(16'h004D,4);
TASK_PP(16'h004E,4);
TASK_PP(16'h004F,4);
TASK_PP(16'h0050,4);
TASK_PP(16'h0051,4);
TASK_PP(16'h0052,4);
TASK_PP(16'h0053,4);
TASK_PP(16'h0054,4);
TASK_PP(16'h0055,4);
TASK_PP(16'h0056,4);
TASK_PP(16'h0057,4);
TASK_PP(16'h0058,4);
TASK_PP(16'h0059,4);
TASK_PP(16'h005A,4);
TASK_PP(16'h005B,4);
TASK_PP(16'h005C,4);
TASK_PP(16'h005D,4);
TASK_PP(16'h005E,4);
TASK_PP(16'h005F,4);
TASK_PP(16'h0060,4);
TASK_PP(16'h0061,4);
TASK_PP(16'h0062,4);
TASK_PP(16'h0063,4);
TASK_PP(16'h0064,4);
TASK_PP(16'h0065,4);
TASK_PP(16'h0066,4);
TASK_PP(16'h0067,4);
TASK_PP(16'h0068,4);
TASK_PP(16'h0069,4);
TASK_PP(16'h006A,4);
TASK_PP(16'h006B,4);
TASK_PP(16'h006C,4);
TASK_PP(16'h006D,4);
TASK_PP(16'h006E,4);
TASK_PP(16'h006F,4);
TASK_PP(16'h0070,4);
TASK_PP(16'h0071,4);
TASK_PP(16'h0072,4);
TASK_PP(16'h0073,4);
TASK_PP(16'h0074,4);
TASK_PP(16'h0075,4);
TASK_PP(16'h0076,4);
TASK_PP(16'h0077,4);
TASK_PP(16'h0078,4);
TASK_PP(16'h0079,4);
TASK_PP(16'h007A,4);
TASK_PP(16'h007B,4);
TASK_PP(16'h007C,4);
TASK_PP(16'h007D,4);
TASK_PP(16'h007E,4);
TASK_PP(16'h007F,4);
TASK_PP(16'h0080,4);
TASK_PP(16'h0081,4);
TASK_PP(16'h0082,4);
TASK_PP(16'h0083,4);
TASK_PP(16'h0084,4);
TASK_PP(16'h0085,4);
TASK_PP(16'h0086,4);
TASK_PP(16'h0087,4);
TASK_PP(16'h0088,4);
TASK_PP(16'h0089,4);
TASK_PP(16'h008A,4);
TASK_PP(16'h008B,4);
TASK_PP(16'h008C,4);
TASK_PP(16'h008D,4);
TASK_PP(16'h008E,4);
TASK_PP(16'h008F,4);
TASK_PP(16'h0090,4);
TASK_PP(16'h0091,4);

// layer 0
TASK_ACCRST;
TASK_MACCYC(0,32'h00000000);
TASK_MACCYC(0,32'h00010001);
TASK_MACCYC(0,32'h00020002);
TASK_MACCYC(0,32'h00030003);
TASK_MACCYC(0,32'h00040004);
TASK_MACCYC(0,32'h00050005);
TASK_MACCYC(0,32'h00060006);
TASK_MACCYC(0,32'h00070007);
TASK_MACCYC(0,32'h00080008);
TASK_MACCYC(0,32'h00090009);
TASK_BIASBUF(4,16'h000A);
TASK_NEURONACT(32'h000003F1);
TASK_NEURONACT(32'h000103F2);
TASK_NEURONACT(32'h000203F3);
TASK_NEURONACT(32'h000303F4);
TASK_ACCRST;
TASK_MACCYC(0,32'h000E0000);
TASK_MACCYC(0,32'h000F0001);
TASK_MACCYC(0,32'h00100002);
TASK_MACCYC(0,32'h00110003);
TASK_MACCYC(0,32'h00120004);
TASK_MACCYC(0,32'h00130005);
TASK_MACCYC(0,32'h00140006);
TASK_MACCYC(0,32'h00150007);
TASK_MACCYC(0,32'h00160008);
TASK_MACCYC(0,32'h00170009);
TASK_BIASBUF(4,16'h0018);
TASK_NEURONACT(32'h000003F5);
TASK_NEURONACT(32'h000103F6);
TASK_NEURONACT(32'h000203F7);
TASK_NEURONACT(32'h000303F8);
TASK_ACCRST;
TASK_MACCYC(0,32'h001C0000);
TASK_MACCYC(0,32'h001D0001);
TASK_MACCYC(0,32'h001E0002);
TASK_MACCYC(0,32'h001F0003);
TASK_MACCYC(0,32'h00200004);
TASK_MACCYC(0,32'h00210005);
TASK_MACCYC(0,32'h00220006);
TASK_MACCYC(0,32'h00230007);
TASK_MACCYC(0,32'h00240008);
TASK_MACCYC(0,32'h00250009);
TASK_BIASBUF(4,16'h0026);
TASK_NEURONACT(32'h000003F9);
TASK_NEURONACT(32'h000103FA);
TASK_NEURONACT(32'h000203FB);
TASK_NEURONACT(32'h000303FC);
TASK_ACCRST;
TASK_MACCYC(0,32'h002A0000);
TASK_MACCYC(0,32'h002B0001);
TASK_MACCYC(0,32'h002C0002);
TASK_MACCYC(0,32'h002D0003);
TASK_MACCYC(0,32'h002E0004);
TASK_MACCYC(0,32'h002F0005);
TASK_MACCYC(0,32'h00300006);
TASK_MACCYC(0,32'h00310007);
TASK_MACCYC(0,32'h00320008);
TASK_MACCYC(0,32'h00330009);
TASK_BIASBUF(4,16'h0034);
TASK_NEURONACT(32'h000003FD);
TASK_NEURONACT(32'h000103FE);
TASK_NEURONACT(32'h000203FF);
TASK_ACCRST;

// layer 1
TASK_ACCRST;
TASK_MACCYC(0,32'h003803F1);
TASK_MACCYC(0,32'h003903F2);
TASK_MACCYC(0,32'h003A03F3);
TASK_MACCYC(0,32'h003B03F4);
TASK_MACCYC(0,32'h003C03F5);
TASK_MACCYC(0,32'h003D03F6);
TASK_MACCYC(0,32'h003E03F7);
TASK_MACCYC(0,32'h003F03F8);
TASK_MACCYC(0,32'h004003F9);
TASK_MACCYC(0,32'h004103FA);
TASK_MACCYC(0,32'h004203FB);
TASK_MACCYC(0,32'h004303FC);
TASK_MACCYC(0,32'h004403FD);
TASK_MACCYC(0,32'h004503FE);
TASK_MACCYC(0,32'h004603FF);
TASK_BIASBUF(4,16'h0047);
TASK_NEURONACT(32'h00000000);
TASK_NEURONACT(32'h00010001);
TASK_NEURONACT(32'h00020002);
TASK_NEURONACT(32'h00030003);
TASK_ACCRST;
TASK_MACCYC(0,32'h004B03F1);
TASK_MACCYC(0,32'h004C03F2);
TASK_MACCYC(0,32'h004D03F3);
TASK_MACCYC(0,32'h004E03F4);
TASK_MACCYC(0,32'h004F03F5);
TASK_MACCYC(0,32'h005003F6);
TASK_MACCYC(0,32'h005103F7);
TASK_MACCYC(0,32'h005203F8);
TASK_MACCYC(0,32'h005303F9);
TASK_MACCYC(0,32'h005403FA);
TASK_MACCYC(0,32'h005503FB);
TASK_MACCYC(0,32'h005603FC);
TASK_MACCYC(0,32'h005703FD);
TASK_MACCYC(0,32'h005803FE);
TASK_MACCYC(0,32'h005903FF);
TASK_BIASBUF(4,16'h005A);
TASK_NEURONACT(32'h00000004);
TASK_NEURONACT(32'h00010005);
TASK_NEURONACT(32'h00020006);
TASK_NEURONACT(32'h00030007);
TASK_ACCRST;

// layer 2
TASK_ACCRST;
TASK_MACCYC(0,32'h005E0000);
TASK_MACCYC(0,32'h005F0001);
TASK_MACCYC(0,32'h00600002);
TASK_MACCYC(0,32'h00610003);
TASK_MACCYC(0,32'h00620004);
TASK_MACCYC(0,32'h00630005);
TASK_MACCYC(0,32'h00640006);
TASK_MACCYC(0,32'h00650007);
TASK_BIASBUF(4,16'h0066);
TASK_NEURONACT(32'h000003F4);
TASK_NEURONACT(32'h000103F5);
TASK_NEURONACT(32'h000203F6);
TASK_NEURONACT(32'h000303F7);
TASK_ACCRST;
TASK_MACCYC(0,32'h006A0000);
TASK_MACCYC(0,32'h006B0001);
TASK_MACCYC(0,32'h006C0002);
TASK_MACCYC(0,32'h006D0003);
TASK_MACCYC(0,32'h006E0004);
TASK_MACCYC(0,32'h006F0005);
TASK_MACCYC(0,32'h00700006);
TASK_MACCYC(0,32'h00710007);
TASK_BIASBUF(4,16'h0072);
TASK_NEURONACT(32'h000003F8);
TASK_NEURONACT(32'h000103F9);
TASK_NEURONACT(32'h000203FA);
TASK_NEURONACT(32'h000303FB);
TASK_ACCRST;
TASK_MACCYC(0,32'h00760000);
TASK_MACCYC(0,32'h00770001);
TASK_MACCYC(0,32'h00780002);
TASK_MACCYC(0,32'h00790003);
TASK_MACCYC(0,32'h007A0004);
TASK_MACCYC(0,32'h007B0005);
TASK_MACCYC(0,32'h007C0006);
TASK_MACCYC(0,32'h007D0007);
TASK_BIASBUF(4,16'h007E);
TASK_NEURONACT(32'h000003FC);
TASK_NEURONACT(32'h000103FD);
TASK_NEURONACT(32'h000203FE);
TASK_NEURONACT(32'h000303FF);
TASK_ACCRST;

// layer 3
TASK_ACCRST;
TASK_MACCYC(0,32'h008203F4);
TASK_MACCYC(0,32'h008303F5);
TASK_MACCYC(0,32'h008403F6);
TASK_MACCYC(0,32'h008503F7);
TASK_MACCYC(0,32'h008603F8);
TASK_MACCYC(0,32'h008703F9);
TASK_MACCYC(0,32'h008803FA);
TASK_MACCYC(0,32'h008903FB);
TASK_MACCYC(0,32'h008A03FC);
TASK_MACCYC(0,32'h008B03FD);
TASK_MACCYC(0,32'h008C03FE);
TASK_MACCYC(0,32'h008D03FF);
TASK_BIASBUF(4,16'h008E);
TASK_NEURONACT(32'h00000000);
TASK_NEURONACT(32'h00010001);
TASK_NEURONACT(32'h00020002);
TASK_NEURONACT(32'h00030003);
TASK_ACCRST;
