`include "./banners/+runP_start.vh"
`include "./banners/+test1.vh"
TASK_RSTEN;
TASK_RST;
TASK_INIT_WRITE_PI;
TASK_LBWR(16'h0000);
TASK_LBWR(16'h0001);
TASK_LBWR(16'h0002);
TASK_LBWR(16'h0003);
TASK_LBWR(16'h0004);
TASK_LBWR(16'h0005);
TASK_LBWR(16'h0006);
TASK_LBWR(16'h0007);
TASK_LBWR(16'h0008);
TASK_LBWR(16'h0009);
TASK_LBWR(16'h000A);
TASK_LBWR(16'h000B);
TASK_LBWR(16'h000C);
TASK_LBWR(16'h000D);
TASK_LBWR(16'h000E);
TASK_LBWR(16'h000F);
TASK_LBWR(16'h0010);
TASK_LBWR(16'h0011);
TASK_LBWR(16'h0012);
TASK_LBWR(16'h0013);
TASK_LBWR(16'h0014);
TASK_LBWR(16'h0015);
TASK_LBWR(16'h0016);
TASK_LBWR(16'h0017);
TASK_LBWR(16'h0018);
TASK_LBWR(16'h0019);
TASK_LBWR(16'h001A);
TASK_LBWR(16'h001B);
TASK_LBWR(16'h001C);
TASK_LBWR(16'h001D);
TASK_LBWR(16'h001E);
TASK_LBWR(16'h001F);
TASK_LBWR(16'h0020);
TASK_LBWR(16'h0021);
TASK_LBWR(16'h0022);
TASK_LBWR(16'h0023);
TASK_LBWR(16'h0024);
TASK_LBWR(16'h0025);
TASK_LBWR(16'h0026);
TASK_LBWR(16'h0027);
TASK_LBWR(16'h0028);
TASK_LBWR(16'h0029);
TASK_LBWR(16'h002A);
TASK_LBWR(16'h002B);
TASK_LBWR(16'h002C);
TASK_LBWR(16'h002D);
TASK_LBWR(16'h002E);
TASK_LBWR(16'h002F);
TASK_LBWR(16'h0030);
TASK_LBWR(16'h0031);
TASK_LBWR(16'h0032);
TASK_LBWR(16'h0033);
TASK_LBWR(16'h0034);
TASK_LBWR(16'h0035);
TASK_LBWR(16'h0036);
TASK_LBWR(16'h0037);
TASK_LBWR(16'h0038);
TASK_LBWR(16'h0039);
TASK_LBWR(16'h003A);
TASK_LBWR(16'h003B);
TASK_LBWR(16'h003C);
TASK_LBWR(16'h003D);
TASK_LBWR(16'h003E);
TASK_LBWR(16'h003F);
TASK_LBWR(16'h0040);
TASK_LBWR(16'h0041);
TASK_LBWR(16'h0042);
TASK_LBWR(16'h0043);
TASK_LBWR(16'h0044);
TASK_LBWR(16'h0045);
TASK_LBWR(16'h0046);
TASK_LBWR(16'h0047);
TASK_LBWR(16'h0048);
TASK_LBWR(16'h0049);
TASK_LBWR(16'h004A);
TASK_LBWR(16'h004B);
TASK_LBWR(16'h004C);
TASK_LBWR(16'h004D);
TASK_LBWR(16'h004E);
TASK_LBWR(16'h004F);
TASK_LBWR(16'h0050);
TASK_LBWR(16'h0051);
TASK_LBWR(16'h0052);
TASK_LBWR(16'h0053);
TASK_LBWR(16'h0054);
TASK_LBWR(16'h0055);
TASK_LBWR(16'h0056);
TASK_LBWR(16'h0057);
TASK_LBWR(16'h0058);
TASK_LBWR(16'h0059);
TASK_LBWR(16'h005A);
TASK_LBWR(16'h005B);
TASK_LBWR(16'h005C);
TASK_LBWR(16'h005D);
TASK_LBWR(16'h005E);
TASK_LBWR(16'h005F);
TASK_LBWR(16'h0060);
TASK_LBWR(16'h0061);
TASK_LBWR(16'h0062);
TASK_LBWR(16'h0063);
TASK_LBWR(16'h0064);
TASK_LBWR(16'h0065);
TASK_LBWR(16'h0066);
TASK_LBWR(16'h0067);
TASK_LBWR(16'h0068);
TASK_LBWR(16'h0069);
TASK_LBWR(16'h006A);
TASK_LBWR(16'h006B);
TASK_LBWR(16'h006C);
TASK_LBWR(16'h006D);
TASK_LBWR(16'h006E);
TASK_LBWR(16'h006F);
TASK_LBWR(16'h0070);
TASK_LBWR(16'h0071);
TASK_LBWR(16'h0072);
TASK_LBWR(16'h0073);
TASK_LBWR(16'h0074);
TASK_LBWR(16'h0075);
TASK_LBWR(16'h0076);
TASK_LBWR(16'h0077);
TASK_LBWR(16'h0078);
TASK_LBWR(16'h0079);
TASK_LBWR(16'h007A);
TASK_LBWR(16'h007B);
TASK_LBWR(16'h007C);
TASK_LBWR(16'h007D);
TASK_LBWR(16'h007E);
TASK_LBWR(16'h007F);
TASK_LBWR(16'h0080);
TASK_LBWR(16'h0081);
TASK_LBWR(16'h0082);
TASK_LBWR(16'h0083);
TASK_LBWR(16'h0084);
TASK_LBWR(16'h0085);
TASK_LBWR(16'h0086);
TASK_LBWR(16'h0087);
TASK_LBWR(16'h0088);
TASK_LBWR(16'h0089);
TASK_LBWR(16'h008A);
TASK_LBWR(16'h008B);
TASK_LBWR(16'h008C);
TASK_LBWR(16'h008D);
TASK_LBWR(16'h008E);
TASK_LBWR(16'h008F);
TASK_LBWR(16'h0090);
TASK_LBWR(16'h0091);
TASK_LBWR(16'h0092);
TASK_LBWR(16'h0093);
TASK_LBWR(16'h0094);
TASK_LBWR(16'h0095);
TASK_LBWR(16'h0096);
TASK_LBWR(16'h0097);
TASK_LBWR(16'h0098);
TASK_LBWR(16'h0099);
TASK_LBWR(16'h009A);
TASK_LBWR(16'h009B);
TASK_LBWR(16'h009C);
TASK_LBWR(16'h009D);
TASK_LBWR(16'h009E);
TASK_LBWR(16'h009F);
TASK_LBWR(16'h00A0);
TASK_LBWR(16'h00A1);
TASK_LBWR(16'h00A2);
TASK_LBWR(16'h00A3);
TASK_LBWR(16'h00A4);
TASK_LBWR(16'h00A5);
TASK_LBWR(16'h00A6);
TASK_LBWR(16'h00A7);
TASK_LBWR(16'h00A8);
TASK_LBWR(16'h00A9);
TASK_LBWR(16'h00AA);
TASK_LBWR(16'h00AB);
TASK_LBWR(16'h00AC);
TASK_LBWR(16'h00AD);
TASK_LBWR(16'h00AE);
TASK_LBWR(16'h00AF);
TASK_LBWR(16'h00B0);
TASK_LBWR(16'h00B1);
TASK_LBWR(16'h00B2);
TASK_LBWR(16'h00B3);
TASK_LBWR(16'h00B4);
TASK_LBWR(16'h00B5);
TASK_LBWR(16'h00B6);
TASK_LBWR(16'h00B7);
TASK_LBWR(16'h00B8);
TASK_LBWR(16'h00B9);
TASK_LBWR(16'h00BA);
TASK_LBWR(16'h00BB);
TASK_LBWR(16'h00BC);
TASK_LBWR(16'h00BD);
TASK_LBWR(16'h00BE);
TASK_LBWR(16'h00BF);
TASK_LBWR(16'h00C0);
TASK_LBWR(16'h00C1);
TASK_LBWR(16'h00C2);
TASK_LBWR(16'h00C3);
TASK_LBWR(16'h00C4);
TASK_LBWR(16'h00C5);
TASK_LBWR(16'h00C6);
TASK_LBWR(16'h00C7);
TASK_LBWR(16'h00C8);
TASK_LBWR(16'h00C9);
TASK_LBWR(16'h00CA);
TASK_LBWR(16'h00CB);
TASK_LBWR(16'h00CC);
TASK_LBWR(16'h00CD);
TASK_LBWR(16'h00CE);
TASK_LBWR(16'h00CF);
TASK_LBWR(16'h00D0);
TASK_LBWR(16'h00D1);
TASK_LBWR(16'h00D2);
TASK_LBWR(16'h00D3);
TASK_LBWR(16'h00D4);
TASK_LBWR(16'h00D5);
TASK_LBWR(16'h00D6);
TASK_LBWR(16'h00D7);
TASK_LBWR(16'h00D8);
TASK_LBWR(16'h00D9);
TASK_LBWR(16'h00DA);
TASK_LBWR(16'h00DB);
TASK_LBWR(16'h00DC);
TASK_LBWR(16'h00DD);
TASK_LBWR(16'h00DE);
TASK_LBWR(16'h00DF);
TASK_LBWR(16'h00E0);
TASK_LBWR(16'h00E1);
TASK_LBWR(16'h00E2);
TASK_LBWR(16'h00E3);
TASK_LBWR(16'h00E4);
TASK_LBWR(16'h00E5);
TASK_LBWR(16'h00E6);
TASK_LBWR(16'h00E7);
TASK_LBWR(16'h00E8);
TASK_LBWR(16'h00E9);
TASK_LBWR(16'h00EA);
TASK_LBWR(16'h00EB);
TASK_LBWR(16'h00EC);
TASK_LBWR(16'h00ED);
TASK_LBWR(16'h00EE);
TASK_LBWR(16'h00EF);
TASK_LBWR(16'h00F0);
TASK_LBWR(16'h00F1);
TASK_LBWR(16'h00F2);
TASK_LBWR(16'h00F3);
TASK_LBWR(16'h00F4);
TASK_LBWR(16'h00F5);
TASK_LBWR(16'h00F6);
TASK_LBWR(16'h00F7);
TASK_LBWR(16'h00F8);
TASK_LBWR(16'h00F9);
TASK_LBWR(16'h00FA);
TASK_LBWR(16'h00FB);
TASK_LBWR(16'h00FC);
TASK_LBWR(16'h00FD);
TASK_LBWR(16'h00FE);
TASK_LBWR(16'h00FF);
TASK_LBWR(16'h0100);
TASK_LBWR(16'h0101);
TASK_LBWR(16'h0102);
TASK_LBWR(16'h0103);
TASK_LBWR(16'h0104);
TASK_LBWR(16'h0105);
TASK_LBWR(16'h0106);
TASK_LBWR(16'h0107);
TASK_LBWR(16'h0108);
TASK_LBWR(16'h0109);
TASK_LBWR(16'h010A);
TASK_LBWR(16'h010B);
TASK_LBWR(16'h010C);
TASK_LBWR(16'h010D);
TASK_LBWR(16'h010E);
TASK_LBWR(16'h010F);
TASK_LBWR(16'h0110);
TASK_LBWR(16'h0111);
TASK_LBWR(16'h0112);
TASK_LBWR(16'h0113);
TASK_LBWR(16'h0114);
TASK_LBWR(16'h0115);
TASK_LBWR(16'h0116);
TASK_LBWR(16'h0117);
TASK_LBWR(16'h0118);
TASK_LBWR(16'h0119);
TASK_LBWR(16'h011A);
TASK_LBWR(16'h011B);
TASK_LBWR(16'h011C);
TASK_LBWR(16'h011D);
TASK_LBWR(16'h011E);
TASK_LBWR(16'h011F);
TASK_LBWR(16'h0120);
TASK_LBWR(16'h0121);
TASK_LBWR(16'h0122);
TASK_LBWR(16'h0123);
TASK_LBWR(16'h0124);
TASK_LBWR(16'h0125);
TASK_LBWR(16'h0126);
TASK_LBWR(16'h0127);
TASK_LBWR(16'h0128);
TASK_LBWR(16'h0129);
TASK_LBWR(16'h012A);
TASK_LBWR(16'h012B);
TASK_LBWR(16'h012C);
TASK_LBWR(16'h012D);
TASK_LBWR(16'h012E);
TASK_LBWR(16'h012F);
TASK_LBWR(16'h0130);
TASK_LBWR(16'h0131);
TASK_LBWR(16'h0132);
TASK_LBWR(16'h0133);
TASK_LBWR(16'h0134);
TASK_LBWR(16'h0135);
TASK_LBWR(16'h0136);
TASK_LBWR(16'h0137);
TASK_LBWR(16'h0138);
TASK_LBWR(16'h0139);
TASK_LBWR(16'h013A);
TASK_LBWR(16'h013B);
TASK_LBWR(16'h013C);
TASK_LBWR(16'h013D);
TASK_LBWR(16'h013E);
TASK_LBWR(16'h013F);
TASK_LBWR(16'h0140);
TASK_LBWR(16'h0141);
TASK_LBWR(16'h0142);
TASK_LBWR(16'h0143);
TASK_LBWR(16'h0144);
TASK_LBWR(16'h0145);
TASK_LBWR(16'h0146);
TASK_LBWR(16'h0147);
TASK_LBWR(16'h0148);
TASK_LBWR(16'h0149);
TASK_LBWR(16'h014A);
TASK_LBWR(16'h014B);
TASK_LBWR(16'h014C);
TASK_LBWR(16'h014D);
TASK_LBWR(16'h014E);
TASK_LBWR(16'h014F);
TASK_LBWR(16'h0150);
TASK_LBWR(16'h0151);
TASK_LBWR(16'h0152);
TASK_LBWR(16'h0153);
TASK_LBWR(16'h0154);
TASK_LBWR(16'h0155);
TASK_LBWR(16'h0156);
TASK_LBWR(16'h0157);
TASK_LBWR(16'h0158);
TASK_LBWR(16'h0159);
TASK_LBWR(16'h015A);
TASK_LBWR(16'h015B);
TASK_LBWR(16'h015C);
TASK_LBWR(16'h015D);
TASK_LBWR(16'h015E);
TASK_LBWR(16'h015F);
TASK_LBWR(16'h0160);
TASK_LBWR(16'h0161);
TASK_LBWR(16'h0162);
TASK_LBWR(16'h0163);
TASK_LBWR(16'h0164);
TASK_LBWR(16'h0165);
TASK_LBWR(16'h0166);
TASK_LBWR(16'h0167);
TASK_LBWR(16'h0168);
TASK_LBWR(16'h0169);
TASK_LBWR(16'h016A);
TASK_LBWR(16'h016B);
TASK_LBWR(16'h016C);
TASK_LBWR(16'h016D);
TASK_LBWR(16'h016E);
TASK_LBWR(16'h016F);
TASK_LBWR(16'h0170);
TASK_LBWR(16'h0171);
TASK_LBWR(16'h0172);
TASK_LBWR(16'h0173);
TASK_LBWR(16'h0174);
TASK_LBWR(16'h0175);
TASK_LBWR(16'h0176);
TASK_LBWR(16'h0177);
TASK_LBWR(16'h0178);
TASK_LBWR(16'h0179);
TASK_LBWR(16'h017A);
TASK_LBWR(16'h017B);
TASK_LBWR(16'h017C);
TASK_LBWR(16'h017D);
TASK_LBWR(16'h017E);
TASK_LBWR(16'h017F);
TASK_LBWR(16'h0180);
TASK_LBWR(16'h0181);
TASK_LBWR(16'h0182);
TASK_LBWR(16'h0183);
TASK_LBWR(16'h0184);
TASK_LBWR(16'h0185);
TASK_LBWR(16'h0186);
TASK_LBWR(16'h0187);
TASK_LBWR(16'h0188);
TASK_LBWR(16'h0189);
TASK_LBWR(16'h018A);
TASK_LBWR(16'h018B);
TASK_LBWR(16'h018C);
TASK_LBWR(16'h018D);
TASK_LBWR(16'h018E);
TASK_LBWR(16'h018F);
TASK_LBWR(16'h0190);
TASK_LBWR(16'h0191);
TASK_LBWR(16'h0192);
TASK_LBWR(16'h0193);
TASK_LBWR(16'h0194);
TASK_LBWR(16'h0195);
TASK_LBWR(16'h0196);
TASK_LBWR(16'h0197);
TASK_LBWR(16'h0198);
TASK_LBWR(16'h0199);
TASK_LBWR(16'h019A);
TASK_LBWR(16'h019B);
TASK_LBWR(16'h019C);
TASK_LBWR(16'h019D);
TASK_LBWR(16'h019E);
TASK_LBWR(16'h019F);
TASK_LBWR(16'h01A0);
TASK_LBWR(16'h01A1);
TASK_LBWR(16'h01A2);
TASK_LBWR(16'h01A3);
TASK_LBWR(16'h01A4);
TASK_LBWR(16'h01A5);
TASK_LBWR(16'h01A6);
TASK_LBWR(16'h01A7);
TASK_LBWR(16'h01A8);
TASK_LBWR(16'h01A9);
TASK_LBWR(16'h01AA);
TASK_LBWR(16'h01AB);
TASK_LBWR(16'h01AC);
TASK_LBWR(16'h01AD);
TASK_LBWR(16'h01AE);
TASK_LBWR(16'h01AF);
TASK_LBWR(16'h01B0);
TASK_LBWR(16'h01B1);
TASK_LBWR(16'h01B2);
TASK_LBWR(16'h01B3);
TASK_LBWR(16'h01B4);
TASK_LBWR(16'h01B5);
TASK_LBWR(16'h01B6);
TASK_LBWR(16'h01B7);
TASK_LBWR(16'h01B8);
TASK_LBWR(16'h01B9);
TASK_LBWR(16'h01BA);
TASK_LBWR(16'h01BB);
TASK_LBWR(16'h01BC);
TASK_LBWR(16'h01BD);
TASK_LBWR(16'h01BE);
TASK_LBWR(16'h01BF);
TASK_LBWR(16'h01C0);
TASK_LBWR(16'h01C1);
TASK_LBWR(16'h01C2);
TASK_LBWR(16'h01C3);
TASK_LBWR(16'h01C4);
TASK_LBWR(16'h01C5);
TASK_LBWR(16'h01C6);
TASK_LBWR(16'h01C7);
TASK_LBWR(16'h01C8);
TASK_LBWR(16'h01C9);
TASK_LBWR(16'h01CA);
TASK_LBWR(16'h01CB);
TASK_LBWR(16'h01CC);
TASK_LBWR(16'h01CD);
TASK_LBWR(16'h01CE);
TASK_LBWR(16'h01CF);
TASK_LBWR(16'h01D0);
TASK_LBWR(16'h01D1);
TASK_LBWR(16'h01D2);
TASK_LBWR(16'h01D3);
TASK_LBWR(16'h01D4);
TASK_LBWR(16'h01D5);
TASK_LBWR(16'h01D6);
TASK_LBWR(16'h01D7);
TASK_LBWR(16'h01D8);
TASK_LBWR(16'h01D9);
TASK_LBWR(16'h01DA);
TASK_LBWR(16'h01DB);
TASK_LBWR(16'h01DC);
TASK_LBWR(16'h01DD);
TASK_LBWR(16'h01DE);
TASK_LBWR(16'h01DF);
TASK_LBWR(16'h01E0);
TASK_LBWR(16'h01E1);
TASK_LBWR(16'h01E2);
TASK_LBWR(16'h01E3);
TASK_LBWR(16'h01E4);
TASK_LBWR(16'h01E5);
TASK_LBWR(16'h01E6);
TASK_LBWR(16'h01E7);
TASK_LBWR(16'h01E8);
TASK_LBWR(16'h01E9);
TASK_LBWR(16'h01EA);
TASK_LBWR(16'h01EB);
TASK_LBWR(16'h01EC);
TASK_LBWR(16'h01ED);
TASK_LBWR(16'h01EE);
TASK_LBWR(16'h01EF);
TASK_LBWR(16'h01F0);
TASK_LBWR(16'h01F1);
TASK_LBWR(16'h01F2);
TASK_LBWR(16'h01F3);
TASK_LBWR(16'h01F4);
TASK_LBWR(16'h01F5);
TASK_LBWR(16'h01F6);
TASK_LBWR(16'h01F7);
TASK_LBWR(16'h01F8);
TASK_LBWR(16'h01F9);
TASK_LBWR(16'h01FA);
TASK_LBWR(16'h01FB);
TASK_LBWR(16'h01FC);
TASK_LBWR(16'h01FD);
TASK_LBWR(16'h01FE);
TASK_LBWR(16'h01FF);
TASK_LBWR(16'h0200);
TASK_LBWR(16'h0201);
TASK_LBWR(16'h0202);
TASK_LBWR(16'h0203);
TASK_LBWR(16'h0204);
TASK_LBWR(16'h0205);
TASK_LBWR(16'h0206);
TASK_LBWR(16'h0207);
TASK_LBWR(16'h0208);
TASK_LBWR(16'h0209);
TASK_LBWR(16'h020A);
TASK_LBWR(16'h020B);
TASK_LBWR(16'h020C);
TASK_LBWR(16'h020D);
TASK_LBWR(16'h020E);
TASK_LBWR(16'h020F);
TASK_LBWR(16'h0210);
TASK_LBWR(16'h0211);
TASK_LBWR(16'h0212);
TASK_LBWR(16'h0213);
TASK_LBWR(16'h0214);
TASK_LBWR(16'h0215);
TASK_LBWR(16'h0216);
TASK_LBWR(16'h0217);
TASK_LBWR(16'h0218);
TASK_LBWR(16'h0219);
TASK_LBWR(16'h021A);
TASK_LBWR(16'h021B);
TASK_LBWR(16'h021C);
TASK_LBWR(16'h021D);
TASK_LBWR(16'h021E);
TASK_LBWR(16'h021F);
TASK_LBWR(16'h0220);
TASK_LBWR(16'h0221);
TASK_LBWR(16'h0222);
TASK_LBWR(16'h0223);
TASK_LBWR(16'h0224);
TASK_LBWR(16'h0225);
TASK_LBWR(16'h0226);
TASK_LBWR(16'h0227);
TASK_LBWR(16'h0228);
TASK_LBWR(16'h0229);
TASK_LBWR(16'h022A);
TASK_LBWR(16'h022B);
TASK_LBWR(16'h022C);
TASK_LBWR(16'h022D);
TASK_LBWR(16'h022E);
TASK_LBWR(16'h022F);
TASK_LBWR(16'h0230);
TASK_LBWR(16'h0231);
TASK_LBWR(16'h0232);
TASK_LBWR(16'h0233);
TASK_LBWR(16'h0234);
TASK_LBWR(16'h0235);
TASK_LBWR(16'h0236);
TASK_LBWR(16'h0237);
TASK_LBWR(16'h0238);
TASK_LBWR(16'h0239);
TASK_LBWR(16'h023A);
TASK_LBWR(16'h023B);
TASK_LBWR(16'h023C);
TASK_LBWR(16'h023D);
TASK_LBWR(16'h023E);
TASK_LBWR(16'h023F);
TASK_LBWR(16'h0240);
TASK_LBWR(16'h0241);
TASK_LBWR(16'h0242);
TASK_LBWR(16'h0243);
TASK_LBWR(16'h0244);
TASK_LBWR(16'h0245);
TASK_LBWR(16'h0246);
TASK_LBWR(16'h0247);
TASK_LBWR(16'h0248);
TASK_LBWR(16'h0249);
TASK_LBWR(16'h024A);
TASK_LBWR(16'h024B);
TASK_LBWR(16'h024C);
TASK_LBWR(16'h024D);
TASK_LBWR(16'h024E);
TASK_LBWR(16'h024F);
TASK_LBWR(16'h0250);
TASK_LBWR(16'h0251);
TASK_LBWR(16'h0252);
TASK_LBWR(16'h0253);
TASK_LBWR(16'h0254);
TASK_LBWR(16'h0255);
TASK_LBWR(16'h0256);
TASK_LBWR(16'h0257);
TASK_LBWR(16'h0258);
TASK_LBWR(16'h0259);
TASK_LBWR(16'h025A);
TASK_LBWR(16'h025B);
TASK_LBWR(16'h025C);
TASK_LBWR(16'h025D);
TASK_LBWR(16'h025E);
TASK_LBWR(16'h025F);
TASK_LBWR(16'h0260);
TASK_LBWR(16'h0261);
TASK_LBWR(16'h0262);
TASK_LBWR(16'h0263);
TASK_LBWR(16'h0264);
TASK_LBWR(16'h0265);
TASK_LBWR(16'h0266);
TASK_LBWR(16'h0267);
TASK_LBWR(16'h0268);
TASK_LBWR(16'h0269);
TASK_LBWR(16'h026A);
TASK_LBWR(16'h026B);
TASK_LBWR(16'h026C);
TASK_LBWR(16'h026D);
TASK_LBWR(16'h026E);
TASK_LBWR(16'h026F);
TASK_LBWR(16'h0270);
TASK_LBWR(16'h0271);
TASK_LBWR(16'h0272);
TASK_LBWR(16'h0273);
TASK_LBWR(16'h0274);
TASK_LBWR(16'h0275);
TASK_LBWR(16'h0276);
TASK_LBWR(16'h0277);
TASK_LBWR(16'h0278);
TASK_LBWR(16'h0279);
TASK_LBWR(16'h027A);
TASK_LBWR(16'h027B);
TASK_LBWR(16'h027C);
TASK_LBWR(16'h027D);
TASK_LBWR(16'h027E);
TASK_LBWR(16'h027F);
TASK_LBWR(16'h0280);
TASK_LBWR(16'h0281);
TASK_LBWR(16'h0282);
TASK_LBWR(16'h0283);
TASK_LBWR(16'h0284);
TASK_LBWR(16'h0285);
TASK_LBWR(16'h0286);
TASK_LBWR(16'h0287);
TASK_LBWR(16'h0288);
TASK_LBWR(16'h0289);
TASK_LBWR(16'h028A);
TASK_LBWR(16'h028B);
TASK_LBWR(16'h028C);
TASK_LBWR(16'h028D);
TASK_LBWR(16'h028E);
TASK_LBWR(16'h028F);
TASK_LBWR(16'h0290);
TASK_LBWR(16'h0291);
TASK_LBWR(16'h0292);
TASK_LBWR(16'h0293);
TASK_LBWR(16'h0294);
TASK_LBWR(16'h0295);
TASK_LBWR(16'h0296);
TASK_LBWR(16'h0297);
TASK_LBWR(16'h0298);
TASK_LBWR(16'h0299);
TASK_LBWR(16'h029A);
TASK_LBWR(16'h029B);
TASK_LBWR(16'h029C);
TASK_LBWR(16'h029D);
TASK_LBWR(16'h029E);
TASK_LBWR(16'h029F);
TASK_LBWR(16'h02A0);
TASK_LBWR(16'h02A1);
TASK_LBWR(16'h02A2);
TASK_LBWR(16'h02A3);
TASK_LBWR(16'h02A4);
TASK_LBWR(16'h02A5);
TASK_LBWR(16'h02A6);
TASK_LBWR(16'h02A7);
TASK_LBWR(16'h02A8);
TASK_LBWR(16'h02A9);
TASK_LBWR(16'h02AA);
TASK_LBWR(16'h02AB);
TASK_LBWR(16'h02AC);
TASK_LBWR(16'h02AD);
TASK_LBWR(16'h02AE);
TASK_LBWR(16'h02AF);
TASK_LBWR(16'h02B0);
TASK_LBWR(16'h02B1);
TASK_LBWR(16'h02B2);
TASK_LBWR(16'h02B3);
TASK_LBWR(16'h02B4);
TASK_LBWR(16'h02B5);
TASK_LBWR(16'h02B6);
TASK_LBWR(16'h02B7);
TASK_LBWR(16'h02B8);
TASK_LBWR(16'h02B9);
TASK_LBWR(16'h02BA);
TASK_LBWR(16'h02BB);
TASK_LBWR(16'h02BC);
TASK_LBWR(16'h02BD);
TASK_LBWR(16'h02BE);
TASK_LBWR(16'h02BF);
TASK_LBWR(16'h02C0);
TASK_LBWR(16'h02C1);
TASK_LBWR(16'h02C2);
TASK_LBWR(16'h02C3);
TASK_LBWR(16'h02C4);
TASK_LBWR(16'h02C5);
TASK_LBWR(16'h02C6);
TASK_LBWR(16'h02C7);
TASK_LBWR(16'h02C8);
TASK_LBWR(16'h02C9);
TASK_LBWR(16'h02CA);
TASK_LBWR(16'h02CB);
TASK_LBWR(16'h02CC);
TASK_LBWR(16'h02CD);
TASK_LBWR(16'h02CE);
TASK_LBWR(16'h02CF);
TASK_LBWR(16'h02D0);
TASK_LBWR(16'h02D1);
TASK_LBWR(16'h02D2);
TASK_LBWR(16'h02D3);
TASK_LBWR(16'h02D4);
TASK_LBWR(16'h02D5);
TASK_LBWR(16'h02D6);
TASK_LBWR(16'h02D7);
TASK_LBWR(16'h02D8);
TASK_LBWR(16'h02D9);
TASK_LBWR(16'h02DA);
TASK_LBWR(16'h02DB);
TASK_LBWR(16'h02DC);
TASK_LBWR(16'h02DD);
TASK_LBWR(16'h02DE);
TASK_LBWR(16'h02DF);
TASK_LBWR(16'h02E0);
TASK_LBWR(16'h02E1);
TASK_LBWR(16'h02E2);
TASK_LBWR(16'h02E3);
TASK_LBWR(16'h02E4);
TASK_LBWR(16'h02E5);
TASK_LBWR(16'h02E6);
TASK_LBWR(16'h02E7);
TASK_LBWR(16'h02E8);
TASK_LBWR(16'h02E9);
TASK_LBWR(16'h02EA);
TASK_LBWR(16'h02EB);
TASK_LBWR(16'h02EC);
TASK_LBWR(16'h02ED);
TASK_LBWR(16'h02EE);
TASK_LBWR(16'h02EF);
TASK_LBWR(16'h02F0);
TASK_LBWR(16'h02F1);
TASK_LBWR(16'h02F2);
TASK_LBWR(16'h02F3);
TASK_LBWR(16'h02F4);
TASK_LBWR(16'h02F5);
TASK_LBWR(16'h02F6);
TASK_LBWR(16'h02F7);
TASK_LBWR(16'h02F8);
TASK_LBWR(16'h02F9);
TASK_LBWR(16'h02FA);
TASK_LBWR(16'h02FB);
TASK_LBWR(16'h02FC);
TASK_LBWR(16'h02FD);
TASK_LBWR(16'h02FE);
TASK_LBWR(16'h02FF);
TASK_LBWR(16'h0300);
TASK_LBWR(16'h0301);
TASK_LBWR(16'h0302);
TASK_LBWR(16'h0303);
TASK_LBWR(16'h0304);
TASK_LBWR(16'h0305);
TASK_LBWR(16'h0306);
TASK_LBWR(16'h0307);
TASK_LBWR(16'h0308);
TASK_LBWR(16'h0309);
TASK_LBWR(16'h030A);
TASK_LBWR(16'h030B);
TASK_LBWR(16'h030C);
TASK_LBWR(16'h030D);
TASK_LBWR(16'h030E);
TASK_LBWR(16'h030F);
TASK_PP(16'h0000,4);
TASK_PP(16'h0001,4);
TASK_PP(16'h0002,4);
TASK_PP(16'h0003,4);
TASK_PP(16'h0004,4);
TASK_PP(16'h0005,4);
TASK_PP(16'h0006,4);
TASK_PP(16'h0007,4);
TASK_PP(16'h0008,4);
TASK_PP(16'h0009,4);
TASK_PP(16'h000A,4);
TASK_PP(16'h000B,4);
TASK_PP(16'h000C,4);
TASK_PP(16'h000D,4);
TASK_PP(16'h000E,4);
TASK_PP(16'h000F,4);
TASK_PP(16'h0010,4);
TASK_PP(16'h0011,4);
TASK_PP(16'h0012,4);
TASK_PP(16'h0013,4);
TASK_PP(16'h0014,4);
TASK_PP(16'h0015,4);
TASK_PP(16'h0016,4);
TASK_PP(16'h0017,4);
TASK_PP(16'h0018,4);
TASK_PP(16'h0019,4);
TASK_PP(16'h001A,4);
TASK_PP(16'h001B,4);
TASK_PP(16'h001C,4);
TASK_PP(16'h001D,4);
TASK_PP(16'h001E,4);
TASK_PP(16'h001F,4);
TASK_PP(16'h0020,4);
TASK_PP(16'h0021,4);
TASK_PP(16'h0022,4);
TASK_PP(16'h0023,4);
TASK_PP(16'h0024,4);
TASK_PP(16'h0025,4);
TASK_PP(16'h0026,4);
TASK_PP(16'h0027,4);
TASK_PP(16'h0028,4);
TASK_PP(16'h0029,4);
TASK_PP(16'h002A,4);
TASK_PP(16'h002B,4);
TASK_PP(16'h002C,4);
TASK_PP(16'h002D,4);
TASK_PP(16'h002E,4);
TASK_PP(16'h002F,4);
TASK_PP(16'h0030,4);
TASK_PP(16'h0031,4);
TASK_PP(16'h0032,4);
TASK_PP(16'h0033,4);
TASK_PP(16'h0034,4);
TASK_PP(16'h0035,4);
TASK_PP(16'h0036,4);
TASK_PP(16'h0037,4);
TASK_PP(16'h0038,4);
TASK_PP(16'h0039,4);
TASK_PP(16'h003A,4);
TASK_PP(16'h003B,4);
TASK_PP(16'h003C,4);
TASK_PP(16'h003D,4);
TASK_PP(16'h003E,4);
TASK_PP(16'h003F,4);
TASK_PP(16'h0040,4);
TASK_PP(16'h0041,4);
TASK_PP(16'h0042,4);
TASK_PP(16'h0043,4);
TASK_PP(16'h0044,4);
TASK_PP(16'h0045,4);
TASK_PP(16'h0046,4);
TASK_PP(16'h0047,4);
TASK_PP(16'h0048,4);
TASK_PP(16'h0049,4);
TASK_PP(16'h004A,4);
TASK_PP(16'h004B,4);
TASK_PP(16'h004C,4);
TASK_PP(16'h004D,4);
TASK_PP(16'h004E,4);
TASK_PP(16'h004F,4);
TASK_PP(16'h0050,4);
TASK_PP(16'h0051,4);
TASK_PP(16'h0052,4);
TASK_PP(16'h0053,4);
TASK_PP(16'h0054,4);
TASK_PP(16'h0055,4);
TASK_PP(16'h0056,4);
TASK_PP(16'h0057,4);
TASK_PP(16'h0058,4);
TASK_PP(16'h0059,4);
TASK_PP(16'h005A,4);
TASK_PP(16'h005B,4);
TASK_PP(16'h005C,4);
TASK_PP(16'h005D,4);
TASK_PP(16'h005E,4);
TASK_PP(16'h005F,4);
TASK_PP(16'h0060,4);
TASK_PP(16'h0061,4);
TASK_PP(16'h0062,4);
TASK_PP(16'h0063,4);
TASK_PP(16'h0064,4);
TASK_PP(16'h0065,4);
TASK_PP(16'h0066,4);
TASK_PP(16'h0067,4);
TASK_PP(16'h0068,4);
TASK_PP(16'h0069,4);
TASK_PP(16'h006A,4);
TASK_PP(16'h006B,4);
TASK_PP(16'h006C,4);
TASK_PP(16'h006D,4);
TASK_PP(16'h006E,4);
TASK_PP(16'h006F,4);
TASK_PP(16'h0070,4);
TASK_PP(16'h0071,4);
TASK_PP(16'h0072,4);
TASK_PP(16'h0073,4);
TASK_PP(16'h0074,4);
TASK_PP(16'h0075,4);
TASK_PP(16'h0076,4);
TASK_PP(16'h0077,4);
TASK_PP(16'h0078,4);
TASK_PP(16'h0079,4);
TASK_PP(16'h007A,4);
TASK_PP(16'h007B,4);
TASK_PP(16'h007C,4);
TASK_PP(16'h007D,4);
TASK_PP(16'h007E,4);
TASK_PP(16'h007F,4);
TASK_PP(16'h0080,4);
TASK_PP(16'h0081,4);
TASK_PP(16'h0082,4);
TASK_PP(16'h0083,4);
TASK_PP(16'h0084,4);
TASK_PP(16'h0085,4);
TASK_PP(16'h0086,4);
TASK_PP(16'h0087,4);
TASK_PP(16'h0088,4);
TASK_PP(16'h0089,4);
TASK_PP(16'h008A,4);
TASK_PP(16'h008B,4);
TASK_PP(16'h008C,4);
TASK_PP(16'h008D,4);
TASK_PP(16'h008E,4);
TASK_PP(16'h008F,4);
TASK_PP(16'h0090,4);
TASK_PP(16'h0091,4);
TASK_PP(16'h0092,4);
TASK_PP(16'h0093,4);
TASK_PP(16'h0094,4);
TASK_PP(16'h0095,4);
TASK_PP(16'h0096,4);
TASK_PP(16'h0097,4);
TASK_PP(16'h0098,4);
TASK_PP(16'h0099,4);
TASK_PP(16'h009A,4);
TASK_PP(16'h009B,4);
TASK_PP(16'h009C,4);
TASK_PP(16'h009D,4);
TASK_PP(16'h009E,4);
TASK_PP(16'h009F,4);
TASK_PP(16'h00A0,4);
TASK_PP(16'h00A1,4);
TASK_PP(16'h00A2,4);
TASK_PP(16'h00A3,4);
TASK_PP(16'h00A4,4);
TASK_PP(16'h00A5,4);
TASK_PP(16'h00A6,4);
TASK_PP(16'h00A7,4);
TASK_PP(16'h00A8,4);
TASK_PP(16'h00A9,4);
TASK_PP(16'h00AA,4);
TASK_PP(16'h00AB,4);
TASK_PP(16'h00AC,4);
TASK_PP(16'h00AD,4);
TASK_PP(16'h00AE,4);
TASK_PP(16'h00AF,4);
TASK_PP(16'h00B0,4);
TASK_PP(16'h00B1,4);
TASK_PP(16'h00B2,4);
TASK_PP(16'h00B3,4);
TASK_PP(16'h00B4,4);
TASK_PP(16'h00B5,4);
TASK_PP(16'h00B6,4);
TASK_PP(16'h00B7,4);
TASK_PP(16'h00B8,4);
TASK_PP(16'h00B9,4);
TASK_PP(16'h00BA,4);
TASK_PP(16'h00BB,4);
TASK_PP(16'h00BC,4);
TASK_PP(16'h00BD,4);
TASK_PP(16'h00BE,4);
TASK_PP(16'h00BF,4);
TASK_PP(16'h00C0,4);
TASK_PP(16'h00C1,4);
TASK_PP(16'h00C2,4);
TASK_PP(16'h00C3,4);
TASK_PP(16'h00C4,4);
TASK_PP(16'h00C5,4);
TASK_PP(16'h00C6,4);
TASK_PP(16'h00C7,4);
TASK_PP(16'h00C8,4);
TASK_PP(16'h00C9,4);
TASK_PP(16'h00CA,4);
TASK_PP(16'h00CB,4);
TASK_PP(16'h00CC,4);
TASK_PP(16'h00CD,4);
TASK_PP(16'h00CE,4);
TASK_PP(16'h00CF,4);
TASK_PP(16'h00D0,4);
TASK_PP(16'h00D1,4);
TASK_PP(16'h00D2,4);
TASK_PP(16'h00D3,4);
TASK_PP(16'h00D4,4);
TASK_PP(16'h00D5,4);
TASK_PP(16'h00D6,4);
TASK_PP(16'h00D7,4);
TASK_PP(16'h00D8,4);
TASK_PP(16'h00D9,4);
TASK_PP(16'h00DA,4);
TASK_PP(16'h00DB,4);
TASK_PP(16'h00DC,4);
TASK_PP(16'h00DD,4);
TASK_PP(16'h00DE,4);
TASK_PP(16'h00DF,4);
TASK_PP(16'h00E0,4);
TASK_PP(16'h00E1,4);
TASK_PP(16'h00E2,4);
TASK_PP(16'h00E3,4);
TASK_PP(16'h00E4,4);
TASK_PP(16'h00E5,4);
TASK_PP(16'h00E6,4);
TASK_PP(16'h00E7,4);
TASK_PP(16'h00E8,4);
TASK_PP(16'h00E9,4);
TASK_PP(16'h00EA,4);
TASK_PP(16'h00EB,4);
TASK_PP(16'h00EC,4);
TASK_PP(16'h00ED,4);
TASK_PP(16'h00EE,4);
TASK_PP(16'h00EF,4);
TASK_PP(16'h00F0,4);
TASK_PP(16'h00F1,4);
TASK_PP(16'h00F2,4);
TASK_PP(16'h00F3,4);
TASK_PP(16'h00F4,4);
TASK_PP(16'h00F5,4);
TASK_PP(16'h00F6,4);
TASK_PP(16'h00F7,4);
TASK_PP(16'h00F8,4);
TASK_PP(16'h00F9,4);
TASK_PP(16'h00FA,4);
TASK_PP(16'h00FB,4);
TASK_PP(16'h00FC,4);
TASK_PP(16'h00FD,4);
TASK_PP(16'h00FE,4);
TASK_PP(16'h00FF,4);
TASK_PP(16'h0100,4);
TASK_PP(16'h0101,4);
TASK_PP(16'h0102,4);
TASK_PP(16'h0103,4);
TASK_PP(16'h0104,4);
TASK_PP(16'h0105,4);
TASK_PP(16'h0106,4);
TASK_PP(16'h0107,4);
TASK_PP(16'h0108,4);
TASK_PP(16'h0109,4);
TASK_PP(16'h010A,4);
TASK_PP(16'h010B,4);
TASK_PP(16'h010C,4);
TASK_PP(16'h010D,4);
TASK_PP(16'h010E,4);
TASK_PP(16'h010F,4);
TASK_PP(16'h0110,4);
TASK_PP(16'h0111,4);
TASK_PP(16'h0112,4);
TASK_PP(16'h0113,4);
TASK_PP(16'h0114,4);
TASK_PP(16'h0115,4);
TASK_PP(16'h0116,4);
TASK_PP(16'h0117,4);
TASK_PP(16'h0118,4);
TASK_PP(16'h0119,4);
TASK_PP(16'h011A,4);
TASK_PP(16'h011B,4);
TASK_PP(16'h011C,4);
TASK_PP(16'h011D,4);
TASK_PP(16'h011E,4);
TASK_PP(16'h011F,4);
TASK_PP(16'h0120,4);
TASK_PP(16'h0121,4);
TASK_PP(16'h0122,4);
TASK_PP(16'h0123,4);
TASK_PP(16'h0124,4);
TASK_PP(16'h0125,4);
TASK_PP(16'h0126,4);
TASK_PP(16'h0127,4);
TASK_PP(16'h0128,4);
TASK_PP(16'h0129,4);
TASK_PP(16'h012A,4);
TASK_PP(16'h012B,4);
TASK_PP(16'h012C,4);
TASK_PP(16'h012D,4);
TASK_PP(16'h012E,4);
TASK_PP(16'h012F,4);
TASK_PP(16'h0130,4);
TASK_PP(16'h0131,4);
TASK_PP(16'h0132,4);
TASK_PP(16'h0133,4);
TASK_PP(16'h0134,4);
TASK_PP(16'h0135,4);
TASK_PP(16'h0136,4);
TASK_PP(16'h0137,4);
TASK_PP(16'h0138,4);
TASK_PP(16'h0139,4);
TASK_PP(16'h013A,4);
TASK_PP(16'h013B,4);
TASK_PP(16'h013C,4);
TASK_PP(16'h013D,4);
TASK_PP(16'h013E,4);
TASK_PP(16'h013F,4);
TASK_PP(16'h0140,4);
TASK_PP(16'h0141,4);
TASK_PP(16'h0142,4);
TASK_PP(16'h0143,4);
TASK_PP(16'h0144,4);
TASK_PP(16'h0145,4);
TASK_PP(16'h0146,4);
TASK_PP(16'h0147,4);
TASK_PP(16'h0148,4);
TASK_PP(16'h0149,4);
TASK_PP(16'h014A,4);
TASK_PP(16'h014B,4);
TASK_PP(16'h014C,4);
TASK_PP(16'h014D,4);
TASK_PP(16'h014E,4);
TASK_PP(16'h014F,4);
TASK_PP(16'h0150,4);
TASK_PP(16'h0151,4);
TASK_PP(16'h0152,4);
TASK_PP(16'h0153,4);
TASK_PP(16'h0154,4);
TASK_PP(16'h0155,4);
TASK_PP(16'h0156,4);
TASK_PP(16'h0157,4);
TASK_PP(16'h0158,4);
TASK_PP(16'h0159,4);
TASK_PP(16'h015A,4);
TASK_PP(16'h015B,4);
TASK_PP(16'h015C,4);
TASK_PP(16'h015D,4);
TASK_PP(16'h015E,4);
TASK_PP(16'h015F,4);
TASK_PP(16'h0160,4);
TASK_PP(16'h0161,4);
TASK_PP(16'h0162,4);
TASK_PP(16'h0163,4);
TASK_PP(16'h0164,4);
TASK_PP(16'h0165,4);
TASK_PP(16'h0166,4);
TASK_PP(16'h0167,4);
TASK_PP(16'h0168,4);
TASK_PP(16'h0169,4);
TASK_PP(16'h016A,4);
TASK_PP(16'h016B,4);
TASK_PP(16'h016C,4);
TASK_PP(16'h016D,4);
TASK_PP(16'h016E,4);
TASK_PP(16'h016F,4);
TASK_PP(16'h0170,4);
TASK_PP(16'h0171,4);
TASK_PP(16'h0172,4);
TASK_PP(16'h0173,4);
TASK_PP(16'h0174,4);
TASK_PP(16'h0175,4);
TASK_PP(16'h0176,4);
TASK_PP(16'h0177,4);
TASK_PP(16'h0178,4);
TASK_PP(16'h0179,4);
TASK_PP(16'h017A,4);
TASK_PP(16'h017B,4);
TASK_PP(16'h017C,4);
TASK_PP(16'h017D,4);
TASK_PP(16'h017E,4);
TASK_PP(16'h017F,4);
TASK_PP(16'h0180,4);
TASK_PP(16'h0181,4);
TASK_PP(16'h0182,4);
TASK_PP(16'h0183,4);
TASK_PP(16'h0184,4);
TASK_PP(16'h0185,4);
TASK_PP(16'h0186,4);
TASK_PP(16'h0187,4);
TASK_PP(16'h0188,4);
TASK_PP(16'h0189,4);
TASK_PP(16'h018A,4);
TASK_PP(16'h018B,4);
TASK_PP(16'h018C,4);
TASK_PP(16'h018D,4);
TASK_PP(16'h018E,4);
TASK_PP(16'h018F,4);
TASK_PP(16'h0190,4);
TASK_PP(16'h0191,4);
TASK_PP(16'h0192,4);
TASK_PP(16'h0193,4);
TASK_PP(16'h0194,4);
TASK_PP(16'h0195,4);
TASK_PP(16'h0196,4);
TASK_PP(16'h0197,4);
TASK_PP(16'h0198,4);
TASK_PP(16'h0199,4);
TASK_PP(16'h019A,4);
TASK_PP(16'h019B,4);
TASK_PP(16'h019C,4);
TASK_PP(16'h019D,4);
TASK_PP(16'h019E,4);
TASK_PP(16'h019F,4);
TASK_PP(16'h01A0,4);
TASK_PP(16'h01A1,4);
TASK_PP(16'h01A2,4);
TASK_PP(16'h01A3,4);
TASK_PP(16'h01A4,4);
TASK_PP(16'h01A5,4);
TASK_PP(16'h01A6,4);
TASK_PP(16'h01A7,4);
TASK_PP(16'h01A8,4);
TASK_PP(16'h01A9,4);
TASK_PP(16'h01AA,4);
TASK_PP(16'h01AB,4);
TASK_PP(16'h01AC,4);
TASK_PP(16'h01AD,4);
TASK_PP(16'h01AE,4);
TASK_PP(16'h01AF,4);
TASK_PP(16'h01B0,4);
TASK_PP(16'h01B1,4);
TASK_PP(16'h01B2,4);
TASK_PP(16'h01B3,4);
TASK_PP(16'h01B4,4);
TASK_PP(16'h01B5,4);
TASK_PP(16'h01B6,4);
TASK_PP(16'h01B7,4);
TASK_PP(16'h01B8,4);
TASK_PP(16'h01B9,4);
TASK_PP(16'h01BA,4);
TASK_PP(16'h01BB,4);
TASK_PP(16'h01BC,4);
TASK_PP(16'h01BD,4);
TASK_PP(16'h01BE,4);
TASK_PP(16'h01BF,4);
TASK_PP(16'h01C0,4);
TASK_PP(16'h01C1,4);
TASK_PP(16'h01C2,4);
TASK_PP(16'h01C3,4);
TASK_PP(16'h01C4,4);
TASK_PP(16'h01C5,4);
TASK_PP(16'h01C6,4);
TASK_PP(16'h01C7,4);
TASK_PP(16'h01C8,4);
TASK_PP(16'h01C9,4);
TASK_PP(16'h01CA,4);
TASK_PP(16'h01CB,4);
TASK_PP(16'h01CC,4);
TASK_PP(16'h01CD,4);
TASK_PP(16'h01CE,4);
TASK_PP(16'h01CF,4);
TASK_PP(16'h01D0,4);
TASK_PP(16'h01D1,4);
TASK_PP(16'h01D2,4);
TASK_PP(16'h01D3,4);
TASK_PP(16'h01D4,4);
TASK_PP(16'h01D5,4);
TASK_PP(16'h01D6,4);
TASK_PP(16'h01D7,4);
TASK_PP(16'h01D8,4);
TASK_PP(16'h01D9,4);
TASK_PP(16'h01DA,4);
TASK_PP(16'h01DB,4);
TASK_PP(16'h01DC,4);
TASK_PP(16'h01DD,4);
TASK_PP(16'h01DE,4);
TASK_PP(16'h01DF,4);
TASK_PP(16'h01E0,4);
TASK_PP(16'h01E1,4);
TASK_PP(16'h01E2,4);
TASK_PP(16'h01E3,4);
TASK_PP(16'h01E4,4);
TASK_PP(16'h01E5,4);
TASK_PP(16'h01E6,4);
TASK_PP(16'h01E7,4);
TASK_PP(16'h01E8,4);
TASK_PP(16'h01E9,4);
TASK_PP(16'h01EA,4);
TASK_PP(16'h01EB,4);
TASK_PP(16'h01EC,4);
TASK_PP(16'h01ED,4);
TASK_PP(16'h01EE,4);
TASK_PP(16'h01EF,4);
TASK_PP(16'h01F0,4);
TASK_PP(16'h01F1,4);
TASK_PP(16'h01F2,4);
TASK_PP(16'h01F3,4);
TASK_PP(16'h01F4,4);
TASK_PP(16'h01F5,4);
TASK_PP(16'h01F6,4);
TASK_PP(16'h01F7,4);
TASK_PP(16'h01F8,4);
TASK_PP(16'h01F9,4);
TASK_PP(16'h01FA,4);
TASK_PP(16'h01FB,4);
TASK_PP(16'h01FC,4);
TASK_PP(16'h01FD,4);
TASK_PP(16'h01FE,4);
TASK_PP(16'h01FF,4);
TASK_PP(16'h0200,4);
TASK_PP(16'h0201,4);
TASK_PP(16'h0202,4);
TASK_PP(16'h0203,4);
TASK_PP(16'h0204,4);
TASK_PP(16'h0205,4);
TASK_PP(16'h0206,4);
TASK_PP(16'h0207,4);
TASK_PP(16'h0208,4);
TASK_PP(16'h0209,4);
TASK_PP(16'h020A,4);
TASK_PP(16'h020B,4);
TASK_PP(16'h020C,4);
TASK_PP(16'h020D,4);
TASK_PP(16'h020E,4);
TASK_PP(16'h020F,4);
TASK_PP(16'h0210,4);
TASK_PP(16'h0211,4);
TASK_PP(16'h0212,4);
TASK_PP(16'h0213,4);
TASK_PP(16'h0214,4);
TASK_PP(16'h0215,4);
TASK_PP(16'h0216,4);
TASK_PP(16'h0217,4);
TASK_PP(16'h0218,4);
TASK_PP(16'h0219,4);
TASK_PP(16'h021A,4);
TASK_PP(16'h021B,4);
TASK_PP(16'h021C,4);
TASK_PP(16'h021D,4);
TASK_PP(16'h021E,4);
TASK_PP(16'h021F,4);
TASK_PP(16'h0220,4);
TASK_PP(16'h0221,4);
TASK_PP(16'h0222,4);
TASK_PP(16'h0223,4);
TASK_PP(16'h0224,4);
TASK_PP(16'h0225,4);
TASK_PP(16'h0226,4);
TASK_PP(16'h0227,4);
TASK_PP(16'h0228,4);
TASK_PP(16'h0229,4);
TASK_PP(16'h022A,4);
TASK_PP(16'h022B,4);
TASK_PP(16'h022C,4);
TASK_PP(16'h022D,4);
TASK_PP(16'h022E,4);
TASK_PP(16'h022F,4);
TASK_PP(16'h0230,4);
TASK_PP(16'h0231,4);
TASK_PP(16'h0232,4);
TASK_PP(16'h0233,4);
TASK_PP(16'h0234,4);
TASK_PP(16'h0235,4);
TASK_PP(16'h0236,4);
TASK_PP(16'h0237,4);
TASK_PP(16'h0238,4);
TASK_PP(16'h0239,4);
TASK_PP(16'h023A,4);
TASK_PP(16'h023B,4);
TASK_PP(16'h023C,4);
TASK_PP(16'h023D,4);
TASK_PP(16'h023E,4);
TASK_PP(16'h023F,4);
TASK_PP(16'h0240,4);
TASK_PP(16'h0241,4);
TASK_PP(16'h0242,4);
TASK_PP(16'h0243,4);
TASK_PP(16'h0244,4);
TASK_PP(16'h0245,4);
TASK_PP(16'h0246,4);
TASK_PP(16'h0247,4);
TASK_PP(16'h0248,4);
TASK_PP(16'h0249,4);
TASK_PP(16'h024A,4);
TASK_PP(16'h024B,4);
TASK_PP(16'h024C,4);
TASK_PP(16'h024D,4);
TASK_PP(16'h024E,4);
TASK_PP(16'h024F,4);
TASK_PP(16'h0250,4);
TASK_PP(16'h0251,4);
TASK_PP(16'h0252,4);
TASK_PP(16'h0253,4);
TASK_PP(16'h0254,4);
TASK_PP(16'h0255,4);
TASK_PP(16'h0256,4);
TASK_PP(16'h0257,4);
TASK_PP(16'h0258,4);
TASK_PP(16'h0259,4);
TASK_PP(16'h025A,4);
TASK_PP(16'h025B,4);
TASK_PP(16'h025C,4);
TASK_PP(16'h025D,4);
TASK_PP(16'h025E,4);
TASK_PP(16'h025F,4);
TASK_PP(16'h0260,4);
TASK_PP(16'h0261,4);
TASK_PP(16'h0262,4);
TASK_PP(16'h0263,4);
TASK_PP(16'h0264,4);
TASK_PP(16'h0265,4);
TASK_PP(16'h0266,4);
TASK_PP(16'h0267,4);
TASK_PP(16'h0268,4);
TASK_PP(16'h0269,4);
TASK_PP(16'h026A,4);
TASK_PP(16'h026B,4);
TASK_PP(16'h026C,4);
TASK_PP(16'h026D,4);
TASK_PP(16'h026E,4);
TASK_PP(16'h026F,4);
TASK_PP(16'h0270,4);
TASK_PP(16'h0271,4);
TASK_PP(16'h0272,4);
TASK_PP(16'h0273,4);
TASK_PP(16'h0274,4);
TASK_PP(16'h0275,4);
TASK_PP(16'h0276,4);
TASK_PP(16'h0277,4);
TASK_PP(16'h0278,4);
TASK_PP(16'h0279,4);
TASK_PP(16'h027A,4);
TASK_PP(16'h027B,4);
TASK_PP(16'h027C,4);
TASK_PP(16'h027D,4);
TASK_PP(16'h027E,4);
TASK_PP(16'h027F,4);
TASK_PP(16'h0280,4);
TASK_PP(16'h0281,4);
TASK_PP(16'h0282,4);
TASK_PP(16'h0283,4);
TASK_PP(16'h0284,4);
TASK_PP(16'h0285,4);
TASK_PP(16'h0286,4);
TASK_PP(16'h0287,4);
TASK_PP(16'h0288,4);
TASK_PP(16'h0289,4);
TASK_PP(16'h028A,4);
TASK_PP(16'h028B,4);
TASK_PP(16'h028C,4);
TASK_PP(16'h028D,4);
TASK_PP(16'h028E,4);
TASK_PP(16'h028F,4);
TASK_PP(16'h0290,4);
TASK_PP(16'h0291,4);
TASK_PP(16'h0292,4);
TASK_PP(16'h0293,4);
TASK_PP(16'h0294,4);
TASK_PP(16'h0295,4);
TASK_PP(16'h0296,4);
TASK_PP(16'h0297,4);
TASK_PP(16'h0298,4);
TASK_PP(16'h0299,4);
TASK_PP(16'h029A,4);
TASK_PP(16'h029B,4);
TASK_PP(16'h029C,4);
TASK_PP(16'h029D,4);
TASK_PP(16'h029E,4);
TASK_PP(16'h029F,4);
TASK_PP(16'h02A0,4);
TASK_PP(16'h02A1,4);
TASK_PP(16'h02A2,4);
TASK_PP(16'h02A3,4);
TASK_PP(16'h02A4,4);
TASK_PP(16'h02A5,4);
TASK_PP(16'h02A6,4);
TASK_PP(16'h02A7,4);
TASK_PP(16'h02A8,4);
TASK_PP(16'h02A9,4);
TASK_PP(16'h02AA,4);
TASK_PP(16'h02AB,4);
TASK_PP(16'h02AC,4);
TASK_PP(16'h02AD,4);
TASK_PP(16'h02AE,4);
TASK_PP(16'h02AF,4);
TASK_PP(16'h02B0,4);
TASK_PP(16'h02B1,4);
TASK_PP(16'h02B2,4);
TASK_PP(16'h02B3,4);
TASK_PP(16'h02B4,4);
TASK_PP(16'h02B5,4);
TASK_PP(16'h02B6,4);
TASK_PP(16'h02B7,4);
TASK_PP(16'h02B8,4);
TASK_PP(16'h02B9,4);
TASK_PP(16'h02BA,4);
TASK_PP(16'h02BB,4);
TASK_PP(16'h02BC,4);
TASK_PP(16'h02BD,4);
TASK_PP(16'h02BE,4);
TASK_PP(16'h02BF,4);
TASK_PP(16'h02C0,4);
TASK_PP(16'h02C1,4);
TASK_PP(16'h02C2,4);
TASK_PP(16'h02C3,4);
TASK_PP(16'h02C4,4);
TASK_PP(16'h02C5,4);
TASK_PP(16'h02C6,4);
TASK_PP(16'h02C7,4);
TASK_PP(16'h02C8,4);
TASK_PP(16'h02C9,4);
TASK_PP(16'h02CA,4);
TASK_PP(16'h02CB,4);
TASK_PP(16'h02CC,4);
TASK_PP(16'h02CD,4);
TASK_PP(16'h02CE,4);
TASK_PP(16'h02CF,4);
TASK_PP(16'h02D0,4);
TASK_PP(16'h02D1,4);
TASK_PP(16'h02D2,4);
TASK_PP(16'h02D3,4);
TASK_PP(16'h02D4,4);
TASK_PP(16'h02D5,4);
TASK_PP(16'h02D6,4);
TASK_PP(16'h02D7,4);
TASK_PP(16'h02D8,4);
TASK_PP(16'h02D9,4);
TASK_PP(16'h02DA,4);
TASK_PP(16'h02DB,4);
TASK_PP(16'h02DC,4);
TASK_PP(16'h02DD,4);
TASK_PP(16'h02DE,4);
TASK_PP(16'h02DF,4);
TASK_PP(16'h02E0,4);
TASK_PP(16'h02E1,4);
TASK_PP(16'h02E2,4);
TASK_PP(16'h02E3,4);
TASK_PP(16'h02E4,4);
TASK_PP(16'h02E5,4);
TASK_PP(16'h02E6,4);
TASK_PP(16'h02E7,4);
TASK_PP(16'h02E8,4);
TASK_PP(16'h02E9,4);
TASK_PP(16'h02EA,4);
TASK_PP(16'h02EB,4);
TASK_PP(16'h02EC,4);
TASK_PP(16'h02ED,4);
TASK_PP(16'h02EE,4);
TASK_PP(16'h02EF,4);
TASK_PP(16'h02F0,4);
TASK_PP(16'h02F1,4);
TASK_PP(16'h02F2,4);
TASK_PP(16'h02F3,4);
TASK_PP(16'h02F4,4);
TASK_PP(16'h02F5,4);
TASK_PP(16'h02F6,4);
TASK_PP(16'h02F7,4);
TASK_PP(16'h02F8,4);
TASK_PP(16'h02F9,4);
TASK_PP(16'h02FA,4);
TASK_PP(16'h02FB,4);
TASK_PP(16'h02FC,4);
TASK_PP(16'h02FD,4);
TASK_PP(16'h02FE,4);
TASK_PP(16'h02FF,4);
TASK_PP(16'h0300,4);
TASK_PP(16'h0301,4);
TASK_PP(16'h0302,4);
TASK_PP(16'h0303,4);
TASK_PP(16'h0304,4);
TASK_PP(16'h0305,4);
TASK_PP(16'h0306,4);
TASK_PP(16'h0307,4);
TASK_PP(16'h0308,4);
TASK_PP(16'h0309,4);
TASK_PP(16'h030A,4);
TASK_PP(16'h030B,4);
TASK_PP(16'h030C,4);
TASK_PP(16'h030D,4);
TASK_PP(16'h030E,4);
TASK_PP(16'h030F,4);
TASK_PP(16'h0310,4);
TASK_PP(16'h0311,4);
TASK_PP(16'h0312,4);
TASK_PP(16'h0313,4);
TASK_PP(16'h0314,4);
TASK_PP(16'h0315,4);
TASK_PP(16'h0316,4);
TASK_PP(16'h0317,4);
TASK_PP(16'h0318,4);
TASK_PP(16'h0319,4);
TASK_PP(16'h031A,4);
TASK_PP(16'h031B,4);
TASK_PP(16'h031C,4);
TASK_PP(16'h031D,4);
TASK_PP(16'h031E,4);
TASK_PP(16'h031F,4);
TASK_PP(16'h0320,4);
TASK_PP(16'h0321,4);
TASK_PP(16'h0322,4);
TASK_PP(16'h0323,4);
TASK_PP(16'h0324,4);
TASK_PP(16'h0325,4);
TASK_PP(16'h0326,4);
TASK_PP(16'h0327,4);
TASK_PP(16'h0328,4);
TASK_PP(16'h0329,4);
TASK_PP(16'h032A,4);
TASK_PP(16'h032B,4);
TASK_PP(16'h032C,4);
TASK_PP(16'h032D,4);
TASK_PP(16'h032E,4);
TASK_PP(16'h032F,4);
TASK_PP(16'h0330,4);
TASK_PP(16'h0331,4);
TASK_PP(16'h0332,4);
TASK_PP(16'h0333,4);
TASK_PP(16'h0334,4);
TASK_PP(16'h0335,4);
TASK_PP(16'h0336,4);
TASK_PP(16'h0337,4);
TASK_PP(16'h0338,4);
TASK_PP(16'h0339,4);
TASK_PP(16'h033A,4);
TASK_PP(16'h033B,4);
TASK_PP(16'h033C,4);
TASK_PP(16'h033D,4);
TASK_PP(16'h033E,4);
TASK_PP(16'h033F,4);
TASK_PP(16'h0340,4);
TASK_PP(16'h0341,4);
TASK_PP(16'h0342,4);
TASK_PP(16'h0343,4);
TASK_PP(16'h0344,4);
TASK_PP(16'h0345,4);
TASK_PP(16'h0346,4);
TASK_PP(16'h0347,4);
TASK_PP(16'h0348,4);
TASK_PP(16'h0349,4);
TASK_PP(16'h034A,4);
TASK_PP(16'h034B,4);
TASK_PP(16'h034C,4);
TASK_PP(16'h034D,4);
TASK_PP(16'h034E,4);
TASK_PP(16'h034F,4);
TASK_PP(16'h0350,4);
TASK_PP(16'h0351,4);
TASK_PP(16'h0352,4);
TASK_PP(16'h0353,4);
TASK_PP(16'h0354,4);
TASK_PP(16'h0355,4);
TASK_PP(16'h0356,4);
TASK_PP(16'h0357,4);
TASK_PP(16'h0358,4);
TASK_PP(16'h0359,4);
TASK_PP(16'h035A,4);
TASK_PP(16'h035B,4);
TASK_PP(16'h035C,4);
TASK_PP(16'h035D,4);
TASK_PP(16'h035E,4);
TASK_PP(16'h035F,4);
TASK_PP(16'h0360,4);
TASK_PP(16'h0361,4);
TASK_PP(16'h0362,4);
TASK_PP(16'h0363,4);
TASK_PP(16'h0364,4);
TASK_PP(16'h0365,4);
TASK_PP(16'h0366,4);
TASK_PP(16'h0367,4);
TASK_PP(16'h0368,4);
TASK_PP(16'h0369,4);
TASK_PP(16'h036A,4);
TASK_PP(16'h036B,4);
TASK_PP(16'h036C,4);
TASK_PP(16'h036D,4);
TASK_PP(16'h036E,4);
TASK_PP(16'h036F,4);
TASK_PP(16'h0370,4);
TASK_PP(16'h0371,4);
TASK_PP(16'h0372,4);
TASK_PP(16'h0373,4);
TASK_PP(16'h0374,4);
TASK_PP(16'h0375,4);
TASK_PP(16'h0376,4);
TASK_PP(16'h0377,4);
TASK_PP(16'h0378,4);
TASK_PP(16'h0379,4);
TASK_PP(16'h037A,4);
TASK_PP(16'h037B,4);
TASK_PP(16'h037C,4);
TASK_PP(16'h037D,4);
TASK_PP(16'h037E,4);
TASK_PP(16'h037F,4);
TASK_PP(16'h0380,4);
TASK_PP(16'h0381,4);
TASK_PP(16'h0382,4);
TASK_PP(16'h0383,4);
TASK_PP(16'h0384,4);
TASK_PP(16'h0385,4);
TASK_PP(16'h0386,4);
TASK_PP(16'h0387,4);
TASK_PP(16'h0388,4);
TASK_PP(16'h0389,4);
TASK_PP(16'h038A,4);
TASK_PP(16'h038B,4);
TASK_PP(16'h038C,4);
TASK_PP(16'h038D,4);
TASK_PP(16'h038E,4);
TASK_PP(16'h038F,4);
TASK_PP(16'h0390,4);
TASK_PP(16'h0391,4);
TASK_PP(16'h0392,4);
TASK_PP(16'h0393,4);
TASK_PP(16'h0394,4);
TASK_PP(16'h0395,4);
TASK_PP(16'h0396,4);
TASK_PP(16'h0397,4);
TASK_PP(16'h0398,4);
TASK_PP(16'h0399,4);
TASK_PP(16'h039A,4);
TASK_PP(16'h039B,4);
TASK_PP(16'h039C,4);
TASK_PP(16'h039D,4);
TASK_PP(16'h039E,4);
TASK_PP(16'h039F,4);
TASK_PP(16'h03A0,4);
TASK_PP(16'h03A1,4);
TASK_PP(16'h03A2,4);
TASK_PP(16'h03A3,4);
TASK_PP(16'h03A4,4);
TASK_PP(16'h03A5,4);
TASK_PP(16'h03A6,4);
TASK_PP(16'h03A7,4);
TASK_PP(16'h03A8,4);
TASK_PP(16'h03A9,4);
TASK_PP(16'h03AA,4);
TASK_PP(16'h03AB,4);
TASK_PP(16'h03AC,4);
TASK_PP(16'h03AD,4);
TASK_PP(16'h03AE,4);
TASK_PP(16'h03AF,4);
TASK_PP(16'h03B0,4);
TASK_PP(16'h03B1,4);
TASK_PP(16'h03B2,4);
TASK_PP(16'h03B3,4);
TASK_PP(16'h03B4,4);
TASK_PP(16'h03B5,4);
TASK_PP(16'h03B6,4);
TASK_PP(16'h03B7,4);
TASK_PP(16'h03B8,4);
TASK_PP(16'h03B9,4);
TASK_PP(16'h03BA,4);
TASK_PP(16'h03BB,4);
TASK_PP(16'h03BC,4);
TASK_PP(16'h03BD,4);
TASK_PP(16'h03BE,4);
TASK_PP(16'h03BF,4);
TASK_PP(16'h03C0,4);
TASK_PP(16'h03C1,4);
TASK_PP(16'h03C2,4);
TASK_PP(16'h03C3,4);
TASK_PP(16'h03C4,4);
TASK_PP(16'h03C5,4);
TASK_PP(16'h03C6,4);
TASK_PP(16'h03C7,4);
TASK_PP(16'h03C8,4);
TASK_PP(16'h03C9,4);
TASK_PP(16'h03CA,4);
TASK_PP(16'h03CB,4);
TASK_PP(16'h03CC,4);
TASK_PP(16'h03CD,4);
TASK_PP(16'h03CE,4);
TASK_PP(16'h03CF,4);
TASK_PP(16'h03D0,4);
TASK_PP(16'h03D1,4);
TASK_PP(16'h03D2,4);
TASK_PP(16'h03D3,4);
TASK_PP(16'h03D4,4);
TASK_PP(16'h03D5,4);
TASK_PP(16'h03D6,4);
TASK_PP(16'h03D7,4);
TASK_PP(16'h03D8,4);
TASK_PP(16'h03D9,4);
TASK_PP(16'h03DA,4);
TASK_PP(16'h03DB,4);
TASK_PP(16'h03DC,4);
TASK_PP(16'h03DD,4);
TASK_PP(16'h03DE,4);
TASK_PP(16'h03DF,4);
TASK_PP(16'h03E0,4);
TASK_PP(16'h03E1,4);
TASK_PP(16'h03E2,4);
TASK_PP(16'h03E3,4);
TASK_PP(16'h03E4,4);
TASK_PP(16'h03E5,4);
TASK_PP(16'h03E6,4);
TASK_PP(16'h03E7,4);
TASK_PP(16'h03E8,4);
TASK_PP(16'h03E9,4);
TASK_PP(16'h03EA,4);
TASK_PP(16'h03EB,4);
TASK_PP(16'h03EC,4);
TASK_PP(16'h03ED,4);
TASK_PP(16'h03EE,4);
TASK_PP(16'h03EF,4);
TASK_PP(16'h03F0,4);
TASK_PP(16'h03F1,4);
TASK_PP(16'h03F2,4);
TASK_PP(16'h03F3,4);
TASK_PP(16'h03F4,4);
TASK_PP(16'h03F5,4);
TASK_PP(16'h03F6,4);
TASK_PP(16'h03F7,4);
TASK_PP(16'h03F8,4);
TASK_PP(16'h03F9,4);
TASK_PP(16'h03FA,4);
TASK_PP(16'h03FB,4);
TASK_PP(16'h03FC,4);
TASK_PP(16'h03FD,4);
TASK_PP(16'h03FE,4);
TASK_PP(16'h03FF,4);
TASK_PP(16'h0400,4);
TASK_PP(16'h0401,4);
TASK_PP(16'h0402,4);
TASK_PP(16'h0403,4);
TASK_PP(16'h0404,4);
TASK_PP(16'h0405,4);
TASK_PP(16'h0406,4);
TASK_PP(16'h0407,4);
TASK_PP(16'h0408,4);
TASK_PP(16'h0409,4);
TASK_PP(16'h040A,4);
TASK_PP(16'h040B,4);
TASK_PP(16'h040C,4);
TASK_PP(16'h040D,4);
TASK_PP(16'h040E,4);
TASK_PP(16'h040F,4);
TASK_PP(16'h0410,4);
TASK_PP(16'h0411,4);
TASK_PP(16'h0412,4);
TASK_PP(16'h0413,4);
TASK_PP(16'h0414,4);
TASK_PP(16'h0415,4);
TASK_PP(16'h0416,4);
TASK_PP(16'h0417,4);
TASK_PP(16'h0418,4);
TASK_PP(16'h0419,4);
TASK_PP(16'h041A,4);
TASK_PP(16'h041B,4);
TASK_PP(16'h041C,4);
TASK_PP(16'h041D,4);
TASK_PP(16'h041E,4);
TASK_PP(16'h041F,4);
TASK_PP(16'h0420,4);
TASK_PP(16'h0421,4);
TASK_PP(16'h0422,4);
TASK_PP(16'h0423,4);
TASK_PP(16'h0424,4);
TASK_PP(16'h0425,4);
TASK_PP(16'h0426,4);
TASK_PP(16'h0427,4);
TASK_PP(16'h0428,4);
TASK_PP(16'h0429,4);
TASK_PP(16'h042A,4);
TASK_PP(16'h042B,4);
TASK_PP(16'h042C,4);
TASK_PP(16'h042D,4);
TASK_PP(16'h042E,4);
TASK_PP(16'h042F,4);
TASK_PP(16'h0430,4);
TASK_PP(16'h0431,4);
TASK_PP(16'h0432,4);
TASK_PP(16'h0433,4);
TASK_PP(16'h0434,4);
TASK_PP(16'h0435,4);
TASK_PP(16'h0436,4);
TASK_PP(16'h0437,4);
TASK_PP(16'h0438,4);
TASK_PP(16'h0439,4);
TASK_PP(16'h043A,4);
TASK_PP(16'h043B,4);
TASK_PP(16'h043C,4);
TASK_PP(16'h043D,4);
TASK_PP(16'h043E,4);
TASK_PP(16'h043F,4);
TASK_PP(16'h0440,4);
TASK_PP(16'h0441,4);
TASK_PP(16'h0442,4);
TASK_PP(16'h0443,4);
TASK_PP(16'h0444,4);
TASK_PP(16'h0445,4);
TASK_PP(16'h0446,4);
TASK_PP(16'h0447,4);
TASK_PP(16'h0448,4);
TASK_PP(16'h0449,4);
TASK_PP(16'h044A,4);
TASK_PP(16'h044B,4);
TASK_PP(16'h044C,4);
TASK_PP(16'h044D,4);
TASK_PP(16'h044E,4);
TASK_PP(16'h044F,4);
TASK_PP(16'h0450,4);
TASK_PP(16'h0451,4);
TASK_PP(16'h0452,4);
TASK_PP(16'h0453,4);
TASK_PP(16'h0454,4);
TASK_PP(16'h0455,4);
TASK_PP(16'h0456,4);
TASK_PP(16'h0457,4);
TASK_PP(16'h0458,4);
TASK_PP(16'h0459,4);
TASK_PP(16'h045A,4);
TASK_PP(16'h045B,4);
TASK_PP(16'h045C,4);
TASK_PP(16'h045D,4);
TASK_PP(16'h045E,4);
TASK_PP(16'h045F,4);
TASK_PP(16'h0460,4);
TASK_PP(16'h0461,4);
TASK_PP(16'h0462,4);
TASK_PP(16'h0463,4);
TASK_PP(16'h0464,4);
TASK_PP(16'h0465,4);
TASK_PP(16'h0466,4);
TASK_PP(16'h0467,4);
TASK_PP(16'h0468,4);
TASK_PP(16'h0469,4);
TASK_PP(16'h046A,4);
TASK_PP(16'h046B,4);
TASK_PP(16'h046C,4);
TASK_PP(16'h046D,4);
TASK_PP(16'h046E,4);
TASK_PP(16'h046F,4);
TASK_PP(16'h0470,4);
TASK_PP(16'h0471,4);
TASK_PP(16'h0472,4);
TASK_PP(16'h0473,4);
TASK_PP(16'h0474,4);
TASK_PP(16'h0475,4);
TASK_PP(16'h0476,4);
TASK_PP(16'h0477,4);
TASK_PP(16'h0478,4);
TASK_PP(16'h0479,4);
TASK_PP(16'h047A,4);
TASK_PP(16'h047B,4);
TASK_PP(16'h047C,4);
TASK_PP(16'h047D,4);
TASK_PP(16'h047E,4);
TASK_PP(16'h047F,4);
TASK_PP(16'h0480,4);
TASK_PP(16'h0481,4);
TASK_PP(16'h0482,4);
TASK_PP(16'h0483,4);
TASK_PP(16'h0484,4);
TASK_PP(16'h0485,4);
TASK_PP(16'h0486,4);
TASK_PP(16'h0487,4);
TASK_PP(16'h0488,4);
TASK_PP(16'h0489,4);
TASK_PP(16'h048A,4);
TASK_PP(16'h048B,4);
TASK_PP(16'h048C,4);
TASK_PP(16'h048D,4);
TASK_PP(16'h048E,4);
TASK_PP(16'h048F,4);
TASK_PP(16'h0490,4);
TASK_PP(16'h0491,4);
TASK_PP(16'h0492,4);
TASK_PP(16'h0493,4);
TASK_PP(16'h0494,4);
TASK_PP(16'h0495,4);
TASK_PP(16'h0496,4);
TASK_PP(16'h0497,4);
TASK_PP(16'h0498,4);
TASK_PP(16'h0499,4);
TASK_PP(16'h049A,4);
TASK_PP(16'h049B,4);
TASK_PP(16'h049C,4);
TASK_PP(16'h049D,4);
TASK_PP(16'h049E,4);
TASK_PP(16'h049F,4);
TASK_PP(16'h04A0,4);
TASK_PP(16'h04A1,4);
TASK_PP(16'h04A2,4);
TASK_PP(16'h04A3,4);
TASK_PP(16'h04A4,4);
TASK_PP(16'h04A5,4);
TASK_PP(16'h04A6,4);
TASK_PP(16'h04A7,4);
TASK_PP(16'h04A8,4);
TASK_PP(16'h04A9,4);
TASK_PP(16'h04AA,4);
TASK_PP(16'h04AB,4);
TASK_PP(16'h04AC,4);
TASK_PP(16'h04AD,4);
TASK_PP(16'h04AE,4);
TASK_PP(16'h04AF,4);
TASK_PP(16'h04B0,4);
TASK_PP(16'h04B1,4);
TASK_PP(16'h04B2,4);
TASK_PP(16'h04B3,4);
TASK_PP(16'h04B4,4);
TASK_PP(16'h04B5,4);
TASK_PP(16'h04B6,4);
TASK_PP(16'h04B7,4);
TASK_PP(16'h04B8,4);
TASK_PP(16'h04B9,4);
TASK_PP(16'h04BA,4);
TASK_PP(16'h04BB,4);
TASK_PP(16'h04BC,4);
TASK_PP(16'h04BD,4);
TASK_PP(16'h04BE,4);
TASK_PP(16'h04BF,4);
TASK_PP(16'h04C0,4);
TASK_PP(16'h04C1,4);
TASK_PP(16'h04C2,4);
TASK_PP(16'h04C3,4);
TASK_PP(16'h04C4,4);
TASK_PP(16'h04C5,4);
TASK_PP(16'h04C6,4);
TASK_PP(16'h04C7,4);
TASK_PP(16'h04C8,4);
TASK_PP(16'h04C9,4);
TASK_PP(16'h04CA,4);
TASK_PP(16'h04CB,4);
TASK_PP(16'h04CC,4);
TASK_PP(16'h04CD,4);
TASK_PP(16'h04CE,4);
TASK_PP(16'h04CF,4);
TASK_PP(16'h04D0,4);
TASK_PP(16'h04D1,4);
TASK_PP(16'h04D2,4);
TASK_PP(16'h04D3,4);
TASK_PP(16'h04D4,4);
TASK_PP(16'h04D5,4);
TASK_PP(16'h04D6,4);
TASK_PP(16'h04D7,4);
TASK_PP(16'h04D8,4);
TASK_PP(16'h04D9,4);
TASK_PP(16'h04DA,4);
TASK_PP(16'h04DB,4);
TASK_PP(16'h04DC,4);
TASK_PP(16'h04DD,4);
TASK_PP(16'h04DE,4);
TASK_PP(16'h04DF,4);
TASK_PP(16'h04E0,4);
TASK_PP(16'h04E1,4);
TASK_PP(16'h04E2,4);
TASK_PP(16'h04E3,4);
TASK_PP(16'h04E4,4);
TASK_PP(16'h04E5,4);
TASK_PP(16'h04E6,4);
TASK_PP(16'h04E7,4);
TASK_PP(16'h04E8,4);
TASK_PP(16'h04E9,4);
TASK_PP(16'h04EA,4);
TASK_PP(16'h04EB,4);
TASK_PP(16'h04EC,4);
TASK_PP(16'h04ED,4);
TASK_PP(16'h04EE,4);
TASK_PP(16'h04EF,4);
TASK_PP(16'h04F0,4);
TASK_PP(16'h04F1,4);
TASK_PP(16'h04F2,4);
TASK_PP(16'h04F3,4);
TASK_PP(16'h04F4,4);
TASK_PP(16'h04F5,4);
TASK_PP(16'h04F6,4);
TASK_PP(16'h04F7,4);
TASK_PP(16'h04F8,4);
TASK_PP(16'h04F9,4);
TASK_PP(16'h04FA,4);
TASK_PP(16'h04FB,4);
TASK_PP(16'h04FC,4);
TASK_PP(16'h04FD,4);
TASK_PP(16'h04FE,4);
TASK_PP(16'h04FF,4);
TASK_PP(16'h0500,4);
TASK_PP(16'h0501,4);
TASK_PP(16'h0502,4);
TASK_PP(16'h0503,4);
TASK_PP(16'h0504,4);
TASK_PP(16'h0505,4);
TASK_PP(16'h0506,4);
TASK_PP(16'h0507,4);
TASK_PP(16'h0508,4);
TASK_PP(16'h0509,4);
TASK_PP(16'h050A,4);
TASK_PP(16'h050B,4);
TASK_PP(16'h050C,4);
TASK_PP(16'h050D,4);
TASK_PP(16'h050E,4);
TASK_PP(16'h050F,4);
TASK_PP(16'h0510,4);
TASK_PP(16'h0511,4);
TASK_PP(16'h0512,4);
TASK_PP(16'h0513,4);
TASK_PP(16'h0514,4);
TASK_PP(16'h0515,4);
TASK_PP(16'h0516,4);
TASK_PP(16'h0517,4);
TASK_PP(16'h0518,4);
TASK_PP(16'h0519,4);
TASK_PP(16'h051A,4);
TASK_PP(16'h051B,4);
TASK_PP(16'h051C,4);
TASK_PP(16'h051D,4);
TASK_PP(16'h051E,4);
TASK_PP(16'h051F,4);
TASK_PP(16'h0520,4);
TASK_PP(16'h0521,4);
TASK_PP(16'h0522,4);
TASK_PP(16'h0523,4);
TASK_PP(16'h0524,4);
TASK_PP(16'h0525,4);
TASK_PP(16'h0526,4);
TASK_PP(16'h0527,4);
TASK_PP(16'h0528,4);
TASK_PP(16'h0529,4);
TASK_PP(16'h052A,4);
TASK_PP(16'h052B,4);
TASK_PP(16'h052C,4);
TASK_PP(16'h052D,4);
TASK_PP(16'h052E,4);
TASK_PP(16'h052F,4);
TASK_PP(16'h0530,4);
TASK_PP(16'h0531,4);
TASK_PP(16'h0532,4);
TASK_PP(16'h0533,4);
TASK_PP(16'h0534,4);
TASK_PP(16'h0535,4);
TASK_PP(16'h0536,4);
TASK_PP(16'h0537,4);
TASK_PP(16'h0538,4);
TASK_PP(16'h0539,4);
TASK_PP(16'h053A,4);
TASK_PP(16'h053B,4);
TASK_PP(16'h053C,4);
TASK_PP(16'h053D,4);
TASK_PP(16'h053E,4);
TASK_PP(16'h053F,4);
TASK_PP(16'h0540,4);
TASK_PP(16'h0541,4);
TASK_PP(16'h0542,4);
TASK_PP(16'h0543,4);
TASK_PP(16'h0544,4);
TASK_PP(16'h0545,4);
TASK_PP(16'h0546,4);
TASK_PP(16'h0547,4);
TASK_PP(16'h0548,4);
TASK_PP(16'h0549,4);
TASK_PP(16'h054A,4);
TASK_PP(16'h054B,4);
TASK_PP(16'h054C,4);
TASK_PP(16'h054D,4);
TASK_PP(16'h054E,4);
TASK_PP(16'h054F,4);
TASK_PP(16'h0550,4);
TASK_PP(16'h0551,4);
TASK_PP(16'h0552,4);
TASK_PP(16'h0553,4);
TASK_PP(16'h0554,4);
TASK_PP(16'h0555,4);
TASK_PP(16'h0556,4);
TASK_PP(16'h0557,4);
TASK_PP(16'h0558,4);
TASK_PP(16'h0559,4);
TASK_PP(16'h055A,4);
TASK_PP(16'h055B,4);
TASK_PP(16'h055C,4);
TASK_PP(16'h055D,4);
TASK_PP(16'h055E,4);
TASK_PP(16'h055F,4);
TASK_PP(16'h0560,4);
TASK_PP(16'h0561,4);
TASK_PP(16'h0562,4);
TASK_PP(16'h0563,4);
TASK_PP(16'h0564,4);
TASK_PP(16'h0565,4);
TASK_PP(16'h0566,4);
TASK_PP(16'h0567,4);
TASK_PP(16'h0568,4);
TASK_PP(16'h0569,4);
TASK_PP(16'h056A,4);
TASK_PP(16'h056B,4);
TASK_PP(16'h056C,4);
TASK_PP(16'h056D,4);
TASK_PP(16'h056E,4);
TASK_PP(16'h056F,4);
TASK_PP(16'h0570,4);
TASK_PP(16'h0571,4);
TASK_PP(16'h0572,4);
TASK_PP(16'h0573,4);
TASK_PP(16'h0574,4);
TASK_PP(16'h0575,4);
TASK_PP(16'h0576,4);
TASK_PP(16'h0577,4);
TASK_PP(16'h0578,4);
TASK_PP(16'h0579,4);
TASK_PP(16'h057A,4);
TASK_PP(16'h057B,4);
TASK_PP(16'h057C,4);
TASK_PP(16'h057D,4);
TASK_PP(16'h057E,4);
TASK_PP(16'h057F,4);
TASK_PP(16'h0580,4);
TASK_PP(16'h0581,4);
TASK_PP(16'h0582,4);
TASK_PP(16'h0583,4);
TASK_PP(16'h0584,4);
TASK_PP(16'h0585,4);
TASK_PP(16'h0586,4);
TASK_PP(16'h0587,4);
TASK_PP(16'h0588,4);
TASK_PP(16'h0589,4);
TASK_PP(16'h058A,4);
TASK_PP(16'h058B,4);
TASK_PP(16'h058C,4);
TASK_PP(16'h058D,4);
TASK_PP(16'h058E,4);
TASK_PP(16'h058F,4);
TASK_PP(16'h0590,4);
TASK_PP(16'h0591,4);
TASK_PP(16'h0592,4);
TASK_PP(16'h0593,4);
TASK_PP(16'h0594,4);
TASK_PP(16'h0595,4);
TASK_PP(16'h0596,4);
TASK_PP(16'h0597,4);
TASK_PP(16'h0598,4);
TASK_PP(16'h0599,4);
TASK_PP(16'h059A,4);
TASK_PP(16'h059B,4);
TASK_PP(16'h059C,4);
TASK_PP(16'h059D,4);
TASK_PP(16'h059E,4);
TASK_PP(16'h059F,4);
TASK_PP(16'h05A0,4);
TASK_PP(16'h05A1,4);
TASK_PP(16'h05A2,4);
TASK_PP(16'h05A3,4);
TASK_PP(16'h05A4,4);
TASK_PP(16'h05A5,4);
TASK_PP(16'h05A6,4);
TASK_PP(16'h05A7,4);
TASK_PP(16'h05A8,4);
TASK_PP(16'h05A9,4);
TASK_PP(16'h05AA,4);
TASK_PP(16'h05AB,4);
TASK_PP(16'h05AC,4);
TASK_PP(16'h05AD,4);
TASK_PP(16'h05AE,4);
TASK_PP(16'h05AF,4);
TASK_PP(16'h05B0,4);
TASK_PP(16'h05B1,4);
TASK_PP(16'h05B2,4);
TASK_PP(16'h05B3,4);
TASK_PP(16'h05B4,4);
TASK_PP(16'h05B5,4);
TASK_PP(16'h05B6,4);
TASK_PP(16'h05B7,4);
TASK_PP(16'h05B8,4);
TASK_PP(16'h05B9,4);
TASK_PP(16'h05BA,4);
TASK_PP(16'h05BB,4);
TASK_PP(16'h05BC,4);
TASK_PP(16'h05BD,4);
TASK_PP(16'h05BE,4);
TASK_PP(16'h05BF,4);
TASK_PP(16'h05C0,4);
TASK_PP(16'h05C1,4);
TASK_PP(16'h05C2,4);
TASK_PP(16'h05C3,4);
TASK_PP(16'h05C4,4);
TASK_PP(16'h05C5,4);
TASK_PP(16'h05C6,4);
TASK_PP(16'h05C7,4);
TASK_PP(16'h05C8,4);
TASK_PP(16'h05C9,4);
TASK_PP(16'h05CA,4);
TASK_PP(16'h05CB,4);
TASK_PP(16'h05CC,4);
TASK_PP(16'h05CD,4);
TASK_PP(16'h05CE,4);
TASK_PP(16'h05CF,4);
TASK_PP(16'h05D0,4);
TASK_PP(16'h05D1,4);
TASK_PP(16'h05D2,4);
TASK_PP(16'h05D3,4);
TASK_PP(16'h05D4,4);
TASK_PP(16'h05D5,4);
TASK_PP(16'h05D6,4);
TASK_PP(16'h05D7,4);
TASK_PP(16'h05D8,4);
TASK_PP(16'h05D9,4);
TASK_PP(16'h05DA,4);
TASK_PP(16'h05DB,4);
TASK_PP(16'h05DC,4);
TASK_PP(16'h05DD,4);
TASK_PP(16'h05DE,4);
TASK_PP(16'h05DF,4);
TASK_PP(16'h05E0,4);
TASK_PP(16'h05E1,4);
TASK_PP(16'h05E2,4);
TASK_PP(16'h05E3,4);
TASK_PP(16'h05E4,4);
TASK_PP(16'h05E5,4);
TASK_PP(16'h05E6,4);
TASK_PP(16'h05E7,4);
TASK_PP(16'h05E8,4);
TASK_PP(16'h05E9,4);
TASK_PP(16'h05EA,4);
TASK_PP(16'h05EB,4);
TASK_PP(16'h05EC,4);
TASK_PP(16'h05ED,4);
TASK_PP(16'h05EE,4);
TASK_PP(16'h05EF,4);
TASK_PP(16'h05F0,4);
TASK_PP(16'h05F1,4);
TASK_PP(16'h05F2,4);
TASK_PP(16'h05F3,4);
TASK_PP(16'h05F4,4);
TASK_PP(16'h05F5,4);
TASK_PP(16'h05F6,4);
TASK_PP(16'h05F7,4);
TASK_PP(16'h05F8,4);
TASK_PP(16'h05F9,4);
TASK_PP(16'h05FA,4);
TASK_PP(16'h05FB,4);
TASK_PP(16'h05FC,4);
TASK_PP(16'h05FD,4);
TASK_PP(16'h05FE,4);
TASK_PP(16'h05FF,4);
TASK_PP(16'h0600,4);
TASK_PP(16'h0601,4);
TASK_PP(16'h0602,4);
TASK_PP(16'h0603,4);
TASK_PP(16'h0604,4);
TASK_PP(16'h0605,4);
TASK_PP(16'h0606,4);
TASK_PP(16'h0607,4);
TASK_PP(16'h0608,4);
TASK_PP(16'h0609,4);
TASK_PP(16'h060A,4);
TASK_PP(16'h060B,4);
TASK_PP(16'h060C,4);
TASK_PP(16'h060D,4);
TASK_PP(16'h060E,4);
TASK_PP(16'h060F,4);
TASK_PP(16'h0610,4);
TASK_PP(16'h0611,4);
TASK_PP(16'h0612,4);
TASK_PP(16'h0613,4);
TASK_PP(16'h0614,4);
TASK_PP(16'h0615,4);
TASK_PP(16'h0616,4);
TASK_PP(16'h0617,4);
TASK_PP(16'h0618,4);
TASK_PP(16'h0619,4);
TASK_PP(16'h061A,4);
TASK_PP(16'h061B,4);
TASK_PP(16'h061C,4);
TASK_PP(16'h061D,4);
TASK_PP(16'h061E,4);
TASK_PP(16'h061F,4);
TASK_PP(16'h0620,4);
TASK_PP(16'h0621,4);
TASK_PP(16'h0622,4);
TASK_PP(16'h0623,4);
TASK_PP(16'h0624,4);
TASK_PP(16'h0625,4);
TASK_PP(16'h0626,4);
TASK_PP(16'h0627,4);
TASK_PP(16'h0628,4);
TASK_PP(16'h0629,4);
TASK_PP(16'h062A,4);
TASK_PP(16'h062B,4);
TASK_PP(16'h062C,4);
TASK_PP(16'h062D,4);
TASK_PP(16'h062E,4);
TASK_PP(16'h062F,4);
TASK_PP(16'h0630,4);
TASK_PP(16'h0631,4);
TASK_PP(16'h0632,4);
TASK_PP(16'h0633,4);
TASK_PP(16'h0634,4);
TASK_PP(16'h0635,4);
TASK_PP(16'h0636,4);
TASK_PP(16'h0637,4);
TASK_PP(16'h0638,4);
TASK_PP(16'h0639,4);
TASK_PP(16'h063A,4);
TASK_PP(16'h063B,4);
TASK_PP(16'h063C,4);
TASK_PP(16'h063D,4);
TASK_PP(16'h063E,4);
TASK_PP(16'h063F,4);
TASK_PP(16'h0640,4);
TASK_PP(16'h0641,4);
TASK_PP(16'h0642,4);
TASK_PP(16'h0643,4);
TASK_PP(16'h0644,4);
TASK_PP(16'h0645,4);
TASK_PP(16'h0646,4);
TASK_PP(16'h0647,4);
TASK_PP(16'h0648,4);
TASK_PP(16'h0649,4);
TASK_PP(16'h064A,4);
TASK_PP(16'h064B,4);
TASK_PP(16'h064C,4);
TASK_PP(16'h064D,4);
TASK_PP(16'h064E,4);
TASK_PP(16'h064F,4);
TASK_PP(16'h0650,4);
TASK_PP(16'h0651,4);
TASK_PP(16'h0652,4);
TASK_PP(16'h0653,4);
TASK_PP(16'h0654,4);
TASK_PP(16'h0655,4);
TASK_PP(16'h0656,4);
TASK_PP(16'h0657,4);
TASK_PP(16'h0658,4);
TASK_PP(16'h0659,4);
TASK_PP(16'h065A,4);
TASK_PP(16'h065B,4);
TASK_PP(16'h065C,4);
TASK_PP(16'h065D,4);
TASK_PP(16'h065E,4);
TASK_PP(16'h065F,4);
TASK_PP(16'h0660,4);
TASK_PP(16'h0661,4);
TASK_PP(16'h0662,4);
TASK_PP(16'h0663,4);
TASK_PP(16'h0664,4);
TASK_PP(16'h0665,4);
TASK_PP(16'h0666,4);
TASK_PP(16'h0667,4);
TASK_PP(16'h0668,4);
TASK_PP(16'h0669,4);
TASK_PP(16'h066A,4);
TASK_PP(16'h066B,4);
TASK_PP(16'h066C,4);
TASK_PP(16'h066D,4);
TASK_PP(16'h066E,4);
TASK_PP(16'h066F,4);
TASK_PP(16'h0670,4);
TASK_PP(16'h0671,4);
TASK_PP(16'h0672,4);
TASK_PP(16'h0673,4);
TASK_PP(16'h0674,4);
TASK_PP(16'h0675,4);
TASK_PP(16'h0676,4);
TASK_PP(16'h0677,4);
TASK_PP(16'h0678,4);
TASK_PP(16'h0679,4);
TASK_PP(16'h067A,4);
TASK_PP(16'h067B,4);
TASK_PP(16'h067C,4);
TASK_PP(16'h067D,4);
TASK_PP(16'h067E,4);
TASK_PP(16'h067F,4);
TASK_PP(16'h0680,4);
TASK_PP(16'h0681,4);
TASK_PP(16'h0682,4);
TASK_PP(16'h0683,4);
TASK_PP(16'h0684,4);
TASK_PP(16'h0685,4);
TASK_PP(16'h0686,4);
TASK_PP(16'h0687,4);
TASK_PP(16'h0688,4);
TASK_PP(16'h0689,4);
TASK_PP(16'h068A,4);
TASK_PP(16'h068B,4);
TASK_PP(16'h068C,4);
TASK_PP(16'h068D,4);
TASK_PP(16'h068E,4);
TASK_PP(16'h068F,4);
TASK_PP(16'h0690,4);
TASK_PP(16'h0691,4);
TASK_PP(16'h0692,4);
TASK_PP(16'h0693,4);
TASK_PP(16'h0694,4);
TASK_PP(16'h0695,4);
TASK_PP(16'h0696,4);
TASK_PP(16'h0697,4);
TASK_PP(16'h0698,4);
TASK_PP(16'h0699,4);
TASK_PP(16'h069A,4);
TASK_PP(16'h069B,4);
TASK_PP(16'h069C,4);
TASK_PP(16'h069D,4);
TASK_PP(16'h069E,4);
TASK_PP(16'h069F,4);
TASK_PP(16'h06A0,4);
TASK_PP(16'h06A1,4);
TASK_PP(16'h06A2,4);
TASK_PP(16'h06A3,4);
TASK_PP(16'h06A4,4);
TASK_PP(16'h06A5,4);
TASK_PP(16'h06A6,4);
TASK_PP(16'h06A7,4);
TASK_PP(16'h06A8,4);
TASK_PP(16'h06A9,4);
TASK_PP(16'h06AA,4);
TASK_PP(16'h06AB,4);
TASK_PP(16'h06AC,4);
TASK_PP(16'h06AD,4);
TASK_PP(16'h06AE,4);
TASK_PP(16'h06AF,4);
TASK_PP(16'h06B0,4);
TASK_PP(16'h06B1,4);
TASK_PP(16'h06B2,4);
TASK_PP(16'h06B3,4);
TASK_PP(16'h06B4,4);
TASK_PP(16'h06B5,4);
TASK_PP(16'h06B6,4);
TASK_PP(16'h06B7,4);
TASK_PP(16'h06B8,4);
TASK_PP(16'h06B9,4);
TASK_PP(16'h06BA,4);
TASK_PP(16'h06BB,4);
TASK_PP(16'h06BC,4);
TASK_PP(16'h06BD,4);
TASK_PP(16'h06BE,4);
TASK_PP(16'h06BF,4);
TASK_PP(16'h06C0,4);
TASK_PP(16'h06C1,4);
TASK_PP(16'h06C2,4);
TASK_PP(16'h06C3,4);
TASK_PP(16'h06C4,4);
TASK_PP(16'h06C5,4);
TASK_PP(16'h06C6,4);
TASK_PP(16'h06C7,4);
TASK_PP(16'h06C8,4);
TASK_PP(16'h06C9,4);
TASK_PP(16'h06CA,4);
TASK_PP(16'h06CB,4);
TASK_PP(16'h06CC,4);
TASK_PP(16'h06CD,4);
TASK_PP(16'h06CE,4);
TASK_PP(16'h06CF,4);
TASK_PP(16'h06D0,4);
TASK_PP(16'h06D1,4);
TASK_PP(16'h06D2,4);
TASK_PP(16'h06D3,4);
TASK_PP(16'h06D4,4);
TASK_PP(16'h06D5,4);
TASK_PP(16'h06D6,4);
TASK_PP(16'h06D7,4);
TASK_PP(16'h06D8,4);
TASK_PP(16'h06D9,4);
TASK_PP(16'h06DA,4);
TASK_PP(16'h06DB,4);
TASK_PP(16'h06DC,4);
TASK_PP(16'h06DD,4);
TASK_PP(16'h06DE,4);
TASK_PP(16'h06DF,4);
TASK_PP(16'h06E0,4);
TASK_PP(16'h06E1,4);
TASK_PP(16'h06E2,4);
TASK_PP(16'h06E3,4);
TASK_PP(16'h06E4,4);
TASK_PP(16'h06E5,4);
TASK_PP(16'h06E6,4);
TASK_PP(16'h06E7,4);
TASK_PP(16'h06E8,4);
TASK_PP(16'h06E9,4);
TASK_PP(16'h06EA,4);
TASK_PP(16'h06EB,4);
TASK_PP(16'h06EC,4);
TASK_PP(16'h06ED,4);
TASK_PP(16'h06EE,4);
TASK_PP(16'h06EF,4);
TASK_PP(16'h06F0,4);
TASK_PP(16'h06F1,4);
TASK_PP(16'h06F2,4);
TASK_PP(16'h06F3,4);
TASK_PP(16'h06F4,4);
TASK_PP(16'h06F5,4);
TASK_PP(16'h06F6,4);
TASK_PP(16'h06F7,4);
TASK_PP(16'h06F8,4);
TASK_PP(16'h06F9,4);
TASK_PP(16'h06FA,4);
TASK_PP(16'h06FB,4);
TASK_PP(16'h06FC,4);
TASK_PP(16'h06FD,4);
TASK_PP(16'h06FE,4);
TASK_PP(16'h06FF,4);
TASK_PP(16'h0700,4);
TASK_PP(16'h0701,4);
TASK_PP(16'h0702,4);
TASK_PP(16'h0703,4);
TASK_PP(16'h0704,4);
TASK_PP(16'h0705,4);
TASK_PP(16'h0706,4);
TASK_PP(16'h0707,4);
TASK_PP(16'h0708,4);
TASK_PP(16'h0709,4);
TASK_PP(16'h070A,4);
TASK_PP(16'h070B,4);
TASK_PP(16'h070C,4);
TASK_PP(16'h070D,4);
TASK_PP(16'h070E,4);
TASK_PP(16'h070F,4);
TASK_PP(16'h0710,4);
TASK_PP(16'h0711,4);
TASK_PP(16'h0712,4);
TASK_PP(16'h0713,4);
TASK_PP(16'h0714,4);
TASK_PP(16'h0715,4);
TASK_PP(16'h0716,4);
TASK_PP(16'h0717,4);
TASK_PP(16'h0718,4);
TASK_PP(16'h0719,4);
TASK_PP(16'h071A,4);
TASK_PP(16'h071B,4);
TASK_PP(16'h071C,4);
TASK_PP(16'h071D,4);
TASK_PP(16'h071E,4);
TASK_PP(16'h071F,4);
TASK_PP(16'h0720,4);
TASK_PP(16'h0721,4);
TASK_PP(16'h0722,4);
TASK_PP(16'h0723,4);
TASK_PP(16'h0724,4);
TASK_PP(16'h0725,4);
TASK_PP(16'h0726,4);
TASK_PP(16'h0727,4);
TASK_PP(16'h0728,4);
TASK_PP(16'h0729,4);
TASK_PP(16'h072A,4);
TASK_PP(16'h072B,4);
TASK_PP(16'h072C,4);
TASK_PP(16'h072D,4);
TASK_PP(16'h072E,4);
TASK_PP(16'h072F,4);
TASK_PP(16'h0730,4);
TASK_PP(16'h0731,4);
TASK_PP(16'h0732,4);
TASK_PP(16'h0733,4);
TASK_PP(16'h0734,4);
TASK_PP(16'h0735,4);
TASK_PP(16'h0736,4);
TASK_PP(16'h0737,4);
TASK_PP(16'h0738,4);
TASK_PP(16'h0739,4);
TASK_PP(16'h073A,4);
TASK_PP(16'h073B,4);
TASK_PP(16'h073C,4);
TASK_PP(16'h073D,4);
TASK_PP(16'h073E,4);
TASK_PP(16'h073F,4);
TASK_PP(16'h0740,4);
TASK_PP(16'h0741,4);
TASK_PP(16'h0742,4);
TASK_PP(16'h0743,4);
TASK_PP(16'h0744,4);
TASK_PP(16'h0745,4);
TASK_PP(16'h0746,4);
TASK_PP(16'h0747,4);
TASK_PP(16'h0748,4);
TASK_PP(16'h0749,4);
TASK_PP(16'h074A,4);
TASK_PP(16'h074B,4);
TASK_PP(16'h074C,4);
TASK_PP(16'h074D,4);
TASK_PP(16'h074E,4);
TASK_PP(16'h074F,4);
TASK_PP(16'h0750,4);
TASK_PP(16'h0751,4);
TASK_PP(16'h0752,4);
TASK_PP(16'h0753,4);
TASK_PP(16'h0754,4);
TASK_PP(16'h0755,4);
TASK_PP(16'h0756,4);
TASK_PP(16'h0757,4);
TASK_PP(16'h0758,4);
TASK_PP(16'h0759,4);
TASK_PP(16'h075A,4);
TASK_PP(16'h075B,4);
TASK_PP(16'h075C,4);
TASK_PP(16'h075D,4);
TASK_PP(16'h075E,4);
TASK_PP(16'h075F,4);
TASK_PP(16'h0760,4);
TASK_PP(16'h0761,4);
TASK_PP(16'h0762,4);
TASK_PP(16'h0763,4);
TASK_PP(16'h0764,4);
TASK_PP(16'h0765,4);
TASK_PP(16'h0766,4);
TASK_PP(16'h0767,4);
TASK_PP(16'h0768,4);
TASK_PP(16'h0769,4);
TASK_PP(16'h076A,4);
TASK_PP(16'h076B,4);
TASK_PP(16'h076C,4);
TASK_PP(16'h076D,4);
TASK_PP(16'h076E,4);
TASK_PP(16'h076F,4);
TASK_PP(16'h0770,4);
TASK_PP(16'h0771,4);
TASK_PP(16'h0772,4);
TASK_PP(16'h0773,4);
TASK_PP(16'h0774,4);
TASK_PP(16'h0775,4);
TASK_PP(16'h0776,4);
TASK_PP(16'h0777,4);
TASK_PP(16'h0778,4);
TASK_PP(16'h0779,4);
TASK_PP(16'h077A,4);
TASK_PP(16'h077B,4);
TASK_PP(16'h077C,4);
TASK_PP(16'h077D,4);
TASK_PP(16'h077E,4);
TASK_PP(16'h077F,4);
TASK_PP(16'h0780,4);
TASK_PP(16'h0781,4);
TASK_PP(16'h0782,4);
TASK_PP(16'h0783,4);
TASK_PP(16'h0784,4);
TASK_PP(16'h0785,4);
TASK_PP(16'h0786,4);
TASK_PP(16'h0787,4);
TASK_PP(16'h0788,4);
TASK_PP(16'h0789,4);
TASK_PP(16'h078A,4);
TASK_PP(16'h078B,4);
TASK_PP(16'h078C,4);
TASK_PP(16'h078D,4);
TASK_PP(16'h078E,4);
TASK_PP(16'h078F,4);
TASK_PP(16'h0790,4);
TASK_PP(16'h0791,4);
TASK_PP(16'h0792,4);
TASK_PP(16'h0793,4);
TASK_PP(16'h0794,4);
TASK_PP(16'h0795,4);
TASK_PP(16'h0796,4);
TASK_PP(16'h0797,4);
TASK_PP(16'h0798,4);
TASK_PP(16'h0799,4);
TASK_PP(16'h079A,4);
TASK_PP(16'h079B,4);
TASK_PP(16'h079C,4);
TASK_PP(16'h079D,4);
TASK_PP(16'h079E,4);
TASK_PP(16'h079F,4);
TASK_PP(16'h07A0,4);
TASK_PP(16'h07A1,4);
TASK_PP(16'h07A2,4);
TASK_PP(16'h07A3,4);
TASK_PP(16'h07A4,4);
TASK_PP(16'h07A5,4);
TASK_PP(16'h07A6,4);
TASK_PP(16'h07A7,4);
TASK_PP(16'h07A8,4);
TASK_PP(16'h07A9,4);
TASK_PP(16'h07AA,4);
TASK_PP(16'h07AB,4);
TASK_PP(16'h07AC,4);
TASK_PP(16'h07AD,4);
TASK_PP(16'h07AE,4);
TASK_PP(16'h07AF,4);
TASK_PP(16'h07B0,4);
TASK_PP(16'h07B1,4);
TASK_PP(16'h07B2,4);
TASK_PP(16'h07B3,4);
TASK_PP(16'h07B4,4);
TASK_PP(16'h07B5,4);
TASK_PP(16'h07B6,4);
TASK_PP(16'h07B7,4);
TASK_PP(16'h07B8,4);
TASK_PP(16'h07B9,4);
TASK_PP(16'h07BA,4);
TASK_PP(16'h07BB,4);
TASK_PP(16'h07BC,4);
TASK_PP(16'h07BD,4);
TASK_PP(16'h07BE,4);
TASK_PP(16'h07BF,4);
TASK_PP(16'h07C0,4);
TASK_PP(16'h07C1,4);
TASK_PP(16'h07C2,4);
TASK_PP(16'h07C3,4);
TASK_PP(16'h07C4,4);
TASK_PP(16'h07C5,4);
TASK_PP(16'h07C6,4);
TASK_PP(16'h07C7,4);
TASK_PP(16'h07C8,4);
TASK_PP(16'h07C9,4);
TASK_PP(16'h07CA,4);
TASK_PP(16'h07CB,4);
TASK_PP(16'h07CC,4);
TASK_PP(16'h07CD,4);
TASK_PP(16'h07CE,4);
TASK_PP(16'h07CF,4);
TASK_PP(16'h07D0,4);
TASK_PP(16'h07D1,4);
TASK_PP(16'h07D2,4);
TASK_PP(16'h07D3,4);
TASK_PP(16'h07D4,4);
TASK_PP(16'h07D5,4);
TASK_PP(16'h07D6,4);
TASK_PP(16'h07D7,4);
TASK_PP(16'h07D8,4);
TASK_PP(16'h07D9,4);
TASK_PP(16'h07DA,4);
TASK_PP(16'h07DB,4);
TASK_PP(16'h07DC,4);
TASK_PP(16'h07DD,4);
TASK_PP(16'h07DE,4);
TASK_PP(16'h07DF,4);
TASK_PP(16'h07E0,4);
TASK_PP(16'h07E1,4);
TASK_PP(16'h07E2,4);
TASK_PP(16'h07E3,4);
TASK_PP(16'h07E4,4);
TASK_PP(16'h07E5,4);
TASK_PP(16'h07E6,4);
TASK_PP(16'h07E7,4);
TASK_PP(16'h07E8,4);
TASK_PP(16'h07E9,4);
TASK_PP(16'h07EA,4);
TASK_PP(16'h07EB,4);
TASK_PP(16'h07EC,4);
TASK_PP(16'h07ED,4);
TASK_PP(16'h07EE,4);
TASK_PP(16'h07EF,4);
TASK_PP(16'h07F0,4);
TASK_PP(16'h07F1,4);
TASK_PP(16'h07F2,4);
TASK_PP(16'h07F3,4);
TASK_PP(16'h07F4,4);
TASK_PP(16'h07F5,4);
TASK_PP(16'h07F6,4);
TASK_PP(16'h07F7,4);
TASK_PP(16'h07F8,4);
TASK_PP(16'h07F9,4);
TASK_PP(16'h07FA,4);
TASK_PP(16'h07FB,4);
TASK_PP(16'h07FC,4);
TASK_PP(16'h07FD,4);
TASK_PP(16'h07FE,4);
TASK_PP(16'h07FF,4);
TASK_PP(16'h0800,4);
TASK_PP(16'h0801,4);
TASK_PP(16'h0802,4);
TASK_PP(16'h0803,4);
TASK_PP(16'h0804,4);
TASK_PP(16'h0805,4);
TASK_PP(16'h0806,4);
TASK_PP(16'h0807,4);
TASK_PP(16'h0808,4);
TASK_PP(16'h0809,4);
TASK_PP(16'h080A,4);
TASK_PP(16'h080B,4);
TASK_PP(16'h080C,4);
TASK_PP(16'h080D,4);
TASK_PP(16'h080E,4);
TASK_PP(16'h080F,4);
TASK_PP(16'h0810,4);
TASK_PP(16'h0811,4);
TASK_PP(16'h0812,4);
TASK_PP(16'h0813,4);
TASK_PP(16'h0814,4);
TASK_PP(16'h0815,4);
TASK_PP(16'h0816,4);
TASK_PP(16'h0817,4);
TASK_PP(16'h0818,4);
TASK_PP(16'h0819,4);
TASK_PP(16'h081A,4);
TASK_PP(16'h081B,4);
TASK_PP(16'h081C,4);
TASK_PP(16'h081D,4);
TASK_PP(16'h081E,4);
TASK_PP(16'h081F,4);
TASK_PP(16'h0820,4);
TASK_PP(16'h0821,4);
TASK_PP(16'h0822,4);
TASK_PP(16'h0823,4);
TASK_PP(16'h0824,4);
TASK_PP(16'h0825,4);
TASK_PP(16'h0826,4);
TASK_PP(16'h0827,4);
TASK_PP(16'h0828,4);
TASK_PP(16'h0829,4);
TASK_PP(16'h082A,4);
TASK_PP(16'h082B,4);
TASK_PP(16'h082C,4);
TASK_PP(16'h082D,4);
TASK_PP(16'h082E,4);
TASK_PP(16'h082F,4);
TASK_PP(16'h0830,4);
TASK_PP(16'h0831,4);
TASK_PP(16'h0832,4);
TASK_PP(16'h0833,4);
TASK_PP(16'h0834,4);
TASK_PP(16'h0835,4);
TASK_PP(16'h0836,4);
TASK_PP(16'h0837,4);
TASK_PP(16'h0838,4);
TASK_PP(16'h0839,4);
TASK_PP(16'h083A,4);
TASK_PP(16'h083B,4);
TASK_PP(16'h083C,4);
TASK_PP(16'h083D,4);
TASK_PP(16'h083E,4);
TASK_PP(16'h083F,4);
TASK_PP(16'h0840,4);
TASK_PP(16'h0841,4);
TASK_PP(16'h0842,4);
TASK_PP(16'h0843,4);
TASK_PP(16'h0844,4);
TASK_PP(16'h0845,4);
TASK_PP(16'h0846,4);
TASK_PP(16'h0847,4);
TASK_PP(16'h0848,4);
TASK_PP(16'h0849,4);
TASK_PP(16'h084A,4);
TASK_PP(16'h084B,4);
TASK_PP(16'h084C,4);
TASK_PP(16'h084D,4);
TASK_PP(16'h084E,4);
TASK_PP(16'h084F,4);
TASK_PP(16'h0850,4);
TASK_PP(16'h0851,4);
TASK_PP(16'h0852,4);
TASK_PP(16'h0853,4);
TASK_PP(16'h0854,4);
TASK_PP(16'h0855,4);
TASK_PP(16'h0856,4);
TASK_PP(16'h0857,4);
TASK_PP(16'h0858,4);
TASK_PP(16'h0859,4);
TASK_PP(16'h085A,4);
TASK_PP(16'h085B,4);
TASK_PP(16'h085C,4);
TASK_PP(16'h085D,4);
TASK_PP(16'h085E,4);
TASK_PP(16'h085F,4);
TASK_PP(16'h0860,4);
TASK_PP(16'h0861,4);
TASK_PP(16'h0862,4);
TASK_PP(16'h0863,4);
TASK_PP(16'h0864,4);
TASK_PP(16'h0865,4);
TASK_PP(16'h0866,4);
TASK_PP(16'h0867,4);
TASK_PP(16'h0868,4);
TASK_PP(16'h0869,4);
TASK_PP(16'h086A,4);
TASK_PP(16'h086B,4);
TASK_PP(16'h086C,4);
TASK_PP(16'h086D,4);
TASK_PP(16'h086E,4);
TASK_PP(16'h086F,4);
TASK_PP(16'h0870,4);
TASK_PP(16'h0871,4);
TASK_PP(16'h0872,4);
TASK_PP(16'h0873,4);
TASK_PP(16'h0874,4);
TASK_PP(16'h0875,4);
TASK_PP(16'h0876,4);
TASK_PP(16'h0877,4);
TASK_PP(16'h0878,4);
TASK_PP(16'h0879,4);
TASK_PP(16'h087A,4);
TASK_PP(16'h087B,4);
TASK_PP(16'h087C,4);
TASK_PP(16'h087D,4);
TASK_PP(16'h087E,4);
TASK_PP(16'h087F,4);
TASK_PP(16'h0880,4);
TASK_PP(16'h0881,4);
TASK_PP(16'h0882,4);
TASK_PP(16'h0883,4);
TASK_PP(16'h0884,4);
TASK_PP(16'h0885,4);
TASK_PP(16'h0886,4);
TASK_PP(16'h0887,4);
TASK_PP(16'h0888,4);
TASK_PP(16'h0889,4);
TASK_PP(16'h088A,4);
TASK_PP(16'h088B,4);
TASK_PP(16'h088C,4);
TASK_PP(16'h088D,4);
TASK_PP(16'h088E,4);
TASK_PP(16'h088F,4);
TASK_PP(16'h0890,4);
TASK_PP(16'h0891,4);
TASK_PP(16'h0892,4);
TASK_PP(16'h0893,4);
TASK_PP(16'h0894,4);
TASK_PP(16'h0895,4);
TASK_PP(16'h0896,4);
TASK_PP(16'h0897,4);
TASK_PP(16'h0898,4);
TASK_PP(16'h0899,4);
TASK_PP(16'h089A,4);
TASK_PP(16'h089B,4);
TASK_PP(16'h089C,4);
TASK_PP(16'h089D,4);
TASK_PP(16'h089E,4);
TASK_PP(16'h089F,4);
TASK_PP(16'h08A0,4);
TASK_PP(16'h08A1,4);
TASK_PP(16'h08A2,4);
TASK_PP(16'h08A3,4);
TASK_PP(16'h08A4,4);
TASK_PP(16'h08A5,4);
TASK_PP(16'h08A6,4);
TASK_PP(16'h08A7,4);
TASK_PP(16'h08A8,4);
TASK_PP(16'h08A9,4);
TASK_PP(16'h08AA,4);
TASK_PP(16'h08AB,4);
TASK_PP(16'h08AC,4);
TASK_PP(16'h08AD,4);
TASK_PP(16'h08AE,4);
TASK_PP(16'h08AF,4);
TASK_PP(16'h08B0,4);
TASK_PP(16'h08B1,4);
TASK_PP(16'h08B2,4);
TASK_PP(16'h08B3,4);
TASK_PP(16'h08B4,4);
TASK_PP(16'h08B5,4);
TASK_PP(16'h08B6,4);
TASK_PP(16'h08B7,4);
TASK_PP(16'h08B8,4);
TASK_PP(16'h08B9,4);
TASK_PP(16'h08BA,4);
TASK_PP(16'h08BB,4);
TASK_PP(16'h08BC,4);
TASK_PP(16'h08BD,4);
TASK_PP(16'h08BE,4);
TASK_PP(16'h08BF,4);
TASK_PP(16'h08C0,4);
TASK_PP(16'h08C1,4);
TASK_PP(16'h08C2,4);
TASK_PP(16'h08C3,4);
TASK_PP(16'h08C4,4);
TASK_PP(16'h08C5,4);
TASK_PP(16'h08C6,4);
TASK_PP(16'h08C7,4);
TASK_PP(16'h08C8,4);
TASK_PP(16'h08C9,4);
TASK_PP(16'h08CA,4);
TASK_PP(16'h08CB,4);
TASK_PP(16'h08CC,4);
TASK_PP(16'h08CD,4);
TASK_PP(16'h08CE,4);
TASK_PP(16'h08CF,4);
TASK_PP(16'h08D0,4);
TASK_PP(16'h08D1,4);
TASK_PP(16'h08D2,4);
TASK_PP(16'h08D3,4);
TASK_PP(16'h08D4,4);
TASK_PP(16'h08D5,4);
TASK_PP(16'h08D6,4);
TASK_PP(16'h08D7,4);
TASK_PP(16'h08D8,4);
TASK_PP(16'h08D9,4);
TASK_PP(16'h08DA,4);
TASK_PP(16'h08DB,4);
TASK_PP(16'h08DC,4);
TASK_PP(16'h08DD,4);
TASK_PP(16'h08DE,4);
TASK_PP(16'h08DF,4);
TASK_PP(16'h08E0,4);
TASK_PP(16'h08E1,4);
TASK_PP(16'h08E2,4);
TASK_PP(16'h08E3,4);
TASK_PP(16'h08E4,4);
TASK_PP(16'h08E5,4);
TASK_PP(16'h08E6,4);
TASK_PP(16'h08E7,4);
TASK_PP(16'h08E8,4);
TASK_PP(16'h08E9,4);
TASK_PP(16'h08EA,4);
TASK_PP(16'h08EB,4);
TASK_PP(16'h08EC,4);
TASK_PP(16'h08ED,4);
TASK_PP(16'h08EE,4);
TASK_PP(16'h08EF,4);
TASK_PP(16'h08F0,4);
TASK_PP(16'h08F1,4);
TASK_PP(16'h08F2,4);
TASK_PP(16'h08F3,4);
TASK_PP(16'h08F4,4);
TASK_PP(16'h08F5,4);
TASK_PP(16'h08F6,4);
TASK_PP(16'h08F7,4);
TASK_PP(16'h08F8,4);
TASK_PP(16'h08F9,4);
TASK_PP(16'h08FA,4);
TASK_PP(16'h08FB,4);
TASK_PP(16'h08FC,4);
TASK_PP(16'h08FD,4);
TASK_PP(16'h08FE,4);
TASK_PP(16'h08FF,4);
TASK_PP(16'h0900,4);
TASK_PP(16'h0901,4);
TASK_PP(16'h0902,4);
TASK_PP(16'h0903,4);
TASK_PP(16'h0904,4);
TASK_PP(16'h0905,4);
TASK_PP(16'h0906,4);
TASK_PP(16'h0907,4);
TASK_PP(16'h0908,4);
TASK_PP(16'h0909,4);
TASK_PP(16'h090A,4);
TASK_PP(16'h090B,4);
TASK_PP(16'h090C,4);
TASK_PP(16'h090D,4);
TASK_PP(16'h090E,4);
TASK_PP(16'h090F,4);
TASK_PP(16'h0910,4);
TASK_PP(16'h0911,4);
TASK_PP(16'h0912,4);
TASK_PP(16'h0913,4);
TASK_PP(16'h0914,4);
TASK_PP(16'h0915,4);
TASK_PP(16'h0916,4);
TASK_PP(16'h0917,4);
TASK_PP(16'h0918,4);
TASK_PP(16'h0919,4);
TASK_PP(16'h091A,4);
TASK_PP(16'h091B,4);
TASK_PP(16'h091C,4);
TASK_PP(16'h091D,4);
TASK_PP(16'h091E,4);
TASK_PP(16'h091F,4);
TASK_PP(16'h0920,4);
TASK_PP(16'h0921,4);
TASK_PP(16'h0922,4);
TASK_PP(16'h0923,4);
TASK_PP(16'h0924,4);
TASK_PP(16'h0925,4);
TASK_PP(16'h0926,4);
TASK_PP(16'h0927,4);
TASK_PP(16'h0928,4);
TASK_PP(16'h0929,4);
TASK_PP(16'h092A,4);
TASK_PP(16'h092B,4);
TASK_PP(16'h092C,4);
TASK_PP(16'h092D,4);
TASK_PP(16'h092E,4);
TASK_PP(16'h092F,4);
TASK_PP(16'h0930,4);
TASK_PP(16'h0931,4);
TASK_PP(16'h0932,4);
TASK_PP(16'h0933,4);
TASK_PP(16'h0934,4);
TASK_PP(16'h0935,4);
TASK_PP(16'h0936,4);
TASK_PP(16'h0937,4);
TASK_PP(16'h0938,4);
TASK_PP(16'h0939,4);
TASK_PP(16'h093A,4);
TASK_PP(16'h093B,4);
TASK_PP(16'h093C,4);
TASK_PP(16'h093D,4);
TASK_PP(16'h093E,4);
TASK_PP(16'h093F,4);
TASK_PP(16'h0940,4);
TASK_PP(16'h0941,4);
TASK_PP(16'h0942,4);
TASK_PP(16'h0943,4);
TASK_PP(16'h0944,4);
TASK_PP(16'h0945,4);
TASK_PP(16'h0946,4);
TASK_PP(16'h0947,4);
TASK_PP(16'h0948,4);
TASK_PP(16'h0949,4);
TASK_PP(16'h094A,4);
TASK_PP(16'h094B,4);
TASK_PP(16'h094C,4);
TASK_PP(16'h094D,4);
TASK_PP(16'h094E,4);
TASK_PP(16'h094F,4);
TASK_PP(16'h0950,4);
TASK_PP(16'h0951,4);
TASK_PP(16'h0952,4);
TASK_PP(16'h0953,4);
TASK_PP(16'h0954,4);
TASK_PP(16'h0955,4);
TASK_PP(16'h0956,4);
TASK_PP(16'h0957,4);
TASK_PP(16'h0958,4);
TASK_PP(16'h0959,4);
TASK_PP(16'h095A,4);
TASK_PP(16'h095B,4);
TASK_PP(16'h095C,4);
TASK_PP(16'h095D,4);
TASK_PP(16'h095E,4);
TASK_PP(16'h095F,4);
TASK_PP(16'h0960,4);
TASK_PP(16'h0961,4);
TASK_PP(16'h0962,4);
TASK_PP(16'h0963,4);
TASK_PP(16'h0964,4);
TASK_PP(16'h0965,4);
TASK_PP(16'h0966,4);
TASK_PP(16'h0967,4);
TASK_PP(16'h0968,4);
TASK_PP(16'h0969,4);
TASK_PP(16'h096A,4);
TASK_PP(16'h096B,4);
TASK_PP(16'h096C,4);
TASK_PP(16'h096D,4);
TASK_PP(16'h096E,4);
TASK_PP(16'h096F,4);
TASK_PP(16'h0970,4);
TASK_PP(16'h0971,4);
TASK_PP(16'h0972,4);
TASK_PP(16'h0973,4);
TASK_PP(16'h0974,4);
TASK_PP(16'h0975,4);
TASK_PP(16'h0976,4);
TASK_PP(16'h0977,4);
TASK_PP(16'h0978,4);
TASK_PP(16'h0979,4);
TASK_PP(16'h097A,4);
TASK_PP(16'h097B,4);
TASK_PP(16'h097C,4);
TASK_PP(16'h097D,4);
TASK_PP(16'h097E,4);
TASK_PP(16'h097F,4);
TASK_PP(16'h0980,4);
TASK_PP(16'h0981,4);
TASK_PP(16'h0982,4);
TASK_PP(16'h0983,4);
TASK_PP(16'h0984,4);
TASK_PP(16'h0985,4);
TASK_PP(16'h0986,4);
TASK_PP(16'h0987,4);
TASK_PP(16'h0988,4);
TASK_PP(16'h0989,4);
TASK_PP(16'h098A,4);
TASK_PP(16'h098B,4);
TASK_PP(16'h098C,4);
TASK_PP(16'h098D,4);
TASK_PP(16'h098E,4);
TASK_PP(16'h098F,4);
TASK_PP(16'h0990,4);
TASK_PP(16'h0991,4);
TASK_PP(16'h0992,4);
TASK_PP(16'h0993,4);
TASK_PP(16'h0994,4);
TASK_PP(16'h0995,4);
TASK_PP(16'h0996,4);
TASK_PP(16'h0997,4);
TASK_PP(16'h0998,4);
TASK_PP(16'h0999,4);
TASK_PP(16'h099A,4);
TASK_PP(16'h099B,4);
TASK_PP(16'h099C,4);
TASK_PP(16'h099D,4);
TASK_PP(16'h099E,4);
TASK_PP(16'h099F,4);
TASK_PP(16'h09A0,4);
TASK_PP(16'h09A1,4);
TASK_PP(16'h09A2,4);
TASK_PP(16'h09A3,4);
TASK_PP(16'h09A4,4);
TASK_PP(16'h09A5,4);
TASK_PP(16'h09A6,4);
TASK_PP(16'h09A7,4);
TASK_PP(16'h09A8,4);
TASK_PP(16'h09A9,4);
TASK_PP(16'h09AA,4);
TASK_PP(16'h09AB,4);
TASK_PP(16'h09AC,4);
TASK_PP(16'h09AD,4);
TASK_PP(16'h09AE,4);
TASK_PP(16'h09AF,4);
TASK_PP(16'h09B0,4);
TASK_PP(16'h09B1,4);
TASK_PP(16'h09B2,4);
TASK_PP(16'h09B3,4);
TASK_PP(16'h09B4,4);
TASK_PP(16'h09B5,4);
TASK_PP(16'h09B6,4);
TASK_PP(16'h09B7,4);
TASK_PP(16'h09B8,4);
TASK_PP(16'h09B9,4);
TASK_PP(16'h09BA,4);
TASK_PP(16'h09BB,4);
TASK_PP(16'h09BC,4);
TASK_PP(16'h09BD,4);
TASK_PP(16'h09BE,4);
TASK_PP(16'h09BF,4);
TASK_PP(16'h09C0,4);
TASK_PP(16'h09C1,4);
TASK_PP(16'h09C2,4);
TASK_PP(16'h09C3,4);
TASK_PP(16'h09C4,4);
TASK_PP(16'h09C5,4);
TASK_PP(16'h09C6,4);
TASK_PP(16'h09C7,4);
TASK_PP(16'h09C8,4);
TASK_PP(16'h09C9,4);
TASK_PP(16'h09CA,4);
TASK_PP(16'h09CB,4);
TASK_PP(16'h09CC,4);
TASK_PP(16'h09CD,4);
TASK_PP(16'h09CE,4);
TASK_PP(16'h09CF,4);
TASK_PP(16'h09D0,4);
TASK_PP(16'h09D1,4);
TASK_PP(16'h09D2,4);
TASK_PP(16'h09D3,4);
TASK_PP(16'h09D4,4);
TASK_PP(16'h09D5,4);
TASK_PP(16'h09D6,4);
TASK_PP(16'h09D7,4);
TASK_PP(16'h09D8,4);
TASK_PP(16'h09D9,4);
TASK_PP(16'h09DA,4);
TASK_PP(16'h09DB,4);
TASK_PP(16'h09DC,4);
TASK_PP(16'h09DD,4);
TASK_PP(16'h09DE,4);
TASK_PP(16'h09DF,4);
TASK_PP(16'h09E0,4);
TASK_PP(16'h09E1,4);
TASK_PP(16'h09E2,4);
TASK_PP(16'h09E3,4);
TASK_PP(16'h09E4,4);
TASK_PP(16'h09E5,4);
TASK_PP(16'h09E6,4);
TASK_PP(16'h09E7,4);
TASK_PP(16'h09E8,4);
TASK_PP(16'h09E9,4);
TASK_PP(16'h09EA,4);
TASK_PP(16'h09EB,4);
TASK_PP(16'h09EC,4);
TASK_PP(16'h09ED,4);
TASK_PP(16'h09EE,4);
TASK_PP(16'h09EF,4);
TASK_PP(16'h09F0,4);
TASK_PP(16'h09F1,4);
TASK_PP(16'h09F2,4);
TASK_PP(16'h09F3,4);
TASK_PP(16'h09F4,4);
TASK_PP(16'h09F5,4);
TASK_PP(16'h09F6,4);
TASK_PP(16'h09F7,4);
TASK_PP(16'h09F8,4);
TASK_PP(16'h09F9,4);
TASK_PP(16'h09FA,4);
TASK_PP(16'h09FB,4);
TASK_PP(16'h09FC,4);
TASK_PP(16'h09FD,4);
TASK_PP(16'h09FE,4);
TASK_PP(16'h09FF,4);
TASK_PP(16'h0A00,4);
TASK_PP(16'h0A01,4);
TASK_PP(16'h0A02,4);
TASK_PP(16'h0A03,4);
TASK_PP(16'h0A04,4);
TASK_PP(16'h0A05,4);
TASK_PP(16'h0A06,4);
TASK_PP(16'h0A07,4);
TASK_PP(16'h0A08,4);
TASK_PP(16'h0A09,4);
TASK_PP(16'h0A0A,4);
TASK_PP(16'h0A0B,4);
TASK_PP(16'h0A0C,4);
TASK_PP(16'h0A0D,4);
TASK_PP(16'h0A0E,4);
TASK_PP(16'h0A0F,4);
TASK_PP(16'h0A10,4);
TASK_PP(16'h0A11,4);
TASK_PP(16'h0A12,4);
TASK_PP(16'h0A13,4);
TASK_PP(16'h0A14,4);
TASK_PP(16'h0A15,4);
TASK_PP(16'h0A16,4);
TASK_PP(16'h0A17,4);
TASK_PP(16'h0A18,4);
TASK_PP(16'h0A19,4);
TASK_PP(16'h0A1A,4);
TASK_PP(16'h0A1B,4);
TASK_PP(16'h0A1C,4);
TASK_PP(16'h0A1D,4);
TASK_PP(16'h0A1E,4);
TASK_PP(16'h0A1F,4);
TASK_PP(16'h0A20,4);
TASK_PP(16'h0A21,4);
TASK_PP(16'h0A22,4);
TASK_PP(16'h0A23,4);
TASK_PP(16'h0A24,4);
TASK_PP(16'h0A25,4);
TASK_PP(16'h0A26,4);
TASK_PP(16'h0A27,4);
TASK_PP(16'h0A28,4);
TASK_PP(16'h0A29,4);
TASK_PP(16'h0A2A,4);
TASK_PP(16'h0A2B,4);
TASK_PP(16'h0A2C,4);
TASK_PP(16'h0A2D,4);
TASK_PP(16'h0A2E,4);
TASK_PP(16'h0A2F,4);
TASK_PP(16'h0A30,4);
TASK_PP(16'h0A31,4);
TASK_PP(16'h0A32,4);
TASK_PP(16'h0A33,4);
TASK_PP(16'h0A34,4);
TASK_PP(16'h0A35,4);
TASK_PP(16'h0A36,4);
TASK_PP(16'h0A37,4);
TASK_PP(16'h0A38,4);
TASK_PP(16'h0A39,4);
TASK_PP(16'h0A3A,4);
TASK_PP(16'h0A3B,4);
TASK_PP(16'h0A3C,4);
TASK_PP(16'h0A3D,4);
TASK_PP(16'h0A3E,4);
TASK_PP(16'h0A3F,4);
TASK_PP(16'h0A40,4);
TASK_PP(16'h0A41,4);
TASK_PP(16'h0A42,4);
TASK_PP(16'h0A43,4);
TASK_PP(16'h0A44,4);
TASK_PP(16'h0A45,4);
TASK_PP(16'h0A46,4);
TASK_PP(16'h0A47,4);
TASK_PP(16'h0A48,4);
TASK_PP(16'h0A49,4);
TASK_PP(16'h0A4A,4);
TASK_PP(16'h0A4B,4);
TASK_PP(16'h0A4C,4);
TASK_PP(16'h0A4D,4);
TASK_PP(16'h0A4E,4);
TASK_PP(16'h0A4F,4);
TASK_PP(16'h0A50,4);
TASK_PP(16'h0A51,4);
TASK_PP(16'h0A52,4);
TASK_PP(16'h0A53,4);
TASK_PP(16'h0A54,4);
TASK_PP(16'h0A55,4);
TASK_PP(16'h0A56,4);
TASK_PP(16'h0A57,4);
TASK_PP(16'h0A58,4);
TASK_PP(16'h0A59,4);
TASK_PP(16'h0A5A,4);
TASK_PP(16'h0A5B,4);
TASK_PP(16'h0A5C,4);
TASK_PP(16'h0A5D,4);
TASK_PP(16'h0A5E,4);
TASK_PP(16'h0A5F,4);
TASK_PP(16'h0A60,4);
TASK_PP(16'h0A61,4);
TASK_PP(16'h0A62,4);
TASK_PP(16'h0A63,4);
TASK_PP(16'h0A64,4);
TASK_PP(16'h0A65,4);
TASK_PP(16'h0A66,4);
TASK_PP(16'h0A67,4);
TASK_PP(16'h0A68,4);
TASK_PP(16'h0A69,4);
TASK_PP(16'h0A6A,4);
TASK_PP(16'h0A6B,4);
TASK_PP(16'h0A6C,4);
TASK_PP(16'h0A6D,4);
TASK_PP(16'h0A6E,4);
TASK_PP(16'h0A6F,4);
TASK_PP(16'h0A70,4);
TASK_PP(16'h0A71,4);
TASK_PP(16'h0A72,4);
TASK_PP(16'h0A73,4);
TASK_PP(16'h0A74,4);
TASK_PP(16'h0A75,4);
TASK_PP(16'h0A76,4);
TASK_PP(16'h0A77,4);
TASK_PP(16'h0A78,4);
TASK_PP(16'h0A79,4);
TASK_PP(16'h0A7A,4);
TASK_PP(16'h0A7B,4);
TASK_PP(16'h0A7C,4);
TASK_PP(16'h0A7D,4);
TASK_PP(16'h0A7E,4);
TASK_PP(16'h0A7F,4);
TASK_PP(16'h0A80,4);
TASK_PP(16'h0A81,4);
TASK_PP(16'h0A82,4);
TASK_PP(16'h0A83,4);
TASK_PP(16'h0A84,4);
TASK_PP(16'h0A85,4);
TASK_PP(16'h0A86,4);
TASK_PP(16'h0A87,4);
TASK_PP(16'h0A88,4);
TASK_PP(16'h0A89,4);
TASK_PP(16'h0A8A,4);
TASK_PP(16'h0A8B,4);
TASK_PP(16'h0A8C,4);
TASK_PP(16'h0A8D,4);
TASK_PP(16'h0A8E,4);
TASK_PP(16'h0A8F,4);
TASK_PP(16'h0A90,4);
TASK_PP(16'h0A91,4);
TASK_PP(16'h0A92,4);
TASK_PP(16'h0A93,4);
TASK_PP(16'h0A94,4);
TASK_PP(16'h0A95,4);
TASK_PP(16'h0A96,4);
TASK_PP(16'h0A97,4);
TASK_PP(16'h0A98,4);
TASK_PP(16'h0A99,4);
TASK_PP(16'h0A9A,4);
TASK_PP(16'h0A9B,4);
TASK_PP(16'h0A9C,4);
TASK_PP(16'h0A9D,4);
TASK_PP(16'h0A9E,4);
TASK_PP(16'h0A9F,4);
TASK_PP(16'h0AA0,4);
TASK_PP(16'h0AA1,4);
TASK_PP(16'h0AA2,4);
TASK_PP(16'h0AA3,4);
TASK_PP(16'h0AA4,4);
TASK_PP(16'h0AA5,4);
TASK_PP(16'h0AA6,4);
TASK_PP(16'h0AA7,4);
TASK_PP(16'h0AA8,4);
TASK_PP(16'h0AA9,4);
TASK_PP(16'h0AAA,4);
TASK_PP(16'h0AAB,4);
TASK_PP(16'h0AAC,4);
TASK_PP(16'h0AAD,4);
TASK_PP(16'h0AAE,4);
TASK_PP(16'h0AAF,4);
TASK_PP(16'h0AB0,4);
TASK_PP(16'h0AB1,4);
TASK_PP(16'h0AB2,4);
TASK_PP(16'h0AB3,4);
TASK_PP(16'h0AB4,4);
TASK_PP(16'h0AB5,4);
TASK_PP(16'h0AB6,4);
TASK_PP(16'h0AB7,4);
TASK_PP(16'h0AB8,4);
TASK_PP(16'h0AB9,4);
TASK_PP(16'h0ABA,4);
TASK_PP(16'h0ABB,4);
TASK_PP(16'h0ABC,4);
TASK_PP(16'h0ABD,4);
TASK_PP(16'h0ABE,4);
TASK_PP(16'h0ABF,4);
TASK_PP(16'h0AC0,4);
TASK_PP(16'h0AC1,4);
TASK_PP(16'h0AC2,4);
TASK_PP(16'h0AC3,4);
TASK_PP(16'h0AC4,4);
TASK_PP(16'h0AC5,4);
TASK_PP(16'h0AC6,4);
TASK_PP(16'h0AC7,4);
TASK_PP(16'h0AC8,4);
TASK_PP(16'h0AC9,4);
TASK_PP(16'h0ACA,4);
TASK_PP(16'h0ACB,4);
TASK_PP(16'h0ACC,4);
TASK_PP(16'h0ACD,4);
TASK_PP(16'h0ACE,4);
TASK_PP(16'h0ACF,4);
TASK_PP(16'h0AD0,4);
TASK_PP(16'h0AD1,4);
TASK_PP(16'h0AD2,4);
TASK_PP(16'h0AD3,4);
TASK_PP(16'h0AD4,4);
TASK_PP(16'h0AD5,4);
TASK_PP(16'h0AD6,4);
TASK_PP(16'h0AD7,4);
TASK_PP(16'h0AD8,4);
TASK_PP(16'h0AD9,4);
TASK_PP(16'h0ADA,4);
TASK_PP(16'h0ADB,4);
TASK_PP(16'h0ADC,4);
TASK_PP(16'h0ADD,4);
TASK_PP(16'h0ADE,4);
TASK_PP(16'h0ADF,4);
TASK_PP(16'h0AE0,4);
TASK_PP(16'h0AE1,4);
TASK_PP(16'h0AE2,4);
TASK_PP(16'h0AE3,4);
TASK_PP(16'h0AE4,4);
TASK_PP(16'h0AE5,4);
TASK_PP(16'h0AE6,4);
TASK_PP(16'h0AE7,4);
TASK_PP(16'h0AE8,4);
TASK_PP(16'h0AE9,4);
TASK_PP(16'h0AEA,4);
TASK_PP(16'h0AEB,4);
TASK_PP(16'h0AEC,4);
TASK_PP(16'h0AED,4);
TASK_PP(16'h0AEE,4);
TASK_PP(16'h0AEF,4);
TASK_PP(16'h0AF0,4);
TASK_PP(16'h0AF1,4);
TASK_PP(16'h0AF2,4);
TASK_PP(16'h0AF3,4);
TASK_PP(16'h0AF4,4);
TASK_PP(16'h0AF5,4);
TASK_PP(16'h0AF6,4);
TASK_PP(16'h0AF7,4);
TASK_PP(16'h0AF8,4);
TASK_PP(16'h0AF9,4);
TASK_PP(16'h0AFA,4);
TASK_PP(16'h0AFB,4);
TASK_PP(16'h0AFC,4);
TASK_PP(16'h0AFD,4);
TASK_PP(16'h0AFE,4);
TASK_PP(16'h0AFF,4);
TASK_PP(16'h0B00,4);
TASK_PP(16'h0B01,4);
TASK_PP(16'h0B02,4);
TASK_PP(16'h0B03,4);
TASK_PP(16'h0B04,4);
TASK_PP(16'h0B05,4);
TASK_PP(16'h0B06,4);
TASK_PP(16'h0B07,4);
TASK_PP(16'h0B08,4);
TASK_PP(16'h0B09,4);
TASK_PP(16'h0B0A,4);
TASK_PP(16'h0B0B,4);
TASK_PP(16'h0B0C,4);
TASK_PP(16'h0B0D,4);
TASK_PP(16'h0B0E,4);
TASK_PP(16'h0B0F,4);
TASK_PP(16'h0B10,4);
TASK_PP(16'h0B11,4);
TASK_PP(16'h0B12,4);
TASK_PP(16'h0B13,4);
TASK_PP(16'h0B14,4);
TASK_PP(16'h0B15,4);
TASK_PP(16'h0B16,4);
TASK_PP(16'h0B17,4);
TASK_PP(16'h0B18,4);
TASK_PP(16'h0B19,4);
TASK_PP(16'h0B1A,4);
TASK_PP(16'h0B1B,4);
TASK_PP(16'h0B1C,4);
TASK_PP(16'h0B1D,4);
TASK_PP(16'h0B1E,4);
TASK_PP(16'h0B1F,4);
TASK_PP(16'h0B20,4);
TASK_PP(16'h0B21,4);
TASK_PP(16'h0B22,4);
TASK_PP(16'h0B23,4);
TASK_PP(16'h0B24,4);
TASK_PP(16'h0B25,4);
TASK_PP(16'h0B26,4);
TASK_PP(16'h0B27,4);
TASK_PP(16'h0B28,4);
TASK_PP(16'h0B29,4);
TASK_PP(16'h0B2A,4);
TASK_PP(16'h0B2B,4);
TASK_PP(16'h0B2C,4);
TASK_PP(16'h0B2D,4);
TASK_PP(16'h0B2E,4);
TASK_PP(16'h0B2F,4);
TASK_PP(16'h0B30,4);
TASK_PP(16'h0B31,4);
TASK_PP(16'h0B32,4);
TASK_PP(16'h0B33,4);
TASK_PP(16'h0B34,4);
TASK_PP(16'h0B35,4);
TASK_PP(16'h0B36,4);
TASK_PP(16'h0B37,4);
TASK_PP(16'h0B38,4);
TASK_PP(16'h0B39,4);
TASK_PP(16'h0B3A,4);
TASK_PP(16'h0B3B,4);
TASK_PP(16'h0B3C,4);
TASK_PP(16'h0B3D,4);
TASK_PP(16'h0B3E,4);
TASK_PP(16'h0B3F,4);
TASK_PP(16'h0B40,4);
TASK_PP(16'h0B41,4);
TASK_PP(16'h0B42,4);
TASK_PP(16'h0B43,4);
TASK_PP(16'h0B44,4);
TASK_PP(16'h0B45,4);
TASK_PP(16'h0B46,4);
TASK_PP(16'h0B47,4);
TASK_PP(16'h0B48,4);
TASK_PP(16'h0B49,4);
TASK_PP(16'h0B4A,4);
TASK_PP(16'h0B4B,4);
TASK_PP(16'h0B4C,4);
TASK_PP(16'h0B4D,4);
TASK_PP(16'h0B4E,4);
TASK_PP(16'h0B4F,4);
TASK_PP(16'h0B50,4);
TASK_PP(16'h0B51,4);
TASK_PP(16'h0B52,4);
TASK_PP(16'h0B53,4);
TASK_PP(16'h0B54,4);
TASK_PP(16'h0B55,4);
TASK_PP(16'h0B56,4);
TASK_PP(16'h0B57,4);
TASK_PP(16'h0B58,4);
TASK_PP(16'h0B59,4);
TASK_PP(16'h0B5A,4);
TASK_PP(16'h0B5B,4);
TASK_PP(16'h0B5C,4);
TASK_PP(16'h0B5D,4);
TASK_PP(16'h0B5E,4);
TASK_PP(16'h0B5F,4);
TASK_PP(16'h0B60,4);
TASK_PP(16'h0B61,4);
TASK_PP(16'h0B62,4);
TASK_PP(16'h0B63,4);
TASK_PP(16'h0B64,4);
TASK_PP(16'h0B65,4);
TASK_PP(16'h0B66,4);
TASK_PP(16'h0B67,4);
TASK_PP(16'h0B68,4);
TASK_PP(16'h0B69,4);
TASK_PP(16'h0B6A,4);
TASK_PP(16'h0B6B,4);
TASK_PP(16'h0B6C,4);
TASK_PP(16'h0B6D,4);
TASK_PP(16'h0B6E,4);
TASK_PP(16'h0B6F,4);
TASK_PP(16'h0B70,4);
TASK_PP(16'h0B71,4);
TASK_PP(16'h0B72,4);
TASK_PP(16'h0B73,4);
TASK_PP(16'h0B74,4);
TASK_PP(16'h0B75,4);
TASK_PP(16'h0B76,4);
TASK_PP(16'h0B77,4);
TASK_PP(16'h0B78,4);
TASK_PP(16'h0B79,4);
TASK_PP(16'h0B7A,4);
TASK_PP(16'h0B7B,4);
TASK_PP(16'h0B7C,4);
TASK_PP(16'h0B7D,4);
TASK_PP(16'h0B7E,4);
TASK_PP(16'h0B7F,4);
TASK_PP(16'h0B80,4);
TASK_PP(16'h0B81,4);
TASK_PP(16'h0B82,4);
TASK_PP(16'h0B83,4);
TASK_PP(16'h0B84,4);
TASK_PP(16'h0B85,4);
TASK_PP(16'h0B86,4);
TASK_PP(16'h0B87,4);
TASK_PP(16'h0B88,4);
TASK_PP(16'h0B89,4);
TASK_PP(16'h0B8A,4);
TASK_PP(16'h0B8B,4);
TASK_PP(16'h0B8C,4);
TASK_PP(16'h0B8D,4);
TASK_PP(16'h0B8E,4);
TASK_PP(16'h0B8F,4);
TASK_PP(16'h0B90,4);
TASK_PP(16'h0B91,4);
TASK_PP(16'h0B92,4);
TASK_PP(16'h0B93,4);
TASK_PP(16'h0B94,4);
TASK_PP(16'h0B95,4);
TASK_PP(16'h0B96,4);
TASK_PP(16'h0B97,4);
TASK_PP(16'h0B98,4);
TASK_PP(16'h0B99,4);
TASK_PP(16'h0B9A,4);
TASK_PP(16'h0B9B,4);
TASK_PP(16'h0B9C,4);
TASK_PP(16'h0B9D,4);
TASK_PP(16'h0B9E,4);
TASK_PP(16'h0B9F,4);
TASK_PP(16'h0BA0,4);
TASK_PP(16'h0BA1,4);
TASK_PP(16'h0BA2,4);
TASK_PP(16'h0BA3,4);
TASK_PP(16'h0BA4,4);
TASK_PP(16'h0BA5,4);
TASK_PP(16'h0BA6,4);
TASK_PP(16'h0BA7,4);
TASK_PP(16'h0BA8,4);
TASK_PP(16'h0BA9,4);
TASK_PP(16'h0BAA,4);
TASK_PP(16'h0BAB,4);
TASK_PP(16'h0BAC,4);
TASK_PP(16'h0BAD,4);
TASK_PP(16'h0BAE,4);
TASK_PP(16'h0BAF,4);
TASK_PP(16'h0BB0,4);
TASK_PP(16'h0BB1,4);
TASK_PP(16'h0BB2,4);
TASK_PP(16'h0BB3,4);
TASK_PP(16'h0BB4,4);
TASK_PP(16'h0BB5,4);
TASK_PP(16'h0BB6,4);
TASK_PP(16'h0BB7,4);
TASK_PP(16'h0BB8,4);
TASK_PP(16'h0BB9,4);
TASK_PP(16'h0BBA,4);
TASK_PP(16'h0BBB,4);
TASK_PP(16'h0BBC,4);
TASK_PP(16'h0BBD,4);
TASK_PP(16'h0BBE,4);
TASK_PP(16'h0BBF,4);
TASK_PP(16'h0BC0,4);
TASK_PP(16'h0BC1,4);
TASK_PP(16'h0BC2,4);
TASK_PP(16'h0BC3,4);
TASK_PP(16'h0BC4,4);
TASK_PP(16'h0BC5,4);
TASK_PP(16'h0BC6,4);
TASK_PP(16'h0BC7,4);
TASK_PP(16'h0BC8,4);
TASK_PP(16'h0BC9,4);
TASK_PP(16'h0BCA,4);
TASK_PP(16'h0BCB,4);
TASK_PP(16'h0BCC,4);
TASK_PP(16'h0BCD,4);
TASK_PP(16'h0BCE,4);
TASK_PP(16'h0BCF,4);
TASK_PP(16'h0BD0,4);
TASK_PP(16'h0BD1,4);
TASK_PP(16'h0BD2,4);
TASK_PP(16'h0BD3,4);
TASK_PP(16'h0BD4,4);
TASK_PP(16'h0BD5,4);
TASK_PP(16'h0BD6,4);
TASK_PP(16'h0BD7,4);
TASK_PP(16'h0BD8,4);
TASK_PP(16'h0BD9,4);
TASK_PP(16'h0BDA,4);
TASK_PP(16'h0BDB,4);
TASK_PP(16'h0BDC,4);
TASK_PP(16'h0BDD,4);
TASK_PP(16'h0BDE,4);
TASK_PP(16'h0BDF,4);
TASK_PP(16'h0BE0,4);
TASK_PP(16'h0BE1,4);
TASK_PP(16'h0BE2,4);
TASK_PP(16'h0BE3,4);
TASK_PP(16'h0BE4,4);
TASK_PP(16'h0BE5,4);
TASK_PP(16'h0BE6,4);
TASK_PP(16'h0BE7,4);
TASK_PP(16'h0BE8,4);
TASK_PP(16'h0BE9,4);
TASK_PP(16'h0BEA,4);
TASK_PP(16'h0BEB,4);
TASK_PP(16'h0BEC,4);
TASK_PP(16'h0BED,4);
TASK_PP(16'h0BEE,4);
TASK_PP(16'h0BEF,4);
TASK_PP(16'h0BF0,4);
TASK_PP(16'h0BF1,4);
TASK_PP(16'h0BF2,4);
TASK_PP(16'h0BF3,4);
TASK_PP(16'h0BF4,4);
TASK_PP(16'h0BF5,4);
TASK_PP(16'h0BF6,4);
TASK_PP(16'h0BF7,4);
TASK_PP(16'h0BF8,4);
TASK_PP(16'h0BF9,4);
TASK_PP(16'h0BFA,4);
TASK_PP(16'h0BFB,4);
TASK_PP(16'h0BFC,4);
TASK_PP(16'h0BFD,4);
TASK_PP(16'h0BFE,4);
TASK_PP(16'h0BFF,4);
TASK_PP(16'h0C00,4);
TASK_PP(16'h0C01,4);
TASK_PP(16'h0C02,4);
TASK_PP(16'h0C03,4);
TASK_PP(16'h0C04,4);
TASK_PP(16'h0C05,4);
TASK_PP(16'h0C06,4);
TASK_PP(16'h0C07,4);
TASK_PP(16'h0C08,4);
TASK_PP(16'h0C09,4);
TASK_PP(16'h0C0A,4);
TASK_PP(16'h0C0B,4);
TASK_PP(16'h0C0C,4);
TASK_PP(16'h0C0D,4);
TASK_PP(16'h0C0E,4);
TASK_PP(16'h0C0F,4);
TASK_PP(16'h0C10,4);
TASK_PP(16'h0C11,4);
TASK_PP(16'h0C12,4);
TASK_PP(16'h0C13,4);
TASK_PP(16'h0C14,4);
TASK_PP(16'h0C15,4);
TASK_PP(16'h0C16,4);
TASK_PP(16'h0C17,4);
TASK_PP(16'h0C18,4);
TASK_PP(16'h0C19,4);
TASK_PP(16'h0C1A,4);
TASK_PP(16'h0C1B,4);
TASK_PP(16'h0C1C,4);
TASK_PP(16'h0C1D,4);
TASK_PP(16'h0C1E,4);
TASK_PP(16'h0C1F,4);
TASK_PP(16'h0C20,4);
TASK_PP(16'h0C21,4);
TASK_PP(16'h0C22,4);
TASK_PP(16'h0C23,4);
TASK_PP(16'h0C24,4);
TASK_PP(16'h0C25,4);
TASK_PP(16'h0C26,4);
TASK_PP(16'h0C27,4);
TASK_PP(16'h0C28,4);
TASK_PP(16'h0C29,4);
TASK_PP(16'h0C2A,4);
TASK_PP(16'h0C2B,4);
TASK_PP(16'h0C2C,4);
TASK_PP(16'h0C2D,4);
TASK_PP(16'h0C2E,4);
TASK_PP(16'h0C2F,4);
TASK_PP(16'h0C30,4);
TASK_PP(16'h0C31,4);
TASK_PP(16'h0C32,4);
TASK_PP(16'h0C33,4);
TASK_PP(16'h0C34,4);
TASK_PP(16'h0C35,4);
TASK_PP(16'h0C36,4);
TASK_PP(16'h0C37,4);
TASK_PP(16'h0C38,4);
TASK_PP(16'h0C39,4);
TASK_PP(16'h0C3A,4);
TASK_PP(16'h0C3B,4);
TASK_PP(16'h0C3C,4);
TASK_PP(16'h0C3D,4);
TASK_PP(16'h0C3E,4);
TASK_PP(16'h0C3F,4);
TASK_PP(16'h0C40,4);
TASK_PP(16'h0C41,4);
TASK_PP(16'h0C42,4);
TASK_PP(16'h0C43,4);
TASK_PP(16'h0C44,4);
TASK_PP(16'h0C45,4);
TASK_PP(16'h0C46,4);
TASK_PP(16'h0C47,4);
TASK_PP(16'h0C48,4);
TASK_PP(16'h0C49,4);
TASK_PP(16'h0C4A,4);
TASK_PP(16'h0C4B,4);
TASK_PP(16'h0C4C,4);
TASK_PP(16'h0C4D,4);
TASK_PP(16'h0C4E,4);
TASK_PP(16'h0C4F,4);
TASK_PP(16'h0C50,4);
TASK_PP(16'h0C51,4);
TASK_PP(16'h0C52,4);
TASK_PP(16'h0C53,4);
TASK_PP(16'h0C54,4);
TASK_PP(16'h0C55,4);
TASK_PP(16'h0C56,4);
TASK_PP(16'h0C57,4);
TASK_PP(16'h0C58,4);
TASK_PP(16'h0C59,4);
TASK_PP(16'h0C5A,4);
TASK_PP(16'h0C5B,4);
TASK_PP(16'h0C5C,4);
TASK_PP(16'h0C5D,4);
TASK_PP(16'h0C5E,4);
TASK_PP(16'h0C5F,4);
TASK_PP(16'h0C60,4);
TASK_PP(16'h0C61,4);
TASK_PP(16'h0C62,4);
TASK_PP(16'h0C63,4);
TASK_PP(16'h0C64,4);
TASK_PP(16'h0C65,4);
TASK_PP(16'h0C66,4);
TASK_PP(16'h0C67,4);
TASK_PP(16'h0C68,4);
TASK_PP(16'h0C69,4);
TASK_PP(16'h0C6A,4);
TASK_PP(16'h0C6B,4);
TASK_PP(16'h0C6C,4);
TASK_PP(16'h0C6D,4);
TASK_PP(16'h0C6E,4);
TASK_PP(16'h0C6F,4);
TASK_PP(16'h0C70,4);
TASK_PP(16'h0C71,4);
TASK_PP(16'h0C72,4);
TASK_PP(16'h0C73,4);
TASK_PP(16'h0C74,4);
TASK_PP(16'h0C75,4);
TASK_PP(16'h0C76,4);
TASK_PP(16'h0C77,4);
TASK_PP(16'h0C78,4);
TASK_PP(16'h0C79,4);
TASK_PP(16'h0C7A,4);
TASK_PP(16'h0C7B,4);
TASK_PP(16'h0C7C,4);
TASK_PP(16'h0C7D,4);
TASK_PP(16'h0C7E,4);
TASK_PP(16'h0C7F,4);
TASK_PP(16'h0C80,4);
TASK_PP(16'h0C81,4);
TASK_PP(16'h0C82,4);
TASK_PP(16'h0C83,4);
TASK_PP(16'h0C84,4);
TASK_PP(16'h0C85,4);
TASK_PP(16'h0C86,4);
TASK_PP(16'h0C87,4);
TASK_PP(16'h0C88,4);
TASK_PP(16'h0C89,4);
TASK_PP(16'h0C8A,4);
TASK_PP(16'h0C8B,4);
TASK_PP(16'h0C8C,4);
TASK_PP(16'h0C8D,4);
TASK_PP(16'h0C8E,4);
TASK_PP(16'h0C8F,4);
TASK_PP(16'h0C90,4);
TASK_PP(16'h0C91,4);
TASK_PP(16'h0C92,4);
TASK_PP(16'h0C93,4);
TASK_PP(16'h0C94,4);
TASK_PP(16'h0C95,4);
TASK_PP(16'h0C96,4);
TASK_PP(16'h0C97,4);
TASK_PP(16'h0C98,4);
TASK_PP(16'h0C99,4);
TASK_PP(16'h0C9A,4);
TASK_PP(16'h0C9B,4);
TASK_PP(16'h0C9C,4);
TASK_PP(16'h0C9D,4);
TASK_PP(16'h0C9E,4);
TASK_PP(16'h0C9F,4);
TASK_PP(16'h0CA0,4);
TASK_PP(16'h0CA1,4);
TASK_PP(16'h0CA2,4);
TASK_PP(16'h0CA3,4);
TASK_PP(16'h0CA4,4);
TASK_PP(16'h0CA5,4);
TASK_PP(16'h0CA6,4);
TASK_PP(16'h0CA7,4);
TASK_PP(16'h0CA8,4);
TASK_PP(16'h0CA9,4);
TASK_PP(16'h0CAA,4);
TASK_PP(16'h0CAB,4);
TASK_PP(16'h0CAC,4);
TASK_PP(16'h0CAD,4);
TASK_PP(16'h0CAE,4);
TASK_PP(16'h0CAF,4);
TASK_PP(16'h0CB0,4);
TASK_PP(16'h0CB1,4);
TASK_PP(16'h0CB2,4);
TASK_PP(16'h0CB3,4);
TASK_PP(16'h0CB4,4);
TASK_PP(16'h0CB5,4);
TASK_PP(16'h0CB6,4);
TASK_PP(16'h0CB7,4);
TASK_PP(16'h0CB8,4);
TASK_PP(16'h0CB9,4);
TASK_PP(16'h0CBA,4);
TASK_PP(16'h0CBB,4);
TASK_PP(16'h0CBC,4);
TASK_PP(16'h0CBD,4);
TASK_PP(16'h0CBE,4);
TASK_PP(16'h0CBF,4);
TASK_PP(16'h0CC0,4);
TASK_PP(16'h0CC1,4);
TASK_PP(16'h0CC2,4);
TASK_PP(16'h0CC3,4);
TASK_PP(16'h0CC4,4);
TASK_PP(16'h0CC5,4);
TASK_PP(16'h0CC6,4);
TASK_PP(16'h0CC7,4);
TASK_PP(16'h0CC8,4);
TASK_PP(16'h0CC9,4);
TASK_PP(16'h0CCA,4);
TASK_PP(16'h0CCB,4);
TASK_PP(16'h0CCC,4);
TASK_PP(16'h0CCD,4);
TASK_PP(16'h0CCE,4);
TASK_PP(16'h0CCF,4);
TASK_PP(16'h0CD0,4);
TASK_PP(16'h0CD1,4);
TASK_PP(16'h0CD2,4);
TASK_PP(16'h0CD3,4);
TASK_PP(16'h0CD4,4);
TASK_PP(16'h0CD5,4);
TASK_PP(16'h0CD6,4);
TASK_PP(16'h0CD7,4);
TASK_PP(16'h0CD8,4);
TASK_PP(16'h0CD9,4);
TASK_PP(16'h0CDA,4);
TASK_PP(16'h0CDB,4);
TASK_PP(16'h0CDC,4);
TASK_PP(16'h0CDD,4);
TASK_PP(16'h0CDE,4);
TASK_PP(16'h0CDF,4);
TASK_PP(16'h0CE0,4);
TASK_PP(16'h0CE1,4);
TASK_PP(16'h0CE2,4);
TASK_PP(16'h0CE3,4);
TASK_PP(16'h0CE4,4);
TASK_PP(16'h0CE5,4);
TASK_PP(16'h0CE6,4);
TASK_PP(16'h0CE7,4);
TASK_PP(16'h0CE8,4);
TASK_PP(16'h0CE9,4);
TASK_PP(16'h0CEA,4);
TASK_PP(16'h0CEB,4);
TASK_PP(16'h0CEC,4);
TASK_PP(16'h0CED,4);
TASK_PP(16'h0CEE,4);
TASK_PP(16'h0CEF,4);
TASK_PP(16'h0CF0,4);
TASK_PP(16'h0CF1,4);
TASK_PP(16'h0CF2,4);
TASK_PP(16'h0CF3,4);
TASK_PP(16'h0CF4,4);
TASK_PP(16'h0CF5,4);
TASK_PP(16'h0CF6,4);
TASK_PP(16'h0CF7,4);
TASK_PP(16'h0CF8,4);
TASK_PP(16'h0CF9,4);
TASK_PP(16'h0CFA,4);
TASK_PP(16'h0CFB,4);
TASK_PP(16'h0CFC,4);
TASK_PP(16'h0CFD,4);
TASK_PP(16'h0CFE,4);
TASK_PP(16'h0CFF,4);
TASK_PP(16'h0D00,4);
TASK_PP(16'h0D01,4);
TASK_PP(16'h0D02,4);
TASK_PP(16'h0D03,4);
TASK_PP(16'h0D04,4);
TASK_PP(16'h0D05,4);
TASK_PP(16'h0D06,4);
TASK_PP(16'h0D07,4);
TASK_PP(16'h0D08,4);
TASK_PP(16'h0D09,4);
TASK_PP(16'h0D0A,4);
TASK_PP(16'h0D0B,4);
TASK_PP(16'h0D0C,4);
TASK_PP(16'h0D0D,4);
TASK_PP(16'h0D0E,4);
TASK_PP(16'h0D0F,4);
TASK_PP(16'h0D10,4);
TASK_PP(16'h0D11,4);
TASK_PP(16'h0D12,4);
TASK_PP(16'h0D13,4);
TASK_PP(16'h0D14,4);
TASK_PP(16'h0D15,4);
TASK_PP(16'h0D16,4);
TASK_PP(16'h0D17,4);
TASK_PP(16'h0D18,4);
TASK_PP(16'h0D19,4);
TASK_PP(16'h0D1A,4);
TASK_PP(16'h0D1B,4);
TASK_PP(16'h0D1C,4);
TASK_PP(16'h0D1D,4);
TASK_PP(16'h0D1E,4);
TASK_PP(16'h0D1F,4);
TASK_PP(16'h0D20,4);
TASK_PP(16'h0D21,4);
TASK_PP(16'h0D22,4);
TASK_PP(16'h0D23,4);
TASK_PP(16'h0D24,4);
TASK_PP(16'h0D25,4);
TASK_PP(16'h0D26,4);
TASK_PP(16'h0D27,4);
TASK_PP(16'h0D28,4);
TASK_PP(16'h0D29,4);
TASK_PP(16'h0D2A,4);
TASK_PP(16'h0D2B,4);
TASK_PP(16'h0D2C,4);
TASK_PP(16'h0D2D,4);
TASK_PP(16'h0D2E,4);
TASK_PP(16'h0D2F,4);
TASK_PP(16'h0D30,4);
TASK_PP(16'h0D31,4);
TASK_PP(16'h0D32,4);
TASK_PP(16'h0D33,4);
TASK_PP(16'h0D34,4);
TASK_PP(16'h0D35,4);
TASK_PP(16'h0D36,4);
TASK_PP(16'h0D37,4);
TASK_PP(16'h0D38,4);
TASK_PP(16'h0D39,4);
TASK_PP(16'h0D3A,4);
TASK_PP(16'h0D3B,4);
TASK_PP(16'h0D3C,4);
TASK_PP(16'h0D3D,4);
TASK_PP(16'h0D3E,4);
TASK_PP(16'h0D3F,4);
TASK_PP(16'h0D40,4);
TASK_PP(16'h0D41,4);
TASK_PP(16'h0D42,4);
TASK_PP(16'h0D43,4);
TASK_PP(16'h0D44,4);
TASK_PP(16'h0D45,4);
TASK_PP(16'h0D46,4);
TASK_PP(16'h0D47,4);
TASK_PP(16'h0D48,4);
TASK_PP(16'h0D49,4);
TASK_PP(16'h0D4A,4);
TASK_PP(16'h0D4B,4);
TASK_PP(16'h0D4C,4);
TASK_PP(16'h0D4D,4);
TASK_PP(16'h0D4E,4);
TASK_PP(16'h0D4F,4);
TASK_PP(16'h0D50,4);
TASK_PP(16'h0D51,4);
TASK_PP(16'h0D52,4);
TASK_PP(16'h0D53,4);
TASK_PP(16'h0D54,4);
TASK_PP(16'h0D55,4);
TASK_PP(16'h0D56,4);
TASK_PP(16'h0D57,4);
TASK_PP(16'h0D58,4);
TASK_PP(16'h0D59,4);
TASK_PP(16'h0D5A,4);
TASK_PP(16'h0D5B,4);
TASK_PP(16'h0D5C,4);
TASK_PP(16'h0D5D,4);
TASK_PP(16'h0D5E,4);
TASK_PP(16'h0D5F,4);
TASK_PP(16'h0D60,4);
TASK_PP(16'h0D61,4);
TASK_PP(16'h0D62,4);
TASK_PP(16'h0D63,4);
TASK_PP(16'h0D64,4);
TASK_PP(16'h0D65,4);
TASK_PP(16'h0D66,4);
TASK_PP(16'h0D67,4);
TASK_PP(16'h0D68,4);
TASK_PP(16'h0D69,4);
TASK_PP(16'h0D6A,4);
TASK_PP(16'h0D6B,4);
TASK_PP(16'h0D6C,4);
TASK_PP(16'h0D6D,4);
TASK_PP(16'h0D6E,4);
TASK_PP(16'h0D6F,4);
TASK_PP(16'h0D70,4);
TASK_PP(16'h0D71,4);
TASK_PP(16'h0D72,4);
TASK_PP(16'h0D73,4);
TASK_PP(16'h0D74,4);
TASK_PP(16'h0D75,4);
TASK_PP(16'h0D76,4);
TASK_PP(16'h0D77,4);
TASK_PP(16'h0D78,4);
TASK_PP(16'h0D79,4);
TASK_PP(16'h0D7A,4);
TASK_PP(16'h0D7B,4);
TASK_PP(16'h0D7C,4);
TASK_PP(16'h0D7D,4);
TASK_PP(16'h0D7E,4);
TASK_PP(16'h0D7F,4);
TASK_PP(16'h0D80,4);
TASK_PP(16'h0D81,4);
TASK_PP(16'h0D82,4);
TASK_PP(16'h0D83,4);
TASK_PP(16'h0D84,4);
TASK_PP(16'h0D85,4);
TASK_PP(16'h0D86,4);
TASK_PP(16'h0D87,4);
TASK_PP(16'h0D88,4);
TASK_PP(16'h0D89,4);
TASK_PP(16'h0D8A,4);
TASK_PP(16'h0D8B,4);
TASK_PP(16'h0D8C,4);
TASK_PP(16'h0D8D,4);
TASK_PP(16'h0D8E,4);
TASK_PP(16'h0D8F,4);
TASK_PP(16'h0D90,4);
TASK_PP(16'h0D91,4);
TASK_PP(16'h0D92,4);
TASK_PP(16'h0D93,4);
TASK_PP(16'h0D94,4);
TASK_PP(16'h0D95,4);
TASK_PP(16'h0D96,4);
TASK_PP(16'h0D97,4);
TASK_PP(16'h0D98,4);
TASK_PP(16'h0D99,4);
TASK_PP(16'h0D9A,4);
TASK_PP(16'h0D9B,4);
TASK_PP(16'h0D9C,4);
TASK_PP(16'h0D9D,4);
TASK_PP(16'h0D9E,4);
TASK_PP(16'h0D9F,4);
TASK_PP(16'h0DA0,4);
TASK_PP(16'h0DA1,4);
TASK_PP(16'h0DA2,4);
TASK_PP(16'h0DA3,4);
TASK_PP(16'h0DA4,4);
TASK_PP(16'h0DA5,4);
TASK_PP(16'h0DA6,4);
TASK_PP(16'h0DA7,4);
TASK_PP(16'h0DA8,4);
TASK_PP(16'h0DA9,4);
TASK_PP(16'h0DAA,4);
TASK_PP(16'h0DAB,4);
TASK_PP(16'h0DAC,4);
TASK_PP(16'h0DAD,4);
TASK_PP(16'h0DAE,4);
TASK_PP(16'h0DAF,4);
TASK_PP(16'h0DB0,4);
TASK_PP(16'h0DB1,4);
TASK_PP(16'h0DB2,4);
TASK_PP(16'h0DB3,4);
TASK_PP(16'h0DB4,4);
TASK_PP(16'h0DB5,4);
TASK_PP(16'h0DB6,4);
TASK_PP(16'h0DB7,4);
TASK_PP(16'h0DB8,4);
TASK_PP(16'h0DB9,4);
TASK_PP(16'h0DBA,4);
TASK_PP(16'h0DBB,4);
TASK_PP(16'h0DBC,4);
TASK_PP(16'h0DBD,4);
TASK_PP(16'h0DBE,4);
TASK_PP(16'h0DBF,4);
TASK_PP(16'h0DC0,4);
TASK_PP(16'h0DC1,4);
TASK_PP(16'h0DC2,4);
TASK_PP(16'h0DC3,4);
TASK_PP(16'h0DC4,4);
TASK_PP(16'h0DC5,4);
TASK_PP(16'h0DC6,4);
TASK_PP(16'h0DC7,4);
TASK_PP(16'h0DC8,4);
TASK_PP(16'h0DC9,4);
TASK_PP(16'h0DCA,4);
TASK_PP(16'h0DCB,4);
TASK_PP(16'h0DCC,4);
TASK_PP(16'h0DCD,4);
TASK_PP(16'h0DCE,4);
TASK_PP(16'h0DCF,4);
TASK_PP(16'h0DD0,4);
TASK_PP(16'h0DD1,4);
TASK_PP(16'h0DD2,4);
TASK_PP(16'h0DD3,4);
TASK_PP(16'h0DD4,4);
TASK_PP(16'h0DD5,4);
TASK_PP(16'h0DD6,4);
TASK_PP(16'h0DD7,4);
TASK_PP(16'h0DD8,4);
TASK_PP(16'h0DD9,4);
TASK_PP(16'h0DDA,4);
TASK_PP(16'h0DDB,4);
TASK_PP(16'h0DDC,4);
TASK_PP(16'h0DDD,4);
TASK_PP(16'h0DDE,4);
TASK_PP(16'h0DDF,4);
TASK_PP(16'h0DE0,4);
TASK_PP(16'h0DE1,4);
TASK_PP(16'h0DE2,4);
TASK_PP(16'h0DE3,4);
TASK_PP(16'h0DE4,4);
TASK_PP(16'h0DE5,4);
TASK_PP(16'h0DE6,4);
TASK_PP(16'h0DE7,4);
TASK_PP(16'h0DE8,4);
TASK_PP(16'h0DE9,4);
TASK_PP(16'h0DEA,4);
TASK_PP(16'h0DEB,4);
TASK_PP(16'h0DEC,4);
TASK_PP(16'h0DED,4);
TASK_PP(16'h0DEE,4);
TASK_PP(16'h0DEF,4);
TASK_PP(16'h0DF0,4);
TASK_PP(16'h0DF1,4);
TASK_PP(16'h0DF2,4);
TASK_PP(16'h0DF3,4);
TASK_PP(16'h0DF4,4);
TASK_PP(16'h0DF5,4);
TASK_PP(16'h0DF6,4);
TASK_PP(16'h0DF7,4);
TASK_PP(16'h0DF8,4);
TASK_PP(16'h0DF9,4);
TASK_PP(16'h0DFA,4);
TASK_PP(16'h0DFB,4);
TASK_PP(16'h0DFC,4);
TASK_PP(16'h0DFD,4);
TASK_PP(16'h0DFE,4);
TASK_PP(16'h0DFF,4);
TASK_PP(16'h0E00,4);
TASK_PP(16'h0E01,4);
TASK_PP(16'h0E02,4);
TASK_PP(16'h0E03,4);
TASK_PP(16'h0E04,4);
TASK_PP(16'h0E05,4);
TASK_PP(16'h0E06,4);
TASK_PP(16'h0E07,4);
TASK_PP(16'h0E08,4);
TASK_PP(16'h0E09,4);
TASK_PP(16'h0E0A,4);
TASK_PP(16'h0E0B,4);
TASK_PP(16'h0E0C,4);
TASK_PP(16'h0E0D,4);
TASK_PP(16'h0E0E,4);
TASK_PP(16'h0E0F,4);
TASK_PP(16'h0E10,4);
TASK_PP(16'h0E11,4);
TASK_PP(16'h0E12,4);
TASK_PP(16'h0E13,4);
TASK_PP(16'h0E14,4);
TASK_PP(16'h0E15,4);
TASK_PP(16'h0E16,4);
TASK_PP(16'h0E17,4);
TASK_PP(16'h0E18,4);
TASK_PP(16'h0E19,4);
TASK_PP(16'h0E1A,4);
TASK_PP(16'h0E1B,4);
TASK_PP(16'h0E1C,4);
TASK_PP(16'h0E1D,4);
TASK_PP(16'h0E1E,4);
TASK_PP(16'h0E1F,4);
TASK_PP(16'h0E20,4);
TASK_PP(16'h0E21,4);
TASK_PP(16'h0E22,4);
TASK_PP(16'h0E23,4);
TASK_PP(16'h0E24,4);
TASK_PP(16'h0E25,4);
TASK_PP(16'h0E26,4);
TASK_PP(16'h0E27,4);
TASK_PP(16'h0E28,4);
TASK_PP(16'h0E29,4);
TASK_PP(16'h0E2A,4);
TASK_PP(16'h0E2B,4);
TASK_PP(16'h0E2C,4);
TASK_PP(16'h0E2D,4);
TASK_PP(16'h0E2E,4);
TASK_PP(16'h0E2F,4);
TASK_PP(16'h0E30,4);
TASK_PP(16'h0E31,4);
TASK_PP(16'h0E32,4);
TASK_PP(16'h0E33,4);
TASK_PP(16'h0E34,4);
TASK_PP(16'h0E35,4);
TASK_PP(16'h0E36,4);
TASK_PP(16'h0E37,4);
TASK_PP(16'h0E38,4);
TASK_PP(16'h0E39,4);
TASK_PP(16'h0E3A,4);
TASK_PP(16'h0E3B,4);
TASK_PP(16'h0E3C,4);
TASK_PP(16'h0E3D,4);
TASK_PP(16'h0E3E,4);
TASK_PP(16'h0E3F,4);
TASK_PP(16'h0E40,4);
TASK_PP(16'h0E41,4);
TASK_PP(16'h0E42,4);
TASK_PP(16'h0E43,4);
TASK_PP(16'h0E44,4);
TASK_PP(16'h0E45,4);
TASK_PP(16'h0E46,4);
TASK_PP(16'h0E47,4);
TASK_PP(16'h0E48,4);
TASK_PP(16'h0E49,4);
TASK_PP(16'h0E4A,4);
TASK_PP(16'h0E4B,4);
TASK_PP(16'h0E4C,4);
TASK_PP(16'h0E4D,4);
TASK_PP(16'h0E4E,4);
TASK_PP(16'h0E4F,4);
TASK_PP(16'h0E50,4);
TASK_PP(16'h0E51,4);
TASK_PP(16'h0E52,4);
TASK_PP(16'h0E53,4);
TASK_PP(16'h0E54,4);
TASK_PP(16'h0E55,4);
TASK_PP(16'h0E56,4);
TASK_PP(16'h0E57,4);
TASK_PP(16'h0E58,4);
TASK_PP(16'h0E59,4);
TASK_PP(16'h0E5A,4);
TASK_PP(16'h0E5B,4);
TASK_PP(16'h0E5C,4);
TASK_PP(16'h0E5D,4);
TASK_PP(16'h0E5E,4);
TASK_PP(16'h0E5F,4);
TASK_PP(16'h0E60,4);
TASK_PP(16'h0E61,4);
TASK_PP(16'h0E62,4);
TASK_PP(16'h0E63,4);
TASK_PP(16'h0E64,4);
TASK_PP(16'h0E65,4);
TASK_PP(16'h0E66,4);
TASK_PP(16'h0E67,4);
TASK_PP(16'h0E68,4);
TASK_PP(16'h0E69,4);
TASK_PP(16'h0E6A,4);
TASK_PP(16'h0E6B,4);
TASK_PP(16'h0E6C,4);
TASK_PP(16'h0E6D,4);
TASK_PP(16'h0E6E,4);
TASK_PP(16'h0E6F,4);
TASK_PP(16'h0E70,4);
TASK_PP(16'h0E71,4);
TASK_PP(16'h0E72,4);
TASK_PP(16'h0E73,4);
TASK_PP(16'h0E74,4);
TASK_PP(16'h0E75,4);
TASK_PP(16'h0E76,4);
TASK_PP(16'h0E77,4);
TASK_PP(16'h0E78,4);
TASK_PP(16'h0E79,4);
TASK_PP(16'h0E7A,4);
TASK_PP(16'h0E7B,4);
TASK_PP(16'h0E7C,4);
TASK_PP(16'h0E7D,4);
TASK_PP(16'h0E7E,4);
TASK_PP(16'h0E7F,4);
TASK_PP(16'h0E80,4);
TASK_PP(16'h0E81,4);
TASK_PP(16'h0E82,4);
TASK_PP(16'h0E83,4);
TASK_PP(16'h0E84,4);
TASK_PP(16'h0E85,4);
TASK_PP(16'h0E86,4);
TASK_PP(16'h0E87,4);
TASK_PP(16'h0E88,4);
TASK_PP(16'h0E89,4);
TASK_PP(16'h0E8A,4);
TASK_PP(16'h0E8B,4);
TASK_PP(16'h0E8C,4);
TASK_PP(16'h0E8D,4);
TASK_PP(16'h0E8E,4);
TASK_PP(16'h0E8F,4);
TASK_PP(16'h0E90,4);
TASK_PP(16'h0E91,4);
TASK_PP(16'h0E92,4);
TASK_PP(16'h0E93,4);
TASK_PP(16'h0E94,4);
TASK_PP(16'h0E95,4);
TASK_PP(16'h0E96,4);
TASK_PP(16'h0E97,4);
TASK_PP(16'h0E98,4);
TASK_PP(16'h0E99,4);
TASK_PP(16'h0E9A,4);
TASK_PP(16'h0E9B,4);
TASK_PP(16'h0E9C,4);
TASK_PP(16'h0E9D,4);
TASK_PP(16'h0E9E,4);
TASK_PP(16'h0E9F,4);
TASK_PP(16'h0EA0,4);
TASK_PP(16'h0EA1,4);
TASK_PP(16'h0EA2,4);
TASK_PP(16'h0EA3,4);
TASK_PP(16'h0EA4,4);
TASK_PP(16'h0EA5,4);
TASK_PP(16'h0EA6,4);
TASK_PP(16'h0EA7,4);
TASK_PP(16'h0EA8,4);
TASK_PP(16'h0EA9,4);
TASK_PP(16'h0EAA,4);
TASK_PP(16'h0EAB,4);
TASK_PP(16'h0EAC,4);
TASK_PP(16'h0EAD,4);
TASK_PP(16'h0EAE,4);
TASK_PP(16'h0EAF,4);
TASK_PP(16'h0EB0,4);
TASK_PP(16'h0EB1,4);
TASK_PP(16'h0EB2,4);
TASK_PP(16'h0EB3,4);
TASK_PP(16'h0EB4,4);
TASK_PP(16'h0EB5,4);
TASK_PP(16'h0EB6,4);
TASK_PP(16'h0EB7,4);
TASK_PP(16'h0EB8,4);
TASK_PP(16'h0EB9,4);
TASK_PP(16'h0EBA,4);
TASK_PP(16'h0EBB,4);
TASK_PP(16'h0EBC,4);
TASK_PP(16'h0EBD,4);
TASK_PP(16'h0EBE,4);
TASK_PP(16'h0EBF,4);
TASK_PP(16'h0EC0,4);
TASK_PP(16'h0EC1,4);
TASK_PP(16'h0EC2,4);
TASK_PP(16'h0EC3,4);
TASK_PP(16'h0EC4,4);
TASK_PP(16'h0EC5,4);
TASK_PP(16'h0EC6,4);
TASK_PP(16'h0EC7,4);
TASK_PP(16'h0EC8,4);
TASK_PP(16'h0EC9,4);
TASK_PP(16'h0ECA,4);
TASK_PP(16'h0ECB,4);
TASK_PP(16'h0ECC,4);
TASK_PP(16'h0ECD,4);
TASK_PP(16'h0ECE,4);
TASK_PP(16'h0ECF,4);
TASK_PP(16'h0ED0,4);
TASK_PP(16'h0ED1,4);
TASK_PP(16'h0ED2,4);
TASK_PP(16'h0ED3,4);
TASK_PP(16'h0ED4,4);
TASK_PP(16'h0ED5,4);
TASK_PP(16'h0ED6,4);
TASK_PP(16'h0ED7,4);
TASK_PP(16'h0ED8,4);
TASK_PP(16'h0ED9,4);
TASK_PP(16'h0EDA,4);
TASK_PP(16'h0EDB,4);
TASK_PP(16'h0EDC,4);
TASK_PP(16'h0EDD,4);
TASK_PP(16'h0EDE,4);
TASK_PP(16'h0EDF,4);
TASK_PP(16'h0EE0,4);
TASK_PP(16'h0EE1,4);
TASK_PP(16'h0EE2,4);
TASK_PP(16'h0EE3,4);
TASK_PP(16'h0EE4,4);
TASK_PP(16'h0EE5,4);
TASK_PP(16'h0EE6,4);
TASK_PP(16'h0EE7,4);
TASK_PP(16'h0EE8,4);
TASK_PP(16'h0EE9,4);
TASK_PP(16'h0EEA,4);
TASK_PP(16'h0EEB,4);
TASK_PP(16'h0EEC,4);
TASK_PP(16'h0EED,4);
TASK_PP(16'h0EEE,4);
TASK_PP(16'h0EEF,4);
TASK_PP(16'h0EF0,4);
TASK_PP(16'h0EF1,4);
TASK_PP(16'h0EF2,4);
TASK_PP(16'h0EF3,4);
TASK_PP(16'h0EF4,4);
TASK_PP(16'h0EF5,4);
TASK_PP(16'h0EF6,4);
TASK_PP(16'h0EF7,4);
TASK_PP(16'h0EF8,4);
TASK_PP(16'h0EF9,4);
TASK_PP(16'h0EFA,4);
TASK_PP(16'h0EFB,4);
TASK_PP(16'h0EFC,4);
TASK_PP(16'h0EFD,4);
TASK_PP(16'h0EFE,4);
TASK_PP(16'h0EFF,4);
TASK_PP(16'h0F00,4);
TASK_PP(16'h0F01,4);
TASK_PP(16'h0F02,4);
TASK_PP(16'h0F03,4);
TASK_PP(16'h0F04,4);
TASK_PP(16'h0F05,4);
TASK_PP(16'h0F06,4);
TASK_PP(16'h0F07,4);
TASK_PP(16'h0F08,4);
TASK_PP(16'h0F09,4);
TASK_PP(16'h0F0A,4);
TASK_PP(16'h0F0B,4);
TASK_PP(16'h0F0C,4);
TASK_PP(16'h0F0D,4);
TASK_PP(16'h0F0E,4);
TASK_PP(16'h0F0F,4);
TASK_PP(16'h0F10,4);
TASK_PP(16'h0F11,4);
TASK_PP(16'h0F12,4);
TASK_PP(16'h0F13,4);
TASK_PP(16'h0F14,4);
TASK_PP(16'h0F15,4);
TASK_PP(16'h0F16,4);
TASK_PP(16'h0F17,4);
TASK_PP(16'h0F18,4);
TASK_PP(16'h0F19,4);
TASK_PP(16'h0F1A,4);
TASK_PP(16'h0F1B,4);
TASK_PP(16'h0F1C,4);
TASK_PP(16'h0F1D,4);
TASK_PP(16'h0F1E,4);
TASK_PP(16'h0F1F,4);
TASK_PP(16'h0F20,4);
TASK_PP(16'h0F21,4);
TASK_PP(16'h0F22,4);
TASK_PP(16'h0F23,4);
TASK_PP(16'h0F24,4);
TASK_PP(16'h0F25,4);
TASK_PP(16'h0F26,4);
TASK_PP(16'h0F27,4);
TASK_PP(16'h0F28,4);
TASK_PP(16'h0F29,4);
TASK_PP(16'h0F2A,4);
TASK_PP(16'h0F2B,4);
TASK_PP(16'h0F2C,4);
TASK_PP(16'h0F2D,4);
TASK_PP(16'h0F2E,4);
TASK_PP(16'h0F2F,4);
TASK_PP(16'h0F30,4);
TASK_PP(16'h0F31,4);
TASK_PP(16'h0F32,4);
TASK_PP(16'h0F33,4);
TASK_PP(16'h0F34,4);
TASK_PP(16'h0F35,4);
TASK_PP(16'h0F36,4);
TASK_PP(16'h0F37,4);
TASK_PP(16'h0F38,4);
TASK_PP(16'h0F39,4);
TASK_PP(16'h0F3A,4);
TASK_PP(16'h0F3B,4);
TASK_PP(16'h0F3C,4);
TASK_PP(16'h0F3D,4);
TASK_PP(16'h0F3E,4);
TASK_PP(16'h0F3F,4);
TASK_PP(16'h0F40,4);
TASK_PP(16'h0F41,4);
TASK_PP(16'h0F42,4);
TASK_PP(16'h0F43,4);
TASK_PP(16'h0F44,4);
TASK_PP(16'h0F45,4);
TASK_PP(16'h0F46,4);
TASK_PP(16'h0F47,4);
TASK_PP(16'h0F48,4);
TASK_PP(16'h0F49,4);
TASK_PP(16'h0F4A,4);
TASK_PP(16'h0F4B,4);
TASK_PP(16'h0F4C,4);
TASK_PP(16'h0F4D,4);
TASK_PP(16'h0F4E,4);
TASK_PP(16'h0F4F,4);
TASK_PP(16'h0F50,4);
TASK_PP(16'h0F51,4);
TASK_PP(16'h0F52,4);
TASK_PP(16'h0F53,4);
TASK_PP(16'h0F54,4);
TASK_PP(16'h0F55,4);
TASK_PP(16'h0F56,4);
TASK_PP(16'h0F57,4);
TASK_PP(16'h0F58,4);
TASK_PP(16'h0F59,4);
TASK_PP(16'h0F5A,4);
TASK_PP(16'h0F5B,4);
TASK_PP(16'h0F5C,4);
TASK_PP(16'h0F5D,4);
TASK_PP(16'h0F5E,4);
TASK_PP(16'h0F5F,4);
TASK_PP(16'h0F60,4);
TASK_PP(16'h0F61,4);
TASK_PP(16'h0F62,4);
TASK_PP(16'h0F63,4);
TASK_PP(16'h0F64,4);
TASK_PP(16'h0F65,4);
TASK_PP(16'h0F66,4);
TASK_PP(16'h0F67,4);
TASK_PP(16'h0F68,4);
TASK_PP(16'h0F69,4);
TASK_PP(16'h0F6A,4);
TASK_PP(16'h0F6B,4);
TASK_PP(16'h0F6C,4);
TASK_PP(16'h0F6D,4);
TASK_PP(16'h0F6E,4);
TASK_PP(16'h0F6F,4);
TASK_PP(16'h0F70,4);
TASK_PP(16'h0F71,4);
TASK_PP(16'h0F72,4);
TASK_PP(16'h0F73,4);
TASK_PP(16'h0F74,4);
TASK_PP(16'h0F75,4);
TASK_PP(16'h0F76,4);
TASK_PP(16'h0F77,4);
TASK_PP(16'h0F78,4);
TASK_PP(16'h0F79,4);
TASK_PP(16'h0F7A,4);
TASK_PP(16'h0F7B,4);
TASK_PP(16'h0F7C,4);
TASK_PP(16'h0F7D,4);
TASK_PP(16'h0F7E,4);
TASK_PP(16'h0F7F,4);
TASK_PP(16'h0F80,4);
TASK_PP(16'h0F81,4);
TASK_PP(16'h0F82,4);
TASK_PP(16'h0F83,4);
TASK_PP(16'h0F84,4);
TASK_PP(16'h0F85,4);
TASK_PP(16'h0F86,4);
TASK_PP(16'h0F87,4);
TASK_PP(16'h0F88,4);
TASK_PP(16'h0F89,4);
TASK_PP(16'h0F8A,4);
TASK_PP(16'h0F8B,4);
TASK_PP(16'h0F8C,4);
TASK_PP(16'h0F8D,4);
TASK_PP(16'h0F8E,4);
TASK_PP(16'h0F8F,4);
TASK_PP(16'h0F90,4);
TASK_PP(16'h0F91,4);
TASK_PP(16'h0F92,4);
TASK_PP(16'h0F93,4);
TASK_PP(16'h0F94,4);
TASK_PP(16'h0F95,4);
TASK_PP(16'h0F96,4);
TASK_PP(16'h0F97,4);
TASK_PP(16'h0F98,4);
TASK_PP(16'h0F99,4);
TASK_PP(16'h0F9A,4);
TASK_PP(16'h0F9B,4);
TASK_PP(16'h0F9C,4);
TASK_PP(16'h0F9D,4);
TASK_PP(16'h0F9E,4);
TASK_PP(16'h0F9F,4);
TASK_PP(16'h0FA0,4);
TASK_PP(16'h0FA1,4);
TASK_PP(16'h0FA2,4);
TASK_PP(16'h0FA3,4);
TASK_PP(16'h0FA4,4);
TASK_PP(16'h0FA5,4);
TASK_PP(16'h0FA6,4);
TASK_PP(16'h0FA7,4);
TASK_PP(16'h0FA8,4);
TASK_PP(16'h0FA9,4);
TASK_PP(16'h0FAA,4);
TASK_PP(16'h0FAB,4);
TASK_PP(16'h0FAC,4);
TASK_PP(16'h0FAD,4);
TASK_PP(16'h0FAE,4);
TASK_PP(16'h0FAF,4);
TASK_PP(16'h0FB0,4);
TASK_PP(16'h0FB1,4);
TASK_PP(16'h0FB2,4);
TASK_PP(16'h0FB3,4);
TASK_PP(16'h0FB4,4);
TASK_PP(16'h0FB5,4);
TASK_PP(16'h0FB6,4);
TASK_PP(16'h0FB7,4);
TASK_PP(16'h0FB8,4);
TASK_PP(16'h0FB9,4);
TASK_PP(16'h0FBA,4);
TASK_PP(16'h0FBB,4);
TASK_PP(16'h0FBC,4);
TASK_PP(16'h0FBD,4);
TASK_PP(16'h0FBE,4);
TASK_PP(16'h0FBF,4);
TASK_PP(16'h0FC0,4);
TASK_PP(16'h0FC1,4);
TASK_PP(16'h0FC2,4);
TASK_PP(16'h0FC3,4);
TASK_PP(16'h0FC4,4);
TASK_PP(16'h0FC5,4);
TASK_PP(16'h0FC6,4);
TASK_PP(16'h0FC7,4);
TASK_PP(16'h0FC8,4);
TASK_PP(16'h0FC9,4);
TASK_PP(16'h0FCA,4);
TASK_PP(16'h0FCB,4);
TASK_PP(16'h0FCC,4);
TASK_PP(16'h0FCD,4);
TASK_PP(16'h0FCE,4);
TASK_PP(16'h0FCF,4);
TASK_PP(16'h0FD0,4);
TASK_PP(16'h0FD1,4);
TASK_PP(16'h0FD2,4);
TASK_PP(16'h0FD3,4);
TASK_PP(16'h0FD4,4);
TASK_PP(16'h0FD5,4);
TASK_PP(16'h0FD6,4);
TASK_PP(16'h0FD7,4);
TASK_PP(16'h0FD8,4);
TASK_PP(16'h0FD9,4);
TASK_PP(16'h0FDA,4);
TASK_PP(16'h0FDB,4);
TASK_PP(16'h0FDC,4);
TASK_PP(16'h0FDD,4);
TASK_PP(16'h0FDE,4);
TASK_PP(16'h0FDF,4);
TASK_PP(16'h0FE0,4);
TASK_PP(16'h0FE1,4);
TASK_PP(16'h0FE2,4);
TASK_PP(16'h0FE3,4);
TASK_PP(16'h0FE4,4);
TASK_PP(16'h0FE5,4);
TASK_PP(16'h0FE6,4);
TASK_PP(16'h0FE7,4);
TASK_PP(16'h0FE8,4);
TASK_PP(16'h0FE9,4);
TASK_PP(16'h0FEA,4);
TASK_PP(16'h0FEB,4);
TASK_PP(16'h0FEC,4);
TASK_PP(16'h0FED,4);
TASK_PP(16'h0FEE,4);
TASK_PP(16'h0FEF,4);
TASK_PP(16'h0FF0,4);
TASK_PP(16'h0FF1,4);
TASK_PP(16'h0FF2,4);
TASK_PP(16'h0FF3,4);
TASK_PP(16'h0FF4,4);
TASK_PP(16'h0FF5,4);
TASK_PP(16'h0FF6,4);
TASK_PP(16'h0FF7,4);
TASK_PP(16'h0FF8,4);
TASK_PP(16'h0FF9,4);
TASK_PP(16'h0FFA,4);
TASK_PP(16'h0FFB,4);
TASK_PP(16'h0FFC,4);
TASK_PP(16'h0FFD,4);
TASK_PP(16'h0FFE,4);
TASK_PP(16'h0FFF,4);
TASK_PP(16'h1000,4);
TASK_PP(16'h1001,4);
TASK_PP(16'h1002,4);
TASK_PP(16'h1003,4);
TASK_PP(16'h1004,4);
TASK_PP(16'h1005,4);
TASK_PP(16'h1006,4);
TASK_PP(16'h1007,4);
TASK_PP(16'h1008,4);
TASK_PP(16'h1009,4);
TASK_PP(16'h100A,4);
TASK_PP(16'h100B,4);
TASK_PP(16'h100C,4);
TASK_PP(16'h100D,4);
TASK_PP(16'h100E,4);
TASK_PP(16'h100F,4);
TASK_PP(16'h1010,4);
TASK_PP(16'h1011,4);
TASK_PP(16'h1012,4);
TASK_PP(16'h1013,4);
TASK_PP(16'h1014,4);
TASK_PP(16'h1015,4);
TASK_PP(16'h1016,4);
TASK_PP(16'h1017,4);
TASK_PP(16'h1018,4);
TASK_PP(16'h1019,4);
TASK_PP(16'h101A,4);
TASK_PP(16'h101B,4);
TASK_PP(16'h101C,4);
TASK_PP(16'h101D,4);
TASK_PP(16'h101E,4);
TASK_PP(16'h101F,4);
TASK_PP(16'h1020,4);
TASK_PP(16'h1021,4);
TASK_PP(16'h1022,4);
TASK_PP(16'h1023,4);
TASK_PP(16'h1024,4);
TASK_PP(16'h1025,4);
TASK_PP(16'h1026,4);
TASK_PP(16'h1027,4);
TASK_PP(16'h1028,4);
TASK_PP(16'h1029,4);
TASK_PP(16'h102A,4);
TASK_PP(16'h102B,4);
TASK_PP(16'h102C,4);
TASK_PP(16'h102D,4);
TASK_PP(16'h102E,4);
TASK_PP(16'h102F,4);
TASK_PP(16'h1030,4);
TASK_PP(16'h1031,4);
TASK_PP(16'h1032,4);
TASK_PP(16'h1033,4);
TASK_PP(16'h1034,4);
TASK_PP(16'h1035,4);
TASK_PP(16'h1036,4);
TASK_PP(16'h1037,4);
TASK_PP(16'h1038,4);
TASK_PP(16'h1039,4);
TASK_PP(16'h103A,4);
TASK_PP(16'h103B,4);
TASK_PP(16'h103C,4);
TASK_PP(16'h103D,4);
TASK_PP(16'h103E,4);
TASK_PP(16'h103F,4);
TASK_PP(16'h1040,4);
TASK_PP(16'h1041,4);
TASK_PP(16'h1042,4);
TASK_PP(16'h1043,4);
TASK_PP(16'h1044,4);
TASK_PP(16'h1045,4);
TASK_PP(16'h1046,4);
TASK_PP(16'h1047,4);
TASK_PP(16'h1048,4);
TASK_PP(16'h1049,4);
TASK_PP(16'h104A,4);
TASK_PP(16'h104B,4);
TASK_PP(16'h104C,4);
TASK_PP(16'h104D,4);
TASK_PP(16'h104E,4);
TASK_PP(16'h104F,4);
TASK_PP(16'h1050,4);
TASK_PP(16'h1051,4);
TASK_PP(16'h1052,4);
TASK_PP(16'h1053,4);
TASK_PP(16'h1054,4);
TASK_PP(16'h1055,4);
TASK_PP(16'h1056,4);
TASK_PP(16'h1057,4);
TASK_PP(16'h1058,4);
TASK_PP(16'h1059,4);
TASK_PP(16'h105A,4);
TASK_PP(16'h105B,4);
TASK_PP(16'h105C,4);
TASK_PP(16'h105D,4);
TASK_PP(16'h105E,4);
TASK_PP(16'h105F,4);
TASK_PP(16'h1060,4);
TASK_PP(16'h1061,4);
TASK_PP(16'h1062,4);
TASK_PP(16'h1063,4);
TASK_PP(16'h1064,4);
TASK_PP(16'h1065,4);
TASK_PP(16'h1066,4);
TASK_PP(16'h1067,4);
TASK_PP(16'h1068,4);
TASK_PP(16'h1069,4);
TASK_PP(16'h106A,4);
TASK_PP(16'h106B,4);
TASK_PP(16'h106C,4);
TASK_PP(16'h106D,4);
TASK_PP(16'h106E,4);
TASK_PP(16'h106F,4);
TASK_PP(16'h1070,4);
TASK_PP(16'h1071,4);
TASK_PP(16'h1072,4);
TASK_PP(16'h1073,4);
TASK_PP(16'h1074,4);
TASK_PP(16'h1075,4);
TASK_PP(16'h1076,4);
TASK_PP(16'h1077,4);
TASK_PP(16'h1078,4);
TASK_PP(16'h1079,4);
TASK_PP(16'h107A,4);
TASK_PP(16'h107B,4);
TASK_PP(16'h107C,4);
TASK_PP(16'h107D,4);
TASK_PP(16'h107E,4);
TASK_PP(16'h107F,4);
TASK_PP(16'h1080,4);
TASK_PP(16'h1081,4);
TASK_PP(16'h1082,4);
TASK_PP(16'h1083,4);
TASK_PP(16'h1084,4);
TASK_PP(16'h1085,4);
TASK_PP(16'h1086,4);
TASK_PP(16'h1087,4);
TASK_PP(16'h1088,4);
TASK_PP(16'h1089,4);
TASK_PP(16'h108A,4);
TASK_PP(16'h108B,4);
TASK_PP(16'h108C,4);
TASK_PP(16'h108D,4);
TASK_PP(16'h108E,4);
TASK_PP(16'h108F,4);
TASK_PP(16'h1090,4);
TASK_PP(16'h1091,4);
TASK_PP(16'h1092,4);
TASK_PP(16'h1093,4);
TASK_PP(16'h1094,4);
TASK_PP(16'h1095,4);
TASK_PP(16'h1096,4);
TASK_PP(16'h1097,4);
TASK_PP(16'h1098,4);
TASK_PP(16'h1099,4);
TASK_PP(16'h109A,4);
TASK_PP(16'h109B,4);
TASK_PP(16'h109C,4);
TASK_PP(16'h109D,4);
TASK_PP(16'h109E,4);
TASK_PP(16'h109F,4);
TASK_PP(16'h10A0,4);
TASK_PP(16'h10A1,4);
TASK_PP(16'h10A2,4);
TASK_PP(16'h10A3,4);
TASK_PP(16'h10A4,4);
TASK_PP(16'h10A5,4);
TASK_PP(16'h10A6,4);
TASK_PP(16'h10A7,4);
TASK_PP(16'h10A8,4);
TASK_PP(16'h10A9,4);
TASK_PP(16'h10AA,4);
TASK_PP(16'h10AB,4);
TASK_PP(16'h10AC,4);
TASK_PP(16'h10AD,4);
TASK_PP(16'h10AE,4);
TASK_PP(16'h10AF,4);
TASK_PP(16'h10B0,4);
TASK_PP(16'h10B1,4);
TASK_PP(16'h10B2,4);
TASK_PP(16'h10B3,4);
TASK_PP(16'h10B4,4);
TASK_PP(16'h10B5,4);
TASK_PP(16'h10B6,4);
TASK_PP(16'h10B7,4);
TASK_PP(16'h10B8,4);
TASK_PP(16'h10B9,4);
TASK_PP(16'h10BA,4);
TASK_PP(16'h10BB,4);
TASK_PP(16'h10BC,4);
TASK_PP(16'h10BD,4);
TASK_PP(16'h10BE,4);
TASK_PP(16'h10BF,4);
TASK_PP(16'h10C0,4);
TASK_PP(16'h10C1,4);
TASK_PP(16'h10C2,4);
TASK_PP(16'h10C3,4);
TASK_PP(16'h10C4,4);
TASK_PP(16'h10C5,4);
TASK_PP(16'h10C6,4);
TASK_PP(16'h10C7,4);
TASK_PP(16'h10C8,4);
TASK_PP(16'h10C9,4);
TASK_PP(16'h10CA,4);
TASK_PP(16'h10CB,4);
TASK_PP(16'h10CC,4);
TASK_PP(16'h10CD,4);
TASK_PP(16'h10CE,4);
TASK_PP(16'h10CF,4);
TASK_PP(16'h10D0,4);
TASK_PP(16'h10D1,4);
TASK_PP(16'h10D2,4);
TASK_PP(16'h10D3,4);
TASK_PP(16'h10D4,4);
TASK_PP(16'h10D5,4);
TASK_PP(16'h10D6,4);
TASK_PP(16'h10D7,4);
TASK_PP(16'h10D8,4);
TASK_PP(16'h10D9,4);
TASK_PP(16'h10DA,4);
TASK_PP(16'h10DB,4);
TASK_PP(16'h10DC,4);
TASK_PP(16'h10DD,4);
TASK_PP(16'h10DE,4);
TASK_PP(16'h10DF,4);
TASK_PP(16'h10E0,4);
TASK_PP(16'h10E1,4);
TASK_PP(16'h10E2,4);
TASK_PP(16'h10E3,4);
TASK_PP(16'h10E4,4);
TASK_PP(16'h10E5,4);
TASK_PP(16'h10E6,4);
TASK_PP(16'h10E7,4);
TASK_PP(16'h10E8,4);
TASK_PP(16'h10E9,4);
TASK_PP(16'h10EA,4);
TASK_PP(16'h10EB,4);
TASK_PP(16'h10EC,4);
TASK_PP(16'h10ED,4);
TASK_PP(16'h10EE,4);
TASK_PP(16'h10EF,4);
TASK_PP(16'h10F0,4);
TASK_PP(16'h10F1,4);
TASK_PP(16'h10F2,4);
TASK_PP(16'h10F3,4);
TASK_PP(16'h10F4,4);
TASK_PP(16'h10F5,4);
TASK_PP(16'h10F6,4);
TASK_PP(16'h10F7,4);
TASK_PP(16'h10F8,4);
TASK_PP(16'h10F9,4);
TASK_PP(16'h10FA,4);
TASK_PP(16'h10FB,4);
TASK_PP(16'h10FC,4);
TASK_PP(16'h10FD,4);
TASK_PP(16'h10FE,4);
TASK_PP(16'h10FF,4);
TASK_PP(16'h1100,4);
TASK_PP(16'h1101,4);
TASK_PP(16'h1102,4);
TASK_PP(16'h1103,4);
TASK_PP(16'h1104,4);
TASK_PP(16'h1105,4);
TASK_PP(16'h1106,4);
TASK_PP(16'h1107,4);
TASK_PP(16'h1108,4);
TASK_PP(16'h1109,4);
TASK_PP(16'h110A,4);
TASK_PP(16'h110B,4);
TASK_PP(16'h110C,4);
TASK_PP(16'h110D,4);
TASK_PP(16'h110E,4);
TASK_PP(16'h110F,4);
TASK_PP(16'h1110,4);
TASK_PP(16'h1111,4);
TASK_PP(16'h1112,4);
TASK_PP(16'h1113,4);
TASK_PP(16'h1114,4);
TASK_PP(16'h1115,4);
TASK_PP(16'h1116,4);
TASK_PP(16'h1117,4);
TASK_PP(16'h1118,4);
TASK_PP(16'h1119,4);
TASK_PP(16'h111A,4);
TASK_PP(16'h111B,4);
TASK_PP(16'h111C,4);
TASK_PP(16'h111D,4);
TASK_PP(16'h111E,4);
TASK_PP(16'h111F,4);
TASK_PP(16'h1120,4);
TASK_PP(16'h1121,4);
TASK_PP(16'h1122,4);
TASK_PP(16'h1123,4);
TASK_PP(16'h1124,4);
TASK_PP(16'h1125,4);
TASK_PP(16'h1126,4);
TASK_PP(16'h1127,4);
TASK_PP(16'h1128,4);
TASK_PP(16'h1129,4);
TASK_PP(16'h112A,4);
TASK_PP(16'h112B,4);
TASK_PP(16'h112C,4);
TASK_PP(16'h112D,4);
TASK_PP(16'h112E,4);
TASK_PP(16'h112F,4);
TASK_PP(16'h1130,4);
TASK_PP(16'h1131,4);
TASK_PP(16'h1132,4);
TASK_PP(16'h1133,4);
TASK_PP(16'h1134,4);
TASK_PP(16'h1135,4);
TASK_PP(16'h1136,4);
TASK_PP(16'h1137,4);
TASK_PP(16'h1138,4);
TASK_PP(16'h1139,4);
TASK_PP(16'h113A,4);
TASK_PP(16'h113B,4);
TASK_PP(16'h113C,4);
TASK_PP(16'h113D,4);
TASK_PP(16'h113E,4);
TASK_PP(16'h113F,4);
TASK_PP(16'h1140,4);
TASK_PP(16'h1141,4);
TASK_PP(16'h1142,4);
TASK_PP(16'h1143,4);
TASK_PP(16'h1144,4);
TASK_PP(16'h1145,4);
TASK_PP(16'h1146,4);
TASK_PP(16'h1147,4);
TASK_PP(16'h1148,4);
TASK_PP(16'h1149,4);
TASK_PP(16'h114A,4);
TASK_PP(16'h114B,4);
TASK_PP(16'h114C,4);
TASK_PP(16'h114D,4);
TASK_PP(16'h114E,4);
TASK_PP(16'h114F,4);
TASK_PP(16'h1150,4);
TASK_PP(16'h1151,4);
TASK_PP(16'h1152,4);
TASK_PP(16'h1153,4);
TASK_PP(16'h1154,4);
TASK_PP(16'h1155,4);
TASK_PP(16'h1156,4);
TASK_PP(16'h1157,4);
TASK_PP(16'h1158,4);
TASK_PP(16'h1159,4);
TASK_PP(16'h115A,4);
TASK_PP(16'h115B,4);
TASK_PP(16'h115C,4);
TASK_PP(16'h115D,4);
TASK_PP(16'h115E,4);
TASK_PP(16'h115F,4);
TASK_PP(16'h1160,4);
TASK_PP(16'h1161,4);
TASK_PP(16'h1162,4);
TASK_PP(16'h1163,4);
TASK_PP(16'h1164,4);
TASK_PP(16'h1165,4);
TASK_PP(16'h1166,4);
TASK_PP(16'h1167,4);
TASK_PP(16'h1168,4);
TASK_PP(16'h1169,4);
TASK_PP(16'h116A,4);
TASK_PP(16'h116B,4);
TASK_PP(16'h116C,4);
TASK_PP(16'h116D,4);
TASK_PP(16'h116E,4);
TASK_PP(16'h116F,4);
TASK_PP(16'h1170,4);
TASK_PP(16'h1171,4);
TASK_PP(16'h1172,4);
TASK_PP(16'h1173,4);
TASK_PP(16'h1174,4);
TASK_PP(16'h1175,4);
TASK_PP(16'h1176,4);
TASK_PP(16'h1177,4);
TASK_PP(16'h1178,4);
TASK_PP(16'h1179,4);
TASK_PP(16'h117A,4);
TASK_PP(16'h117B,4);
TASK_PP(16'h117C,4);
TASK_PP(16'h117D,4);
TASK_PP(16'h117E,4);
TASK_PP(16'h117F,4);
TASK_PP(16'h1180,4);
TASK_PP(16'h1181,4);
TASK_PP(16'h1182,4);
TASK_PP(16'h1183,4);
TASK_PP(16'h1184,4);
TASK_PP(16'h1185,4);
TASK_PP(16'h1186,4);
TASK_PP(16'h1187,4);
TASK_PP(16'h1188,4);
TASK_PP(16'h1189,4);
TASK_PP(16'h118A,4);
TASK_PP(16'h118B,4);
TASK_PP(16'h118C,4);
TASK_PP(16'h118D,4);
TASK_PP(16'h118E,4);
TASK_PP(16'h118F,4);
TASK_PP(16'h1190,4);
TASK_PP(16'h1191,4);
TASK_PP(16'h1192,4);
TASK_PP(16'h1193,4);
TASK_PP(16'h1194,4);
TASK_PP(16'h1195,4);
TASK_PP(16'h1196,4);
TASK_PP(16'h1197,4);
TASK_PP(16'h1198,4);
TASK_PP(16'h1199,4);
TASK_PP(16'h119A,4);
TASK_PP(16'h119B,4);
TASK_PP(16'h119C,4);
TASK_PP(16'h119D,4);
TASK_PP(16'h119E,4);
TASK_PP(16'h119F,4);
TASK_PP(16'h11A0,4);
TASK_PP(16'h11A1,4);
TASK_PP(16'h11A2,4);
TASK_PP(16'h11A3,4);
TASK_PP(16'h11A4,4);
TASK_PP(16'h11A5,4);
TASK_PP(16'h11A6,4);
TASK_PP(16'h11A7,4);
TASK_PP(16'h11A8,4);
TASK_PP(16'h11A9,4);
TASK_PP(16'h11AA,4);
TASK_PP(16'h11AB,4);
TASK_PP(16'h11AC,4);
TASK_PP(16'h11AD,4);
TASK_PP(16'h11AE,4);
TASK_PP(16'h11AF,4);
TASK_PP(16'h11B0,4);
TASK_PP(16'h11B1,4);
TASK_PP(16'h11B2,4);
TASK_PP(16'h11B3,4);
TASK_PP(16'h11B4,4);
TASK_PP(16'h11B5,4);
TASK_PP(16'h11B6,4);
TASK_PP(16'h11B7,4);
TASK_PP(16'h11B8,4);
TASK_PP(16'h11B9,4);
TASK_PP(16'h11BA,4);
TASK_PP(16'h11BB,4);
TASK_PP(16'h11BC,4);
TASK_PP(16'h11BD,4);
TASK_PP(16'h11BE,4);
TASK_PP(16'h11BF,4);
TASK_PP(16'h11C0,4);
TASK_PP(16'h11C1,4);
TASK_PP(16'h11C2,4);
TASK_PP(16'h11C3,4);
TASK_PP(16'h11C4,4);
TASK_PP(16'h11C5,4);
TASK_PP(16'h11C6,4);
TASK_PP(16'h11C7,4);
TASK_PP(16'h11C8,4);
TASK_PP(16'h11C9,4);
TASK_PP(16'h11CA,4);
TASK_PP(16'h11CB,4);
TASK_PP(16'h11CC,4);
TASK_PP(16'h11CD,4);
TASK_PP(16'h11CE,4);
TASK_PP(16'h11CF,4);
TASK_PP(16'h11D0,4);
TASK_PP(16'h11D1,4);
TASK_PP(16'h11D2,4);
TASK_PP(16'h11D3,4);
TASK_PP(16'h11D4,4);
TASK_PP(16'h11D5,4);
TASK_PP(16'h11D6,4);
TASK_PP(16'h11D7,4);
TASK_PP(16'h11D8,4);
TASK_PP(16'h11D9,4);
TASK_PP(16'h11DA,4);
TASK_PP(16'h11DB,4);
TASK_PP(16'h11DC,4);
TASK_PP(16'h11DD,4);
TASK_PP(16'h11DE,4);
TASK_PP(16'h11DF,4);
TASK_PP(16'h11E0,4);
TASK_PP(16'h11E1,4);
TASK_PP(16'h11E2,4);
TASK_PP(16'h11E3,4);
TASK_PP(16'h11E4,4);
TASK_PP(16'h11E5,4);
TASK_PP(16'h11E6,4);
TASK_PP(16'h11E7,4);
TASK_PP(16'h11E8,4);
TASK_PP(16'h11E9,4);
TASK_PP(16'h11EA,4);
TASK_PP(16'h11EB,4);
TASK_PP(16'h11EC,4);
TASK_PP(16'h11ED,4);
TASK_PP(16'h11EE,4);
TASK_PP(16'h11EF,4);
TASK_PP(16'h11F0,4);
TASK_PP(16'h11F1,4);
TASK_PP(16'h11F2,4);
TASK_PP(16'h11F3,4);
TASK_PP(16'h11F4,4);
TASK_PP(16'h11F5,4);
TASK_PP(16'h11F6,4);
TASK_PP(16'h11F7,4);
TASK_PP(16'h11F8,4);
TASK_PP(16'h11F9,4);
TASK_PP(16'h11FA,4);
TASK_PP(16'h11FB,4);
TASK_PP(16'h11FC,4);
TASK_PP(16'h11FD,4);
TASK_PP(16'h11FE,4);
TASK_PP(16'h11FF,4);
TASK_PP(16'h1200,4);
TASK_PP(16'h1201,4);
TASK_PP(16'h1202,4);
TASK_PP(16'h1203,4);
TASK_PP(16'h1204,4);
TASK_PP(16'h1205,4);
TASK_PP(16'h1206,4);
TASK_PP(16'h1207,4);
TASK_PP(16'h1208,4);
TASK_PP(16'h1209,4);
TASK_PP(16'h120A,4);
TASK_PP(16'h120B,4);
TASK_PP(16'h120C,4);
TASK_PP(16'h120D,4);
TASK_PP(16'h120E,4);
TASK_PP(16'h120F,4);
TASK_PP(16'h1210,4);
TASK_PP(16'h1211,4);
TASK_PP(16'h1212,4);
TASK_PP(16'h1213,4);
TASK_PP(16'h1214,4);
TASK_PP(16'h1215,4);
TASK_PP(16'h1216,4);
TASK_PP(16'h1217,4);
TASK_PP(16'h1218,4);
TASK_PP(16'h1219,4);
TASK_PP(16'h121A,4);
TASK_PP(16'h121B,4);
TASK_PP(16'h121C,4);
TASK_PP(16'h121D,4);
TASK_PP(16'h121E,4);
TASK_PP(16'h121F,4);
TASK_PP(16'h1220,4);
TASK_PP(16'h1221,4);
TASK_PP(16'h1222,4);
TASK_PP(16'h1223,4);
TASK_PP(16'h1224,4);
TASK_PP(16'h1225,4);
TASK_PP(16'h1226,4);
TASK_PP(16'h1227,4);
TASK_PP(16'h1228,4);
TASK_PP(16'h1229,4);
TASK_PP(16'h122A,4);
TASK_PP(16'h122B,4);
TASK_PP(16'h122C,4);
TASK_PP(16'h122D,4);
TASK_PP(16'h122E,4);
TASK_PP(16'h122F,4);
TASK_PP(16'h1230,4);
TASK_PP(16'h1231,4);
TASK_PP(16'h1232,4);
TASK_PP(16'h1233,4);
TASK_PP(16'h1234,4);
TASK_PP(16'h1235,4);
TASK_PP(16'h1236,4);
TASK_PP(16'h1237,4);
TASK_PP(16'h1238,4);
TASK_PP(16'h1239,4);
TASK_PP(16'h123A,4);
TASK_PP(16'h123B,4);
TASK_PP(16'h123C,4);
TASK_PP(16'h123D,4);
TASK_PP(16'h123E,4);
TASK_PP(16'h123F,4);
TASK_PP(16'h1240,4);
TASK_PP(16'h1241,4);
TASK_PP(16'h1242,4);
TASK_PP(16'h1243,4);
TASK_PP(16'h1244,4);
TASK_PP(16'h1245,4);
TASK_PP(16'h1246,4);
TASK_PP(16'h1247,4);
TASK_PP(16'h1248,4);
TASK_PP(16'h1249,4);
TASK_PP(16'h124A,4);
TASK_PP(16'h124B,4);
TASK_PP(16'h124C,4);
TASK_PP(16'h124D,4);
TASK_PP(16'h124E,4);
TASK_PP(16'h124F,4);
TASK_PP(16'h1250,4);
TASK_PP(16'h1251,4);
TASK_PP(16'h1252,4);
TASK_PP(16'h1253,4);
TASK_PP(16'h1254,4);
TASK_PP(16'h1255,4);
TASK_PP(16'h1256,4);
TASK_PP(16'h1257,4);
TASK_PP(16'h1258,4);
TASK_PP(16'h1259,4);
TASK_PP(16'h125A,4);
TASK_PP(16'h125B,4);
TASK_PP(16'h125C,4);
TASK_PP(16'h125D,4);
TASK_PP(16'h125E,4);
TASK_PP(16'h125F,4);
TASK_PP(16'h1260,4);
TASK_PP(16'h1261,4);
TASK_PP(16'h1262,4);
TASK_PP(16'h1263,4);
TASK_PP(16'h1264,4);
TASK_PP(16'h1265,4);
TASK_PP(16'h1266,4);
TASK_PP(16'h1267,4);
TASK_PP(16'h1268,4);
TASK_PP(16'h1269,4);
TASK_PP(16'h126A,4);
TASK_PP(16'h126B,4);
TASK_PP(16'h126C,4);
TASK_PP(16'h126D,4);
TASK_PP(16'h126E,4);
TASK_PP(16'h126F,4);
TASK_PP(16'h1270,4);
TASK_PP(16'h1271,4);
TASK_PP(16'h1272,4);
TASK_PP(16'h1273,4);
TASK_PP(16'h1274,4);
TASK_PP(16'h1275,4);
TASK_PP(16'h1276,4);
TASK_PP(16'h1277,4);
TASK_PP(16'h1278,4);
TASK_PP(16'h1279,4);
TASK_PP(16'h127A,4);
TASK_PP(16'h127B,4);
TASK_PP(16'h127C,4);
TASK_PP(16'h127D,4);
TASK_PP(16'h127E,4);
TASK_PP(16'h127F,4);
TASK_PP(16'h1280,4);
TASK_PP(16'h1281,4);
TASK_PP(16'h1282,4);
TASK_PP(16'h1283,4);
TASK_PP(16'h1284,4);
TASK_PP(16'h1285,4);
TASK_PP(16'h1286,4);
TASK_PP(16'h1287,4);
TASK_PP(16'h1288,4);
TASK_PP(16'h1289,4);
TASK_PP(16'h128A,4);
TASK_PP(16'h128B,4);
TASK_PP(16'h128C,4);
TASK_PP(16'h128D,4);
TASK_PP(16'h128E,4);
TASK_PP(16'h128F,4);
TASK_PP(16'h1290,4);
TASK_PP(16'h1291,4);
TASK_PP(16'h1292,4);
TASK_PP(16'h1293,4);
TASK_PP(16'h1294,4);
TASK_PP(16'h1295,4);
TASK_PP(16'h1296,4);
TASK_PP(16'h1297,4);
TASK_PP(16'h1298,4);
TASK_PP(16'h1299,4);
TASK_PP(16'h129A,4);
TASK_PP(16'h129B,4);
TASK_PP(16'h129C,4);
TASK_PP(16'h129D,4);
TASK_PP(16'h129E,4);
TASK_PP(16'h129F,4);
TASK_PP(16'h12A0,4);
TASK_PP(16'h12A1,4);
TASK_PP(16'h12A2,4);
TASK_PP(16'h12A3,4);
TASK_PP(16'h12A4,4);
TASK_PP(16'h12A5,4);
TASK_PP(16'h12A6,4);
TASK_PP(16'h12A7,4);
TASK_PP(16'h12A8,4);
TASK_PP(16'h12A9,4);
TASK_PP(16'h12AA,4);
TASK_PP(16'h12AB,4);
TASK_PP(16'h12AC,4);
TASK_PP(16'h12AD,4);
TASK_PP(16'h12AE,4);
TASK_PP(16'h12AF,4);
TASK_PP(16'h12B0,4);
TASK_PP(16'h12B1,4);
TASK_PP(16'h12B2,4);
TASK_PP(16'h12B3,4);
TASK_PP(16'h12B4,4);
TASK_PP(16'h12B5,4);
TASK_PP(16'h12B6,4);
TASK_PP(16'h12B7,4);
TASK_PP(16'h12B8,4);
TASK_PP(16'h12B9,4);
TASK_PP(16'h12BA,4);
TASK_PP(16'h12BB,4);
TASK_PP(16'h12BC,4);
TASK_PP(16'h12BD,4);
TASK_PP(16'h12BE,4);
TASK_PP(16'h12BF,4);
TASK_PP(16'h12C0,4);
TASK_PP(16'h12C1,4);
TASK_PP(16'h12C2,4);
TASK_PP(16'h12C3,4);
TASK_PP(16'h12C4,4);
TASK_PP(16'h12C5,4);
TASK_PP(16'h12C6,4);
TASK_PP(16'h12C7,4);
TASK_PP(16'h12C8,4);
TASK_PP(16'h12C9,4);
TASK_PP(16'h12CA,4);
TASK_PP(16'h12CB,4);
TASK_PP(16'h12CC,4);
TASK_PP(16'h12CD,4);
TASK_PP(16'h12CE,4);
TASK_PP(16'h12CF,4);
TASK_PP(16'h12D0,4);
TASK_PP(16'h12D1,4);
TASK_PP(16'h12D2,4);
TASK_PP(16'h12D3,4);
TASK_PP(16'h12D4,4);
TASK_PP(16'h12D5,4);
TASK_PP(16'h12D6,4);
TASK_PP(16'h12D7,4);
TASK_PP(16'h12D8,4);
TASK_PP(16'h12D9,4);
TASK_PP(16'h12DA,4);
TASK_PP(16'h12DB,4);
TASK_PP(16'h12DC,4);
TASK_PP(16'h12DD,4);
TASK_PP(16'h12DE,4);
TASK_PP(16'h12DF,4);
TASK_PP(16'h12E0,4);
TASK_PP(16'h12E1,4);
TASK_PP(16'h12E2,4);
TASK_PP(16'h12E3,4);
TASK_PP(16'h12E4,4);
TASK_PP(16'h12E5,4);
TASK_PP(16'h12E6,4);
TASK_PP(16'h12E7,4);
TASK_PP(16'h12E8,4);
TASK_PP(16'h12E9,4);
TASK_PP(16'h12EA,4);
TASK_PP(16'h12EB,4);
TASK_PP(16'h12EC,4);
TASK_PP(16'h12ED,4);
TASK_PP(16'h12EE,4);
TASK_PP(16'h12EF,4);
TASK_PP(16'h12F0,4);
TASK_PP(16'h12F1,4);
TASK_PP(16'h12F2,4);
TASK_PP(16'h12F3,4);
TASK_PP(16'h12F4,4);
TASK_PP(16'h12F5,4);
TASK_PP(16'h12F6,4);
TASK_PP(16'h12F7,4);
TASK_PP(16'h12F8,4);
TASK_PP(16'h12F9,4);
TASK_PP(16'h12FA,4);
TASK_PP(16'h12FB,4);
TASK_PP(16'h12FC,4);
TASK_PP(16'h12FD,4);
TASK_PP(16'h12FE,4);
TASK_PP(16'h12FF,4);
TASK_PP(16'h1300,4);
TASK_PP(16'h1301,4);
TASK_PP(16'h1302,4);
TASK_PP(16'h1303,4);
TASK_PP(16'h1304,4);
TASK_PP(16'h1305,4);
TASK_PP(16'h1306,4);
TASK_PP(16'h1307,4);
TASK_PP(16'h1308,4);
TASK_PP(16'h1309,4);
TASK_PP(16'h130A,4);
TASK_PP(16'h130B,4);
TASK_PP(16'h130C,4);
TASK_PP(16'h130D,4);
TASK_PP(16'h130E,4);
TASK_PP(16'h130F,4);
TASK_PP(16'h1310,4);
TASK_PP(16'h1311,4);
TASK_PP(16'h1312,4);
TASK_PP(16'h1313,4);
TASK_PP(16'h1314,4);
TASK_PP(16'h1315,4);
TASK_PP(16'h1316,4);
TASK_PP(16'h1317,4);
TASK_PP(16'h1318,4);
TASK_PP(16'h1319,4);
TASK_PP(16'h131A,4);
TASK_PP(16'h131B,4);
TASK_PP(16'h131C,4);
TASK_PP(16'h131D,4);
TASK_PP(16'h131E,4);
TASK_PP(16'h131F,4);
TASK_PP(16'h1320,4);
TASK_PP(16'h1321,4);
TASK_PP(16'h1322,4);
TASK_PP(16'h1323,4);
TASK_PP(16'h1324,4);
TASK_PP(16'h1325,4);
TASK_PP(16'h1326,4);
TASK_PP(16'h1327,4);
TASK_PP(16'h1328,4);
TASK_PP(16'h1329,4);
TASK_PP(16'h132A,4);
TASK_PP(16'h132B,4);
TASK_PP(16'h132C,4);
TASK_PP(16'h132D,4);
TASK_PP(16'h132E,4);
TASK_PP(16'h132F,4);
TASK_PP(16'h1330,4);
TASK_PP(16'h1331,4);
TASK_PP(16'h1332,4);
TASK_PP(16'h1333,4);
TASK_PP(16'h1334,4);
TASK_PP(16'h1335,4);
TASK_PP(16'h1336,4);
TASK_PP(16'h1337,4);
TASK_PP(16'h1338,4);
TASK_PP(16'h1339,4);
TASK_PP(16'h133A,4);
TASK_PP(16'h133B,4);
TASK_PP(16'h133C,4);
TASK_PP(16'h133D,4);
TASK_PP(16'h133E,4);
TASK_PP(16'h133F,4);
TASK_PP(16'h1340,4);
TASK_PP(16'h1341,4);
TASK_PP(16'h1342,4);
TASK_PP(16'h1343,4);
TASK_PP(16'h1344,4);
TASK_PP(16'h1345,4);
TASK_PP(16'h1346,4);
TASK_PP(16'h1347,4);
TASK_PP(16'h1348,4);
TASK_PP(16'h1349,4);
TASK_PP(16'h134A,4);
TASK_PP(16'h134B,4);
TASK_PP(16'h134C,4);
TASK_PP(16'h134D,4);
TASK_PP(16'h134E,4);
TASK_PP(16'h134F,4);
TASK_PP(16'h1350,4);
TASK_PP(16'h1351,4);
TASK_PP(16'h1352,4);
TASK_PP(16'h1353,4);
TASK_PP(16'h1354,4);
TASK_PP(16'h1355,4);
TASK_PP(16'h1356,4);
TASK_PP(16'h1357,4);
TASK_PP(16'h1358,4);
TASK_PP(16'h1359,4);
TASK_PP(16'h135A,4);
TASK_PP(16'h135B,4);
TASK_PP(16'h135C,4);
TASK_PP(16'h135D,4);
TASK_PP(16'h135E,4);
TASK_PP(16'h135F,4);
TASK_PP(16'h1360,4);
TASK_PP(16'h1361,4);
TASK_PP(16'h1362,4);
TASK_PP(16'h1363,4);
TASK_PP(16'h1364,4);
TASK_PP(16'h1365,4);
TASK_PP(16'h1366,4);
TASK_PP(16'h1367,4);
TASK_PP(16'h1368,4);
TASK_PP(16'h1369,4);
TASK_PP(16'h136A,4);
TASK_PP(16'h136B,4);
TASK_PP(16'h136C,4);
TASK_PP(16'h136D,4);
TASK_PP(16'h136E,4);
TASK_PP(16'h136F,4);
TASK_PP(16'h1370,4);
TASK_PP(16'h1371,4);
TASK_PP(16'h1372,4);
TASK_PP(16'h1373,4);
TASK_PP(16'h1374,4);
TASK_PP(16'h1375,4);
TASK_PP(16'h1376,4);
TASK_PP(16'h1377,4);
TASK_PP(16'h1378,4);
TASK_PP(16'h1379,4);
TASK_PP(16'h137A,4);
TASK_PP(16'h137B,4);
TASK_PP(16'h137C,4);
TASK_PP(16'h137D,4);
TASK_PP(16'h137E,4);
TASK_PP(16'h137F,4);
TASK_PP(16'h1380,4);
TASK_PP(16'h1381,4);
TASK_PP(16'h1382,4);
TASK_PP(16'h1383,4);
TASK_PP(16'h1384,4);
TASK_PP(16'h1385,4);
TASK_PP(16'h1386,4);
TASK_PP(16'h1387,4);
TASK_PP(16'h1388,4);
TASK_PP(16'h1389,4);
TASK_PP(16'h138A,4);
TASK_PP(16'h138B,4);
TASK_PP(16'h138C,4);
TASK_PP(16'h138D,4);
TASK_PP(16'h138E,4);
TASK_PP(16'h138F,4);
TASK_PP(16'h1390,4);
TASK_PP(16'h1391,4);
TASK_PP(16'h1392,4);
TASK_PP(16'h1393,4);
TASK_PP(16'h1394,4);
TASK_PP(16'h1395,4);
TASK_PP(16'h1396,4);
TASK_PP(16'h1397,4);
TASK_PP(16'h1398,4);
TASK_PP(16'h1399,4);
TASK_PP(16'h139A,4);
TASK_PP(16'h139B,4);
TASK_PP(16'h139C,4);
TASK_PP(16'h139D,4);
TASK_PP(16'h139E,4);
TASK_PP(16'h139F,4);
TASK_PP(16'h13A0,4);
TASK_PP(16'h13A1,4);
TASK_PP(16'h13A2,4);
TASK_PP(16'h13A3,4);
TASK_PP(16'h13A4,4);
TASK_PP(16'h13A5,4);
TASK_PP(16'h13A6,4);
TASK_PP(16'h13A7,4);
TASK_PP(16'h13A8,4);
TASK_PP(16'h13A9,4);
TASK_PP(16'h13AA,4);
TASK_PP(16'h13AB,4);
TASK_PP(16'h13AC,4);
TASK_PP(16'h13AD,4);
TASK_PP(16'h13AE,4);
TASK_PP(16'h13AF,4);
TASK_PP(16'h13B0,4);
TASK_PP(16'h13B1,4);
TASK_PP(16'h13B2,4);
TASK_PP(16'h13B3,4);
TASK_PP(16'h13B4,4);
TASK_PP(16'h13B5,4);
TASK_PP(16'h13B6,4);
TASK_PP(16'h13B7,4);
TASK_PP(16'h13B8,4);
TASK_PP(16'h13B9,4);
TASK_PP(16'h13BA,4);
TASK_PP(16'h13BB,4);
TASK_PP(16'h13BC,4);
TASK_PP(16'h13BD,4);
TASK_PP(16'h13BE,4);
TASK_PP(16'h13BF,4);
TASK_PP(16'h13C0,4);
TASK_PP(16'h13C1,4);
TASK_PP(16'h13C2,4);
TASK_PP(16'h13C3,4);
TASK_PP(16'h13C4,4);
TASK_PP(16'h13C5,4);
TASK_PP(16'h13C6,4);
TASK_PP(16'h13C7,4);
TASK_PP(16'h13C8,4);
TASK_PP(16'h13C9,4);
TASK_PP(16'h13CA,4);
TASK_PP(16'h13CB,4);
TASK_PP(16'h13CC,4);
TASK_PP(16'h13CD,4);
TASK_PP(16'h13CE,4);
TASK_PP(16'h13CF,4);
TASK_PP(16'h13D0,4);
TASK_PP(16'h13D1,4);
TASK_PP(16'h13D2,4);
TASK_PP(16'h13D3,4);
TASK_PP(16'h13D4,4);
TASK_PP(16'h13D5,4);
TASK_PP(16'h13D6,4);
TASK_PP(16'h13D7,4);
TASK_PP(16'h13D8,4);
TASK_PP(16'h13D9,4);
TASK_PP(16'h13DA,4);
TASK_PP(16'h13DB,4);
TASK_PP(16'h13DC,4);
TASK_PP(16'h13DD,4);
TASK_PP(16'h13DE,4);
TASK_PP(16'h13DF,4);
TASK_PP(16'h13E0,4);
TASK_PP(16'h13E1,4);
TASK_PP(16'h13E2,4);
TASK_PP(16'h13E3,4);
TASK_PP(16'h13E4,4);
TASK_PP(16'h13E5,4);
TASK_PP(16'h13E6,4);
TASK_PP(16'h13E7,4);
TASK_PP(16'h13E8,4);
TASK_PP(16'h13E9,4);
TASK_PP(16'h13EA,4);
TASK_PP(16'h13EB,4);
TASK_PP(16'h13EC,4);
TASK_PP(16'h13ED,4);
TASK_PP(16'h13EE,4);
TASK_PP(16'h13EF,4);
TASK_PP(16'h13F0,4);
TASK_PP(16'h13F1,4);
TASK_PP(16'h13F2,4);
TASK_PP(16'h13F3,4);
TASK_PP(16'h13F4,4);
TASK_PP(16'h13F5,4);
TASK_PP(16'h13F6,4);
TASK_PP(16'h13F7,4);
TASK_PP(16'h13F8,4);
TASK_PP(16'h13F9,4);
TASK_PP(16'h13FA,4);
TASK_PP(16'h13FB,4);
TASK_PP(16'h13FC,4);
TASK_PP(16'h13FD,4);
TASK_PP(16'h13FE,4);
TASK_PP(16'h13FF,4);
TASK_PP(16'h1400,4);
TASK_PP(16'h1401,4);
TASK_PP(16'h1402,4);
TASK_PP(16'h1403,4);
TASK_PP(16'h1404,4);
TASK_PP(16'h1405,4);
TASK_PP(16'h1406,4);
TASK_PP(16'h1407,4);
TASK_PP(16'h1408,4);
TASK_PP(16'h1409,4);
TASK_PP(16'h140A,4);
TASK_PP(16'h140B,4);
TASK_PP(16'h140C,4);
TASK_PP(16'h140D,4);
TASK_PP(16'h140E,4);
TASK_PP(16'h140F,4);
TASK_PP(16'h1410,4);
TASK_PP(16'h1411,4);
TASK_PP(16'h1412,4);
TASK_PP(16'h1413,4);
TASK_PP(16'h1414,4);
TASK_PP(16'h1415,4);
TASK_PP(16'h1416,4);
TASK_PP(16'h1417,4);
TASK_PP(16'h1418,4);
TASK_PP(16'h1419,4);
TASK_PP(16'h141A,4);
TASK_PP(16'h141B,4);
TASK_PP(16'h141C,4);
TASK_PP(16'h141D,4);
TASK_PP(16'h141E,4);
TASK_PP(16'h141F,4);
TASK_PP(16'h1420,4);
TASK_PP(16'h1421,4);
TASK_PP(16'h1422,4);
TASK_PP(16'h1423,4);
TASK_PP(16'h1424,4);
TASK_PP(16'h1425,4);
TASK_PP(16'h1426,4);
TASK_PP(16'h1427,4);
TASK_PP(16'h1428,4);
TASK_PP(16'h1429,4);
TASK_PP(16'h142A,4);
TASK_PP(16'h142B,4);
TASK_PP(16'h142C,4);
TASK_PP(16'h142D,4);
TASK_PP(16'h142E,4);
TASK_PP(16'h142F,4);
TASK_PP(16'h1430,4);
TASK_PP(16'h1431,4);
TASK_PP(16'h1432,4);
TASK_PP(16'h1433,4);
TASK_PP(16'h1434,4);
TASK_PP(16'h1435,4);
TASK_PP(16'h1436,4);
TASK_PP(16'h1437,4);
TASK_PP(16'h1438,4);
TASK_PP(16'h1439,4);
TASK_PP(16'h143A,4);
TASK_PP(16'h143B,4);
TASK_PP(16'h143C,4);
TASK_PP(16'h143D,4);
TASK_PP(16'h143E,4);
TASK_PP(16'h143F,4);
TASK_PP(16'h1440,4);
TASK_PP(16'h1441,4);
TASK_PP(16'h1442,4);
TASK_PP(16'h1443,4);
TASK_PP(16'h1444,4);
TASK_PP(16'h1445,4);
TASK_PP(16'h1446,4);
TASK_PP(16'h1447,4);
TASK_PP(16'h1448,4);
TASK_PP(16'h1449,4);
TASK_PP(16'h144A,4);
TASK_PP(16'h144B,4);
TASK_PP(16'h144C,4);
TASK_PP(16'h144D,4);
TASK_PP(16'h144E,4);
TASK_PP(16'h144F,4);
TASK_PP(16'h1450,4);
TASK_PP(16'h1451,4);
TASK_PP(16'h1452,4);
TASK_PP(16'h1453,4);
TASK_PP(16'h1454,4);
TASK_PP(16'h1455,4);
TASK_PP(16'h1456,4);
TASK_PP(16'h1457,4);
TASK_PP(16'h1458,4);
TASK_PP(16'h1459,4);
TASK_PP(16'h145A,4);
TASK_PP(16'h145B,4);
TASK_PP(16'h145C,4);
TASK_PP(16'h145D,4);
TASK_PP(16'h145E,4);
TASK_PP(16'h145F,4);
TASK_PP(16'h1460,4);
TASK_PP(16'h1461,4);
TASK_PP(16'h1462,4);
TASK_PP(16'h1463,4);
TASK_PP(16'h1464,4);
TASK_PP(16'h1465,4);
TASK_PP(16'h1466,4);
TASK_PP(16'h1467,4);
TASK_PP(16'h1468,4);
TASK_PP(16'h1469,4);
TASK_PP(16'h146A,4);
TASK_PP(16'h146B,4);
TASK_PP(16'h146C,4);
TASK_PP(16'h146D,4);
TASK_PP(16'h146E,4);
TASK_PP(16'h146F,4);
TASK_PP(16'h1470,4);
TASK_PP(16'h1471,4);
TASK_PP(16'h1472,4);
TASK_PP(16'h1473,4);
TASK_PP(16'h1474,4);
TASK_PP(16'h1475,4);
TASK_PP(16'h1476,4);
TASK_PP(16'h1477,4);
TASK_PP(16'h1478,4);
TASK_PP(16'h1479,4);
TASK_PP(16'h147A,4);
TASK_PP(16'h147B,4);
TASK_PP(16'h147C,4);
TASK_PP(16'h147D,4);
TASK_PP(16'h147E,4);
TASK_PP(16'h147F,4);
TASK_PP(16'h1480,4);
TASK_PP(16'h1481,4);
TASK_PP(16'h1482,4);
TASK_PP(16'h1483,4);
TASK_PP(16'h1484,4);
TASK_PP(16'h1485,4);
TASK_PP(16'h1486,4);
TASK_PP(16'h1487,4);
TASK_PP(16'h1488,4);
TASK_PP(16'h1489,4);
TASK_PP(16'h148A,4);
TASK_PP(16'h148B,4);
TASK_PP(16'h148C,4);
TASK_PP(16'h148D,4);
TASK_PP(16'h148E,4);
TASK_PP(16'h148F,4);
TASK_PP(16'h1490,4);
TASK_PP(16'h1491,4);
TASK_PP(16'h1492,4);
TASK_PP(16'h1493,4);
TASK_PP(16'h1494,4);
TASK_PP(16'h1495,4);
TASK_PP(16'h1496,4);
TASK_PP(16'h1497,4);
TASK_PP(16'h1498,4);
TASK_PP(16'h1499,4);
TASK_PP(16'h149A,4);
TASK_PP(16'h149B,4);
TASK_PP(16'h149C,4);
TASK_PP(16'h149D,4);
TASK_PP(16'h149E,4);
TASK_PP(16'h149F,4);
TASK_PP(16'h14A0,4);
TASK_PP(16'h14A1,4);
TASK_PP(16'h14A2,4);
TASK_PP(16'h14A3,4);
TASK_PP(16'h14A4,4);
TASK_PP(16'h14A5,4);
TASK_PP(16'h14A6,4);
TASK_PP(16'h14A7,4);
TASK_PP(16'h14A8,4);
TASK_PP(16'h14A9,4);
TASK_PP(16'h14AA,4);
TASK_PP(16'h14AB,4);
TASK_PP(16'h14AC,4);
TASK_PP(16'h14AD,4);
TASK_PP(16'h14AE,4);
TASK_PP(16'h14AF,4);
TASK_PP(16'h14B0,4);
TASK_PP(16'h14B1,4);
TASK_PP(16'h14B2,4);
TASK_PP(16'h14B3,4);
TASK_PP(16'h14B4,4);
TASK_PP(16'h14B5,4);
TASK_PP(16'h14B6,4);
TASK_PP(16'h14B7,4);
TASK_PP(16'h14B8,4);
TASK_PP(16'h14B9,4);
TASK_PP(16'h14BA,4);
TASK_PP(16'h14BB,4);
TASK_PP(16'h14BC,4);
TASK_PP(16'h14BD,4);
TASK_PP(16'h14BE,4);
TASK_PP(16'h14BF,4);
TASK_PP(16'h14C0,4);
TASK_PP(16'h14C1,4);
TASK_PP(16'h14C2,4);
TASK_PP(16'h14C3,4);
TASK_PP(16'h14C4,4);
TASK_PP(16'h14C5,4);
TASK_PP(16'h14C6,4);
TASK_PP(16'h14C7,4);
TASK_PP(16'h14C8,4);
TASK_PP(16'h14C9,4);
TASK_PP(16'h14CA,4);
TASK_PP(16'h14CB,4);
TASK_PP(16'h14CC,4);
TASK_PP(16'h14CD,4);
TASK_PP(16'h14CE,4);
TASK_PP(16'h14CF,4);
TASK_PP(16'h14D0,4);
TASK_PP(16'h14D1,4);
TASK_PP(16'h14D2,4);
TASK_PP(16'h14D3,4);
TASK_PP(16'h14D4,4);
TASK_PP(16'h14D5,4);
TASK_PP(16'h14D6,4);
TASK_PP(16'h14D7,4);
TASK_PP(16'h14D8,4);
TASK_PP(16'h14D9,4);
TASK_PP(16'h14DA,4);
TASK_PP(16'h14DB,4);
TASK_PP(16'h14DC,4);
TASK_PP(16'h14DD,4);
TASK_PP(16'h14DE,4);
TASK_PP(16'h14DF,4);
TASK_PP(16'h14E0,4);
TASK_PP(16'h14E1,4);
TASK_PP(16'h14E2,4);
TASK_PP(16'h14E3,4);
TASK_PP(16'h14E4,4);
TASK_PP(16'h14E5,4);
TASK_PP(16'h14E6,4);
TASK_PP(16'h14E7,4);
TASK_PP(16'h14E8,4);
TASK_PP(16'h14E9,4);
TASK_PP(16'h14EA,4);
TASK_PP(16'h14EB,4);
TASK_PP(16'h14EC,4);
TASK_PP(16'h14ED,4);
TASK_PP(16'h14EE,4);
TASK_PP(16'h14EF,4);
TASK_PP(16'h14F0,4);
TASK_PP(16'h14F1,4);
TASK_PP(16'h14F2,4);
TASK_PP(16'h14F3,4);
TASK_PP(16'h14F4,4);
TASK_PP(16'h14F5,4);
TASK_PP(16'h14F6,4);
TASK_PP(16'h14F7,4);
TASK_PP(16'h14F8,4);
TASK_PP(16'h14F9,4);
TASK_PP(16'h14FA,4);
TASK_PP(16'h14FB,4);
TASK_PP(16'h14FC,4);
TASK_PP(16'h14FD,4);
TASK_PP(16'h14FE,4);
TASK_PP(16'h14FF,4);
TASK_PP(16'h1500,4);
TASK_PP(16'h1501,4);
TASK_PP(16'h1502,4);
TASK_PP(16'h1503,4);
TASK_PP(16'h1504,4);
TASK_PP(16'h1505,4);
TASK_PP(16'h1506,4);
TASK_PP(16'h1507,4);
TASK_PP(16'h1508,4);
TASK_PP(16'h1509,4);
TASK_PP(16'h150A,4);
TASK_PP(16'h150B,4);
TASK_PP(16'h150C,4);
TASK_PP(16'h150D,4);
TASK_PP(16'h150E,4);
TASK_PP(16'h150F,4);
TASK_PP(16'h1510,4);
TASK_PP(16'h1511,4);
TASK_PP(16'h1512,4);
TASK_PP(16'h1513,4);
TASK_PP(16'h1514,4);
TASK_PP(16'h1515,4);
TASK_PP(16'h1516,4);
TASK_PP(16'h1517,4);
TASK_PP(16'h1518,4);
TASK_PP(16'h1519,4);
TASK_PP(16'h151A,4);
TASK_PP(16'h151B,4);
TASK_PP(16'h151C,4);
TASK_PP(16'h151D,4);
TASK_PP(16'h151E,4);
TASK_PP(16'h151F,4);
TASK_PP(16'h1520,4);
TASK_PP(16'h1521,4);
TASK_PP(16'h1522,4);
TASK_PP(16'h1523,4);
TASK_PP(16'h1524,4);
TASK_PP(16'h1525,4);
TASK_PP(16'h1526,4);
TASK_PP(16'h1527,4);
TASK_PP(16'h1528,4);
TASK_PP(16'h1529,4);
TASK_PP(16'h152A,4);
TASK_PP(16'h152B,4);
TASK_PP(16'h152C,4);
TASK_PP(16'h152D,4);
TASK_PP(16'h152E,4);
TASK_PP(16'h152F,4);
TASK_PP(16'h1530,4);
TASK_PP(16'h1531,4);
TASK_PP(16'h1532,4);
TASK_PP(16'h1533,4);
TASK_PP(16'h1534,4);
TASK_PP(16'h1535,4);
TASK_PP(16'h1536,4);
TASK_PP(16'h1537,4);
TASK_PP(16'h1538,4);
TASK_PP(16'h1539,4);
TASK_PP(16'h153A,4);
TASK_PP(16'h153B,4);
TASK_PP(16'h153C,4);
TASK_PP(16'h153D,4);
TASK_PP(16'h153E,4);
TASK_PP(16'h153F,4);
TASK_PP(16'h1540,4);
TASK_PP(16'h1541,4);
TASK_PP(16'h1542,4);
TASK_PP(16'h1543,4);
TASK_PP(16'h1544,4);
TASK_PP(16'h1545,4);
TASK_PP(16'h1546,4);
TASK_PP(16'h1547,4);
TASK_PP(16'h1548,4);
TASK_PP(16'h1549,4);
TASK_PP(16'h154A,4);
TASK_PP(16'h154B,4);
TASK_PP(16'h154C,4);
TASK_PP(16'h154D,4);
TASK_PP(16'h154E,4);
TASK_PP(16'h154F,4);
TASK_PP(16'h1550,4);
TASK_PP(16'h1551,4);
TASK_PP(16'h1552,4);
TASK_PP(16'h1553,4);
TASK_PP(16'h1554,4);
TASK_PP(16'h1555,4);
TASK_PP(16'h1556,4);
TASK_PP(16'h1557,4);
TASK_PP(16'h1558,4);
TASK_PP(16'h1559,4);
TASK_PP(16'h155A,4);
TASK_PP(16'h155B,4);
TASK_PP(16'h155C,4);
TASK_PP(16'h155D,4);
TASK_PP(16'h155E,4);
TASK_PP(16'h155F,4);
TASK_PP(16'h1560,4);
TASK_PP(16'h1561,4);
TASK_PP(16'h1562,4);
TASK_PP(16'h1563,4);
TASK_PP(16'h1564,4);
TASK_PP(16'h1565,4);
TASK_PP(16'h1566,4);
TASK_PP(16'h1567,4);
TASK_PP(16'h1568,4);
TASK_PP(16'h1569,4);
TASK_PP(16'h156A,4);
TASK_PP(16'h156B,4);
TASK_PP(16'h156C,4);
TASK_PP(16'h156D,4);
TASK_PP(16'h156E,4);
TASK_PP(16'h156F,4);
TASK_PP(16'h1570,4);
TASK_PP(16'h1571,4);
TASK_PP(16'h1572,4);
TASK_PP(16'h1573,4);
TASK_PP(16'h1574,4);
TASK_PP(16'h1575,4);
TASK_PP(16'h1576,4);
TASK_PP(16'h1577,4);
TASK_PP(16'h1578,4);
TASK_PP(16'h1579,4);
TASK_PP(16'h157A,4);
TASK_PP(16'h157B,4);
TASK_PP(16'h157C,4);
TASK_PP(16'h157D,4);
TASK_PP(16'h157E,4);
TASK_PP(16'h157F,4);
TASK_PP(16'h1580,4);
TASK_PP(16'h1581,4);
TASK_PP(16'h1582,4);
TASK_PP(16'h1583,4);
TASK_PP(16'h1584,4);
TASK_PP(16'h1585,4);
TASK_PP(16'h1586,4);
TASK_PP(16'h1587,4);
TASK_PP(16'h1588,4);
TASK_PP(16'h1589,4);
TASK_PP(16'h158A,4);
TASK_PP(16'h158B,4);
TASK_PP(16'h158C,4);
TASK_PP(16'h158D,4);
TASK_PP(16'h158E,4);
TASK_PP(16'h158F,4);
TASK_PP(16'h1590,4);
TASK_PP(16'h1591,4);
TASK_PP(16'h1592,4);
TASK_PP(16'h1593,4);
TASK_PP(16'h1594,4);
TASK_PP(16'h1595,4);
TASK_PP(16'h1596,4);
TASK_PP(16'h1597,4);
TASK_PP(16'h1598,4);
TASK_PP(16'h1599,4);
TASK_PP(16'h159A,4);
TASK_PP(16'h159B,4);
TASK_PP(16'h159C,4);
TASK_PP(16'h159D,4);
TASK_PP(16'h159E,4);
TASK_PP(16'h159F,4);
TASK_PP(16'h15A0,4);
TASK_PP(16'h15A1,4);
TASK_PP(16'h15A2,4);
TASK_PP(16'h15A3,4);
TASK_PP(16'h15A4,4);
TASK_PP(16'h15A5,4);
TASK_PP(16'h15A6,4);
TASK_PP(16'h15A7,4);
TASK_PP(16'h15A8,4);
TASK_PP(16'h15A9,4);
TASK_PP(16'h15AA,4);
TASK_PP(16'h15AB,4);
TASK_PP(16'h15AC,4);
TASK_PP(16'h15AD,4);
TASK_PP(16'h15AE,4);
TASK_PP(16'h15AF,4);
TASK_PP(16'h15B0,4);
TASK_PP(16'h15B1,4);
TASK_PP(16'h15B2,4);
TASK_PP(16'h15B3,4);
TASK_PP(16'h15B4,4);
TASK_PP(16'h15B5,4);
TASK_PP(16'h15B6,4);
TASK_PP(16'h15B7,4);
TASK_PP(16'h15B8,4);
TASK_PP(16'h15B9,4);
TASK_PP(16'h15BA,4);
TASK_PP(16'h15BB,4);
TASK_PP(16'h15BC,4);
TASK_PP(16'h15BD,4);
TASK_PP(16'h15BE,4);
TASK_PP(16'h15BF,4);
TASK_PP(16'h15C0,4);
TASK_PP(16'h15C1,4);
TASK_PP(16'h15C2,4);
TASK_PP(16'h15C3,4);
TASK_PP(16'h15C4,4);
TASK_PP(16'h15C5,4);
TASK_PP(16'h15C6,4);
TASK_PP(16'h15C7,4);
TASK_PP(16'h15C8,4);
TASK_PP(16'h15C9,4);
TASK_PP(16'h15CA,4);
TASK_PP(16'h15CB,4);
TASK_PP(16'h15CC,4);
TASK_PP(16'h15CD,4);
TASK_PP(16'h15CE,4);
TASK_PP(16'h15CF,4);
TASK_PP(16'h15D0,4);
TASK_PP(16'h15D1,4);
TASK_PP(16'h15D2,4);
TASK_PP(16'h15D3,4);
TASK_PP(16'h15D4,4);
TASK_PP(16'h15D5,4);
TASK_PP(16'h15D6,4);
TASK_PP(16'h15D7,4);
TASK_PP(16'h15D8,4);
TASK_PP(16'h15D9,4);
TASK_PP(16'h15DA,4);
TASK_PP(16'h15DB,4);
TASK_PP(16'h15DC,4);
TASK_PP(16'h15DD,4);
TASK_PP(16'h15DE,4);
TASK_PP(16'h15DF,4);
TASK_PP(16'h15E0,4);
TASK_PP(16'h15E1,4);
TASK_PP(16'h15E2,4);
TASK_PP(16'h15E3,4);
TASK_PP(16'h15E4,4);
TASK_PP(16'h15E5,4);
TASK_PP(16'h15E6,4);
TASK_PP(16'h15E7,4);
TASK_PP(16'h15E8,4);
TASK_PP(16'h15E9,4);
TASK_PP(16'h15EA,4);
TASK_PP(16'h15EB,4);
TASK_PP(16'h15EC,4);
TASK_PP(16'h15ED,4);
TASK_PP(16'h15EE,4);
TASK_PP(16'h15EF,4);
TASK_PP(16'h15F0,4);
TASK_PP(16'h15F1,4);
TASK_PP(16'h15F2,4);
TASK_PP(16'h15F3,4);
TASK_PP(16'h15F4,4);
TASK_PP(16'h15F5,4);
TASK_PP(16'h15F6,4);
TASK_PP(16'h15F7,4);
TASK_PP(16'h15F8,4);
TASK_PP(16'h15F9,4);
TASK_PP(16'h15FA,4);
TASK_PP(16'h15FB,4);
TASK_PP(16'h15FC,4);
TASK_PP(16'h15FD,4);
TASK_PP(16'h15FE,4);
TASK_PP(16'h15FF,4);
TASK_PP(16'h1600,4);
TASK_PP(16'h1601,4);
TASK_PP(16'h1602,4);
TASK_PP(16'h1603,4);
TASK_PP(16'h1604,4);
TASK_PP(16'h1605,4);
TASK_PP(16'h1606,4);
TASK_PP(16'h1607,4);
TASK_PP(16'h1608,4);
TASK_PP(16'h1609,4);
TASK_PP(16'h160A,4);
TASK_PP(16'h160B,4);
TASK_PP(16'h160C,4);
TASK_PP(16'h160D,4);
TASK_PP(16'h160E,4);
TASK_PP(16'h160F,4);
TASK_PP(16'h1610,4);
TASK_PP(16'h1611,4);
TASK_PP(16'h1612,4);
TASK_PP(16'h1613,4);
TASK_PP(16'h1614,4);
TASK_PP(16'h1615,4);
TASK_PP(16'h1616,4);
TASK_PP(16'h1617,4);
TASK_PP(16'h1618,4);
TASK_PP(16'h1619,4);
TASK_PP(16'h161A,4);
TASK_PP(16'h161B,4);
TASK_PP(16'h161C,4);
TASK_PP(16'h161D,4);
TASK_PP(16'h161E,4);
TASK_PP(16'h161F,4);
TASK_PP(16'h1620,4);
TASK_PP(16'h1621,4);
TASK_PP(16'h1622,4);
TASK_PP(16'h1623,4);
TASK_PP(16'h1624,4);
TASK_PP(16'h1625,4);
TASK_PP(16'h1626,4);
TASK_PP(16'h1627,4);
TASK_PP(16'h1628,4);
TASK_PP(16'h1629,4);
TASK_PP(16'h162A,4);
TASK_PP(16'h162B,4);
TASK_PP(16'h162C,4);
TASK_PP(16'h162D,4);
TASK_PP(16'h162E,4);
TASK_PP(16'h162F,4);
TASK_PP(16'h1630,4);
TASK_PP(16'h1631,4);
TASK_PP(16'h1632,4);
TASK_PP(16'h1633,4);
TASK_PP(16'h1634,4);
TASK_PP(16'h1635,4);
TASK_PP(16'h1636,4);
TASK_PP(16'h1637,4);
TASK_PP(16'h1638,4);
TASK_PP(16'h1639,4);
TASK_PP(16'h163A,4);
TASK_PP(16'h163B,4);
TASK_PP(16'h163C,4);
TASK_PP(16'h163D,4);
TASK_PP(16'h163E,4);
TASK_PP(16'h163F,4);
TASK_PP(16'h1640,4);
TASK_PP(16'h1641,4);
TASK_PP(16'h1642,4);
TASK_PP(16'h1643,4);
TASK_PP(16'h1644,4);
TASK_PP(16'h1645,4);
TASK_PP(16'h1646,4);
TASK_PP(16'h1647,4);
TASK_PP(16'h1648,4);
TASK_PP(16'h1649,4);
TASK_PP(16'h164A,4);
TASK_PP(16'h164B,4);
TASK_PP(16'h164C,4);
TASK_PP(16'h164D,4);
TASK_PP(16'h164E,4);
TASK_PP(16'h164F,4);
TASK_PP(16'h1650,4);
TASK_PP(16'h1651,4);
TASK_PP(16'h1652,4);
TASK_PP(16'h1653,4);
TASK_PP(16'h1654,4);
TASK_PP(16'h1655,4);
TASK_PP(16'h1656,4);
TASK_PP(16'h1657,4);
TASK_PP(16'h1658,4);
TASK_PP(16'h1659,4);
TASK_PP(16'h165A,4);
TASK_PP(16'h165B,4);
TASK_PP(16'h165C,4);
TASK_PP(16'h165D,4);
TASK_PP(16'h165E,4);
TASK_PP(16'h165F,4);
TASK_PP(16'h1660,4);
TASK_PP(16'h1661,4);
TASK_PP(16'h1662,4);
TASK_PP(16'h1663,4);
TASK_PP(16'h1664,4);
TASK_PP(16'h1665,4);
TASK_PP(16'h1666,4);
TASK_PP(16'h1667,4);
TASK_PP(16'h1668,4);
TASK_PP(16'h1669,4);
TASK_PP(16'h166A,4);
TASK_PP(16'h166B,4);
TASK_PP(16'h166C,4);
TASK_PP(16'h166D,4);
TASK_PP(16'h166E,4);
TASK_PP(16'h166F,4);
TASK_PP(16'h1670,4);
TASK_PP(16'h1671,4);
TASK_PP(16'h1672,4);
TASK_PP(16'h1673,4);
TASK_PP(16'h1674,4);
TASK_PP(16'h1675,4);
TASK_PP(16'h1676,4);
TASK_PP(16'h1677,4);
TASK_PP(16'h1678,4);
TASK_PP(16'h1679,4);
TASK_PP(16'h167A,4);
TASK_PP(16'h167B,4);
TASK_PP(16'h167C,4);
TASK_PP(16'h167D,4);
TASK_PP(16'h167E,4);
TASK_PP(16'h167F,4);
TASK_PP(16'h1680,4);
TASK_PP(16'h1681,4);
TASK_PP(16'h1682,4);
TASK_PP(16'h1683,4);
TASK_PP(16'h1684,4);
TASK_PP(16'h1685,4);
TASK_PP(16'h1686,4);
TASK_PP(16'h1687,4);
TASK_PP(16'h1688,4);
TASK_PP(16'h1689,4);
TASK_PP(16'h168A,4);
TASK_PP(16'h168B,4);
TASK_PP(16'h168C,4);
TASK_PP(16'h168D,4);
TASK_PP(16'h168E,4);
TASK_PP(16'h168F,4);
TASK_PP(16'h1690,4);
TASK_PP(16'h1691,4);
TASK_PP(16'h1692,4);
TASK_PP(16'h1693,4);
TASK_PP(16'h1694,4);
TASK_PP(16'h1695,4);
TASK_PP(16'h1696,4);
TASK_PP(16'h1697,4);
TASK_PP(16'h1698,4);
TASK_PP(16'h1699,4);
TASK_PP(16'h169A,4);
TASK_PP(16'h169B,4);
TASK_PP(16'h169C,4);
TASK_PP(16'h169D,4);
TASK_PP(16'h169E,4);
TASK_PP(16'h169F,4);
TASK_PP(16'h16A0,4);
TASK_PP(16'h16A1,4);
TASK_PP(16'h16A2,4);
TASK_PP(16'h16A3,4);
TASK_PP(16'h16A4,4);
TASK_PP(16'h16A5,4);
TASK_PP(16'h16A6,4);
TASK_PP(16'h16A7,4);
TASK_PP(16'h16A8,4);
TASK_PP(16'h16A9,4);
TASK_PP(16'h16AA,4);
TASK_PP(16'h16AB,4);
TASK_PP(16'h16AC,4);
TASK_PP(16'h16AD,4);
TASK_PP(16'h16AE,4);
TASK_PP(16'h16AF,4);
TASK_PP(16'h16B0,4);
TASK_PP(16'h16B1,4);
TASK_PP(16'h16B2,4);
TASK_PP(16'h16B3,4);
TASK_PP(16'h16B4,4);
TASK_PP(16'h16B5,4);
TASK_PP(16'h16B6,4);
TASK_PP(16'h16B7,4);
TASK_PP(16'h16B8,4);
TASK_PP(16'h16B9,4);
TASK_PP(16'h16BA,4);
TASK_PP(16'h16BB,4);
TASK_PP(16'h16BC,4);
TASK_PP(16'h16BD,4);
TASK_PP(16'h16BE,4);
TASK_PP(16'h16BF,4);
TASK_PP(16'h16C0,4);
TASK_PP(16'h16C1,4);
TASK_PP(16'h16C2,4);
TASK_PP(16'h16C3,4);
TASK_PP(16'h16C4,4);
TASK_PP(16'h16C5,4);
TASK_PP(16'h16C6,4);
TASK_PP(16'h16C7,4);
TASK_PP(16'h16C8,4);
TASK_PP(16'h16C9,4);
TASK_PP(16'h16CA,4);
TASK_PP(16'h16CB,4);
TASK_PP(16'h16CC,4);
TASK_PP(16'h16CD,4);
TASK_PP(16'h16CE,4);
TASK_PP(16'h16CF,4);
TASK_PP(16'h16D0,4);
TASK_PP(16'h16D1,4);
TASK_PP(16'h16D2,4);
TASK_PP(16'h16D3,4);
TASK_PP(16'h16D4,4);
TASK_PP(16'h16D5,4);
TASK_PP(16'h16D6,4);
TASK_PP(16'h16D7,4);
TASK_PP(16'h16D8,4);
TASK_PP(16'h16D9,4);
TASK_PP(16'h16DA,4);
TASK_PP(16'h16DB,4);
TASK_PP(16'h16DC,4);
TASK_PP(16'h16DD,4);
TASK_PP(16'h16DE,4);
TASK_PP(16'h16DF,4);
TASK_PP(16'h16E0,4);
TASK_PP(16'h16E1,4);
TASK_PP(16'h16E2,4);
TASK_PP(16'h16E3,4);
TASK_PP(16'h16E4,4);
TASK_PP(16'h16E5,4);
TASK_PP(16'h16E6,4);
TASK_PP(16'h16E7,4);
TASK_PP(16'h16E8,4);
TASK_PP(16'h16E9,4);
TASK_PP(16'h16EA,4);
TASK_PP(16'h16EB,4);
TASK_PP(16'h16EC,4);
TASK_PP(16'h16ED,4);
TASK_PP(16'h16EE,4);
TASK_PP(16'h16EF,4);
TASK_PP(16'h16F0,4);
TASK_PP(16'h16F1,4);
TASK_PP(16'h16F2,4);
TASK_PP(16'h16F3,4);
TASK_PP(16'h16F4,4);
TASK_PP(16'h16F5,4);
TASK_PP(16'h16F6,4);
TASK_PP(16'h16F7,4);
TASK_PP(16'h16F8,4);
TASK_PP(16'h16F9,4);
TASK_PP(16'h16FA,4);
TASK_PP(16'h16FB,4);
TASK_PP(16'h16FC,4);
TASK_PP(16'h16FD,4);
TASK_PP(16'h16FE,4);
TASK_PP(16'h16FF,4);
TASK_PP(16'h1700,4);
TASK_PP(16'h1701,4);
TASK_PP(16'h1702,4);
TASK_PP(16'h1703,4);
TASK_PP(16'h1704,4);
TASK_PP(16'h1705,4);
TASK_PP(16'h1706,4);
TASK_PP(16'h1707,4);
TASK_PP(16'h1708,4);
TASK_PP(16'h1709,4);
TASK_PP(16'h170A,4);
TASK_PP(16'h170B,4);
TASK_PP(16'h170C,4);
TASK_PP(16'h170D,4);
TASK_PP(16'h170E,4);
TASK_PP(16'h170F,4);
TASK_PP(16'h1710,4);
TASK_PP(16'h1711,4);
TASK_PP(16'h1712,4);
TASK_PP(16'h1713,4);
TASK_PP(16'h1714,4);
TASK_PP(16'h1715,4);
TASK_PP(16'h1716,4);
TASK_PP(16'h1717,4);
TASK_PP(16'h1718,4);
TASK_PP(16'h1719,4);
TASK_PP(16'h171A,4);
TASK_PP(16'h171B,4);
TASK_PP(16'h171C,4);
TASK_PP(16'h171D,4);
TASK_PP(16'h171E,4);
TASK_PP(16'h171F,4);
TASK_PP(16'h1720,4);
TASK_PP(16'h1721,4);
TASK_PP(16'h1722,4);
TASK_PP(16'h1723,4);
TASK_PP(16'h1724,4);
TASK_PP(16'h1725,4);
TASK_PP(16'h1726,4);
TASK_PP(16'h1727,4);
TASK_PP(16'h1728,4);
TASK_PP(16'h1729,4);
TASK_PP(16'h172A,4);
TASK_PP(16'h172B,4);
TASK_PP(16'h172C,4);
TASK_PP(16'h172D,4);
TASK_PP(16'h172E,4);
TASK_PP(16'h172F,4);
TASK_PP(16'h1730,4);
TASK_PP(16'h1731,4);
TASK_PP(16'h1732,4);
TASK_PP(16'h1733,4);
TASK_PP(16'h1734,4);
TASK_PP(16'h1735,4);
TASK_PP(16'h1736,4);
TASK_PP(16'h1737,4);
TASK_PP(16'h1738,4);
TASK_PP(16'h1739,4);
TASK_PP(16'h173A,4);
TASK_PP(16'h173B,4);
TASK_PP(16'h173C,4);
TASK_PP(16'h173D,4);
TASK_PP(16'h173E,4);
TASK_PP(16'h173F,4);
TASK_PP(16'h1740,4);
TASK_PP(16'h1741,4);
TASK_PP(16'h1742,4);
TASK_PP(16'h1743,4);
TASK_PP(16'h1744,4);
TASK_PP(16'h1745,4);
TASK_PP(16'h1746,4);
TASK_PP(16'h1747,4);
TASK_PP(16'h1748,4);
TASK_PP(16'h1749,4);
TASK_PP(16'h174A,4);
TASK_PP(16'h174B,4);
TASK_PP(16'h174C,4);
TASK_PP(16'h174D,4);
TASK_PP(16'h174E,4);
TASK_PP(16'h174F,4);
TASK_PP(16'h1750,4);
TASK_PP(16'h1751,4);
TASK_PP(16'h1752,4);
TASK_PP(16'h1753,4);
TASK_PP(16'h1754,4);
TASK_PP(16'h1755,4);
TASK_PP(16'h1756,4);
TASK_PP(16'h1757,4);
TASK_PP(16'h1758,4);
TASK_PP(16'h1759,4);
TASK_PP(16'h175A,4);
TASK_PP(16'h175B,4);
TASK_PP(16'h175C,4);
TASK_PP(16'h175D,4);
TASK_PP(16'h175E,4);
TASK_PP(16'h175F,4);
TASK_PP(16'h1760,4);
TASK_PP(16'h1761,4);
TASK_PP(16'h1762,4);
TASK_PP(16'h1763,4);
TASK_PP(16'h1764,4);
TASK_PP(16'h1765,4);
TASK_PP(16'h1766,4);
TASK_PP(16'h1767,4);
TASK_PP(16'h1768,4);
TASK_PP(16'h1769,4);
TASK_PP(16'h176A,4);
TASK_PP(16'h176B,4);
TASK_PP(16'h176C,4);
TASK_PP(16'h176D,4);
TASK_PP(16'h176E,4);
TASK_PP(16'h176F,4);
TASK_PP(16'h1770,4);
TASK_PP(16'h1771,4);
TASK_PP(16'h1772,4);
TASK_PP(16'h1773,4);
TASK_PP(16'h1774,4);
TASK_PP(16'h1775,4);
TASK_PP(16'h1776,4);
TASK_PP(16'h1777,4);
TASK_PP(16'h1778,4);
TASK_PP(16'h1779,4);
TASK_PP(16'h177A,4);
TASK_PP(16'h177B,4);
TASK_PP(16'h177C,4);
TASK_PP(16'h177D,4);
TASK_PP(16'h177E,4);
TASK_PP(16'h177F,4);
TASK_PP(16'h1780,4);
TASK_PP(16'h1781,4);
TASK_PP(16'h1782,4);
TASK_PP(16'h1783,4);
TASK_PP(16'h1784,4);
TASK_PP(16'h1785,4);
TASK_PP(16'h1786,4);
TASK_PP(16'h1787,4);
TASK_PP(16'h1788,4);
TASK_PP(16'h1789,4);
TASK_PP(16'h178A,4);
TASK_PP(16'h178B,4);
TASK_PP(16'h178C,4);
TASK_PP(16'h178D,4);
TASK_PP(16'h178E,4);
TASK_PP(16'h178F,4);
TASK_PP(16'h1790,4);
TASK_PP(16'h1791,4);
TASK_PP(16'h1792,4);
TASK_PP(16'h1793,4);
TASK_PP(16'h1794,4);
TASK_PP(16'h1795,4);
TASK_PP(16'h1796,4);
TASK_PP(16'h1797,4);
TASK_PP(16'h1798,4);
TASK_PP(16'h1799,4);
TASK_PP(16'h179A,4);
TASK_PP(16'h179B,4);
TASK_PP(16'h179C,4);
TASK_PP(16'h179D,4);
TASK_PP(16'h179E,4);
TASK_PP(16'h179F,4);
TASK_PP(16'h17A0,4);
TASK_PP(16'h17A1,4);
TASK_PP(16'h17A2,4);
TASK_PP(16'h17A3,4);
TASK_PP(16'h17A4,4);
TASK_PP(16'h17A5,4);
TASK_PP(16'h17A6,4);
TASK_PP(16'h17A7,4);
TASK_PP(16'h17A8,4);
TASK_PP(16'h17A9,4);
TASK_PP(16'h17AA,4);
TASK_PP(16'h17AB,4);
TASK_PP(16'h17AC,4);
TASK_PP(16'h17AD,4);
TASK_PP(16'h17AE,4);
TASK_PP(16'h17AF,4);
TASK_PP(16'h17B0,4);
TASK_PP(16'h17B1,4);
TASK_PP(16'h17B2,4);
TASK_PP(16'h17B3,4);
TASK_PP(16'h17B4,4);
TASK_PP(16'h17B5,4);
TASK_PP(16'h17B6,4);
TASK_PP(16'h17B7,4);
TASK_PP(16'h17B8,4);
TASK_PP(16'h17B9,4);
TASK_PP(16'h17BA,4);
TASK_PP(16'h17BB,4);
TASK_PP(16'h17BC,4);
TASK_PP(16'h17BD,4);
TASK_PP(16'h17BE,4);
TASK_PP(16'h17BF,4);
TASK_PP(16'h17C0,4);
TASK_PP(16'h17C1,4);
TASK_PP(16'h17C2,4);
TASK_PP(16'h17C3,4);
TASK_PP(16'h17C4,4);
TASK_PP(16'h17C5,4);
TASK_PP(16'h17C6,4);
TASK_PP(16'h17C7,4);
TASK_PP(16'h17C8,4);
TASK_PP(16'h17C9,4);
TASK_PP(16'h17CA,4);
TASK_PP(16'h17CB,4);
TASK_PP(16'h17CC,4);
TASK_PP(16'h17CD,4);
TASK_PP(16'h17CE,4);
TASK_PP(16'h17CF,4);
TASK_PP(16'h17D0,4);
TASK_PP(16'h17D1,4);
TASK_PP(16'h17D2,4);
TASK_PP(16'h17D3,4);
TASK_PP(16'h17D4,4);
TASK_PP(16'h17D5,4);
TASK_PP(16'h17D6,4);
TASK_PP(16'h17D7,4);
TASK_PP(16'h17D8,4);
TASK_PP(16'h17D9,4);
TASK_PP(16'h17DA,4);
TASK_PP(16'h17DB,4);
TASK_PP(16'h17DC,4);
TASK_PP(16'h17DD,4);
TASK_PP(16'h17DE,4);
TASK_PP(16'h17DF,4);
TASK_PP(16'h17E0,4);
TASK_PP(16'h17E1,4);
TASK_PP(16'h17E2,4);
TASK_PP(16'h17E3,4);
TASK_PP(16'h17E4,4);
TASK_PP(16'h17E5,4);
TASK_PP(16'h17E6,4);
TASK_PP(16'h17E7,4);
TASK_PP(16'h17E8,4);
TASK_PP(16'h17E9,4);
TASK_PP(16'h17EA,4);
TASK_PP(16'h17EB,4);
TASK_PP(16'h17EC,4);
TASK_PP(16'h17ED,4);
TASK_PP(16'h17EE,4);
TASK_PP(16'h17EF,4);
TASK_PP(16'h17F0,4);
TASK_PP(16'h17F1,4);
TASK_PP(16'h17F2,4);
TASK_PP(16'h17F3,4);
TASK_PP(16'h17F4,4);
TASK_PP(16'h17F5,4);
TASK_PP(16'h17F6,4);
TASK_PP(16'h17F7,4);
TASK_PP(16'h17F8,4);
TASK_PP(16'h17F9,4);
TASK_PP(16'h17FA,4);
TASK_PP(16'h17FB,4);
TASK_PP(16'h17FC,4);
TASK_PP(16'h17FD,4);
TASK_PP(16'h17FE,4);
TASK_PP(16'h17FF,4);
TASK_PP(16'h1800,4);
TASK_PP(16'h1801,4);
TASK_PP(16'h1802,4);
TASK_PP(16'h1803,4);
TASK_PP(16'h1804,4);
TASK_PP(16'h1805,4);
TASK_PP(16'h1806,4);
TASK_PP(16'h1807,4);
TASK_PP(16'h1808,4);
TASK_PP(16'h1809,4);
TASK_PP(16'h180A,4);
TASK_PP(16'h180B,4);
TASK_PP(16'h180C,4);
TASK_PP(16'h180D,4);
TASK_PP(16'h180E,4);
TASK_PP(16'h180F,4);
TASK_PP(16'h1810,4);
TASK_PP(16'h1811,4);
TASK_PP(16'h1812,4);
TASK_PP(16'h1813,4);
TASK_PP(16'h1814,4);
TASK_PP(16'h1815,4);
TASK_PP(16'h1816,4);
TASK_PP(16'h1817,4);
TASK_PP(16'h1818,4);
TASK_PP(16'h1819,4);
TASK_PP(16'h181A,4);
TASK_PP(16'h181B,4);
TASK_PP(16'h181C,4);
TASK_PP(16'h181D,4);
TASK_PP(16'h181E,4);
TASK_PP(16'h181F,4);
TASK_PP(16'h1820,4);
TASK_PP(16'h1821,4);
TASK_PP(16'h1822,4);
TASK_PP(16'h1823,4);
TASK_PP(16'h1824,4);
TASK_PP(16'h1825,4);
TASK_PP(16'h1826,4);
TASK_PP(16'h1827,4);
TASK_PP(16'h1828,4);
TASK_PP(16'h1829,4);
TASK_PP(16'h182A,4);
TASK_PP(16'h182B,4);
TASK_PP(16'h182C,4);
TASK_PP(16'h182D,4);
TASK_PP(16'h182E,4);
TASK_PP(16'h182F,4);
TASK_PP(16'h1830,4);
TASK_PP(16'h1831,4);
TASK_PP(16'h1832,4);
TASK_PP(16'h1833,4);
TASK_PP(16'h1834,4);
TASK_PP(16'h1835,4);
TASK_PP(16'h1836,4);
TASK_PP(16'h1837,4);
TASK_PP(16'h1838,4);
TASK_PP(16'h1839,4);
TASK_PP(16'h183A,4);
TASK_PP(16'h183B,4);
TASK_PP(16'h183C,4);
TASK_PP(16'h183D,4);
TASK_PP(16'h183E,4);
TASK_PP(16'h183F,4);
TASK_PP(16'h1840,4);
TASK_PP(16'h1841,4);
TASK_PP(16'h1842,4);
TASK_PP(16'h1843,4);
TASK_PP(16'h1844,4);
TASK_PP(16'h1845,4);
TASK_PP(16'h1846,4);
TASK_PP(16'h1847,4);
TASK_PP(16'h1848,4);
TASK_PP(16'h1849,4);
TASK_PP(16'h184A,4);
TASK_PP(16'h184B,4);
TASK_PP(16'h184C,4);
TASK_PP(16'h184D,4);
TASK_PP(16'h184E,4);
TASK_PP(16'h184F,4);
TASK_PP(16'h1850,4);
TASK_PP(16'h1851,4);
TASK_PP(16'h1852,4);
TASK_PP(16'h1853,4);
TASK_PP(16'h1854,4);
TASK_PP(16'h1855,4);
TASK_PP(16'h1856,4);
TASK_PP(16'h1857,4);
TASK_PP(16'h1858,4);
TASK_PP(16'h1859,4);
TASK_PP(16'h185A,4);
TASK_PP(16'h185B,4);
TASK_PP(16'h185C,4);
TASK_PP(16'h185D,4);
TASK_PP(16'h185E,4);
TASK_PP(16'h185F,4);
TASK_PP(16'h1860,4);
TASK_PP(16'h1861,4);
TASK_PP(16'h1862,4);
TASK_PP(16'h1863,4);
TASK_PP(16'h1864,4);
TASK_PP(16'h1865,4);
TASK_PP(16'h1866,4);
TASK_PP(16'h1867,4);
TASK_PP(16'h1868,4);
TASK_PP(16'h1869,4);
TASK_PP(16'h186A,4);
TASK_PP(16'h186B,4);
TASK_PP(16'h186C,4);
TASK_PP(16'h186D,4);
TASK_PP(16'h186E,4);
TASK_PP(16'h186F,4);
TASK_PP(16'h1870,4);
TASK_PP(16'h1871,4);
TASK_PP(16'h1872,4);
TASK_PP(16'h1873,4);
TASK_PP(16'h1874,4);
TASK_PP(16'h1875,4);
TASK_PP(16'h1876,4);
TASK_PP(16'h1877,4);
TASK_PP(16'h1878,4);
TASK_PP(16'h1879,4);
TASK_PP(16'h187A,4);
TASK_PP(16'h187B,4);
TASK_PP(16'h187C,4);
TASK_PP(16'h187D,4);
TASK_PP(16'h187E,4);
TASK_PP(16'h187F,4);
TASK_PP(16'h1880,4);
TASK_PP(16'h1881,4);
TASK_PP(16'h1882,4);
TASK_PP(16'h1883,4);
TASK_PP(16'h1884,4);
TASK_PP(16'h1885,4);
TASK_PP(16'h1886,4);
TASK_PP(16'h1887,4);
TASK_PP(16'h1888,4);
TASK_PP(16'h1889,4);
TASK_PP(16'h188A,4);
TASK_PP(16'h188B,4);
TASK_PP(16'h188C,4);
TASK_PP(16'h188D,4);
TASK_PP(16'h188E,4);
TASK_PP(16'h188F,4);
TASK_PP(16'h1890,4);
TASK_PP(16'h1891,4);
TASK_PP(16'h1892,4);
TASK_PP(16'h1893,4);
TASK_PP(16'h1894,4);
TASK_PP(16'h1895,4);
TASK_PP(16'h1896,4);
TASK_PP(16'h1897,4);
TASK_PP(16'h1898,4);
TASK_PP(16'h1899,4);
TASK_PP(16'h189A,4);
TASK_PP(16'h189B,4);
TASK_PP(16'h189C,4);
TASK_PP(16'h189D,4);
TASK_PP(16'h189E,4);
TASK_PP(16'h189F,4);
TASK_PP(16'h18A0,4);
TASK_PP(16'h18A1,4);
TASK_PP(16'h18A2,4);
TASK_PP(16'h18A3,4);
TASK_PP(16'h18A4,4);
TASK_PP(16'h18A5,4);
TASK_PP(16'h18A6,4);
TASK_PP(16'h18A7,4);
TASK_PP(16'h18A8,4);
TASK_PP(16'h18A9,4);
TASK_PP(16'h18AA,4);
TASK_PP(16'h18AB,4);
TASK_PP(16'h18AC,4);
TASK_PP(16'h18AD,4);
TASK_PP(16'h18AE,4);
TASK_PP(16'h18AF,4);
TASK_PP(16'h18B0,4);
TASK_PP(16'h18B1,4);
TASK_PP(16'h18B2,4);
TASK_PP(16'h18B3,4);
TASK_PP(16'h18B4,4);
TASK_PP(16'h18B5,4);
TASK_PP(16'h18B6,4);
TASK_PP(16'h18B7,4);
TASK_PP(16'h18B8,4);
TASK_PP(16'h18B9,4);
TASK_PP(16'h18BA,4);
TASK_PP(16'h18BB,4);
TASK_PP(16'h18BC,4);
TASK_PP(16'h18BD,4);
TASK_PP(16'h18BE,4);
TASK_PP(16'h18BF,4);
TASK_PP(16'h18C0,4);
TASK_PP(16'h18C1,4);
TASK_PP(16'h18C2,4);
TASK_PP(16'h18C3,4);
TASK_PP(16'h18C4,4);
TASK_PP(16'h18C5,4);
TASK_PP(16'h18C6,4);
TASK_PP(16'h18C7,4);
TASK_PP(16'h18C8,4);
TASK_PP(16'h18C9,4);
TASK_PP(16'h18CA,4);
TASK_PP(16'h18CB,4);
TASK_PP(16'h18CC,4);
TASK_PP(16'h18CD,4);
TASK_PP(16'h18CE,4);
TASK_PP(16'h18CF,4);
TASK_PP(16'h18D0,4);
TASK_PP(16'h18D1,4);
TASK_PP(16'h18D2,4);
TASK_PP(16'h18D3,4);
TASK_PP(16'h18D4,4);
TASK_PP(16'h18D5,4);
TASK_PP(16'h18D6,4);
TASK_PP(16'h18D7,4);
TASK_PP(16'h18D8,4);
TASK_PP(16'h18D9,4);
TASK_PP(16'h18DA,4);
TASK_PP(16'h18DB,4);
TASK_PP(16'h18DC,4);
TASK_PP(16'h18DD,4);
TASK_PP(16'h18DE,4);
TASK_PP(16'h18DF,4);
TASK_PP(16'h18E0,4);
TASK_PP(16'h18E1,4);
TASK_PP(16'h18E2,4);
TASK_PP(16'h18E3,4);
TASK_PP(16'h18E4,4);
TASK_PP(16'h18E5,4);
TASK_PP(16'h18E6,4);
TASK_PP(16'h18E7,4);
TASK_PP(16'h18E8,4);
TASK_PP(16'h18E9,4);
TASK_PP(16'h18EA,4);
TASK_PP(16'h18EB,4);
TASK_PP(16'h18EC,4);
TASK_PP(16'h18ED,4);
TASK_PP(16'h18EE,4);
TASK_PP(16'h18EF,4);
TASK_PP(16'h18F0,4);
TASK_PP(16'h18F1,4);
TASK_PP(16'h18F2,4);
TASK_PP(16'h18F3,4);
TASK_PP(16'h18F4,4);
TASK_PP(16'h18F5,4);
TASK_PP(16'h18F6,4);
TASK_PP(16'h18F7,4);
TASK_PP(16'h18F8,4);
TASK_PP(16'h18F9,4);
TASK_PP(16'h18FA,4);
TASK_PP(16'h18FB,4);
TASK_PP(16'h18FC,4);
TASK_PP(16'h18FD,4);
TASK_PP(16'h18FE,4);
TASK_PP(16'h18FF,4);
TASK_PP(16'h1900,4);
TASK_PP(16'h1901,4);
TASK_PP(16'h1902,4);
TASK_PP(16'h1903,4);
TASK_PP(16'h1904,4);
TASK_PP(16'h1905,4);
TASK_PP(16'h1906,4);
TASK_PP(16'h1907,4);
TASK_PP(16'h1908,4);
TASK_PP(16'h1909,4);
TASK_PP(16'h190A,4);
TASK_PP(16'h190B,4);
TASK_PP(16'h190C,4);
TASK_PP(16'h190D,4);
TASK_PP(16'h190E,4);
TASK_PP(16'h190F,4);
TASK_PP(16'h1910,4);
TASK_PP(16'h1911,4);
TASK_PP(16'h1912,4);
TASK_PP(16'h1913,4);
TASK_PP(16'h1914,4);
TASK_PP(16'h1915,4);
TASK_PP(16'h1916,4);
TASK_PP(16'h1917,4);
TASK_PP(16'h1918,4);
TASK_PP(16'h1919,4);
TASK_PP(16'h191A,4);
TASK_PP(16'h191B,4);
TASK_PP(16'h191C,4);
TASK_PP(16'h191D,4);
TASK_PP(16'h191E,4);
TASK_PP(16'h191F,4);
TASK_PP(16'h1920,4);
TASK_PP(16'h1921,4);
TASK_PP(16'h1922,4);
TASK_PP(16'h1923,4);
TASK_PP(16'h1924,4);
TASK_PP(16'h1925,4);
TASK_PP(16'h1926,4);
TASK_PP(16'h1927,4);
TASK_PP(16'h1928,4);
TASK_PP(16'h1929,4);
TASK_PP(16'h192A,4);
TASK_PP(16'h192B,4);
TASK_PP(16'h192C,4);
TASK_PP(16'h192D,4);
TASK_PP(16'h192E,4);
TASK_PP(16'h192F,4);
TASK_PP(16'h1930,4);
TASK_PP(16'h1931,4);
TASK_PP(16'h1932,4);
TASK_PP(16'h1933,4);
TASK_PP(16'h1934,4);
TASK_PP(16'h1935,4);
TASK_PP(16'h1936,4);
TASK_PP(16'h1937,4);
TASK_PP(16'h1938,4);
TASK_PP(16'h1939,4);
TASK_PP(16'h193A,4);
TASK_PP(16'h193B,4);
TASK_PP(16'h193C,4);
TASK_PP(16'h193D,4);
TASK_PP(16'h193E,4);
TASK_PP(16'h193F,4);
TASK_PP(16'h1940,4);
TASK_PP(16'h1941,4);
TASK_PP(16'h1942,4);
TASK_PP(16'h1943,4);
TASK_PP(16'h1944,4);
TASK_PP(16'h1945,4);
TASK_PP(16'h1946,4);
TASK_PP(16'h1947,4);
TASK_PP(16'h1948,4);
TASK_PP(16'h1949,4);
TASK_PP(16'h194A,4);
TASK_PP(16'h194B,4);
TASK_PP(16'h194C,4);
TASK_PP(16'h194D,4);
TASK_PP(16'h194E,4);
TASK_PP(16'h194F,4);
TASK_PP(16'h1950,4);
TASK_PP(16'h1951,4);
TASK_PP(16'h1952,4);
TASK_PP(16'h1953,4);
TASK_PP(16'h1954,4);
TASK_PP(16'h1955,4);
TASK_PP(16'h1956,4);
TASK_PP(16'h1957,4);
TASK_PP(16'h1958,4);
TASK_PP(16'h1959,4);
TASK_PP(16'h195A,4);
TASK_PP(16'h195B,4);
TASK_PP(16'h195C,4);
TASK_PP(16'h195D,4);
TASK_PP(16'h195E,4);
TASK_PP(16'h195F,4);
TASK_PP(16'h1960,4);
TASK_PP(16'h1961,4);
TASK_PP(16'h1962,4);
TASK_PP(16'h1963,4);
TASK_PP(16'h1964,4);
TASK_PP(16'h1965,4);
TASK_PP(16'h1966,4);
TASK_PP(16'h1967,4);
TASK_PP(16'h1968,4);
TASK_PP(16'h1969,4);
TASK_PP(16'h196A,4);
TASK_PP(16'h196B,4);
TASK_PP(16'h196C,4);
TASK_PP(16'h196D,4);
TASK_PP(16'h196E,4);
TASK_PP(16'h196F,4);
TASK_PP(16'h1970,4);
TASK_PP(16'h1971,4);
TASK_PP(16'h1972,4);
TASK_PP(16'h1973,4);
TASK_PP(16'h1974,4);
TASK_PP(16'h1975,4);
TASK_PP(16'h1976,4);
TASK_PP(16'h1977,4);
TASK_PP(16'h1978,4);
TASK_PP(16'h1979,4);
TASK_PP(16'h197A,4);
TASK_PP(16'h197B,4);
TASK_PP(16'h197C,4);
TASK_PP(16'h197D,4);
TASK_PP(16'h197E,4);
TASK_PP(16'h197F,4);
TASK_PP(16'h1980,4);
TASK_PP(16'h1981,4);
TASK_PP(16'h1982,4);
TASK_PP(16'h1983,4);
TASK_PP(16'h1984,4);
TASK_PP(16'h1985,4);
TASK_PP(16'h1986,4);
TASK_PP(16'h1987,4);
TASK_PP(16'h1988,4);
TASK_PP(16'h1989,4);
TASK_PP(16'h198A,4);
TASK_PP(16'h198B,4);
TASK_PP(16'h198C,4);
TASK_PP(16'h198D,4);
TASK_PP(16'h198E,4);
TASK_PP(16'h198F,4);
TASK_PP(16'h1990,4);
TASK_PP(16'h1991,4);
TASK_PP(16'h1992,4);
TASK_PP(16'h1993,4);
TASK_PP(16'h1994,4);
TASK_PP(16'h1995,4);
TASK_PP(16'h1996,4);
TASK_PP(16'h1997,4);
TASK_PP(16'h1998,4);
TASK_PP(16'h1999,4);
TASK_PP(16'h199A,4);
TASK_PP(16'h199B,4);
TASK_PP(16'h199C,4);
TASK_PP(16'h199D,4);
TASK_PP(16'h199E,4);
TASK_PP(16'h199F,4);
TASK_PP(16'h19A0,4);
TASK_PP(16'h19A1,4);
TASK_PP(16'h19A2,4);
TASK_PP(16'h19A3,4);
TASK_PP(16'h19A4,4);
TASK_PP(16'h19A5,4);
TASK_PP(16'h19A6,4);
TASK_PP(16'h19A7,4);
TASK_PP(16'h19A8,4);
TASK_PP(16'h19A9,4);
TASK_PP(16'h19AA,4);
TASK_PP(16'h19AB,4);
TASK_PP(16'h19AC,4);
TASK_PP(16'h19AD,4);
TASK_PP(16'h19AE,4);
TASK_PP(16'h19AF,4);
TASK_PP(16'h19B0,4);
TASK_PP(16'h19B1,4);
TASK_PP(16'h19B2,4);
TASK_PP(16'h19B3,4);
TASK_PP(16'h19B4,4);
TASK_PP(16'h19B5,4);
TASK_PP(16'h19B6,4);
TASK_PP(16'h19B7,4);
TASK_PP(16'h19B8,4);
TASK_PP(16'h19B9,4);
TASK_PP(16'h19BA,4);
TASK_PP(16'h19BB,4);
TASK_PP(16'h19BC,4);
TASK_PP(16'h19BD,4);
TASK_PP(16'h19BE,4);
TASK_PP(16'h19BF,4);
TASK_PP(16'h19C0,4);
TASK_PP(16'h19C1,4);
TASK_PP(16'h19C2,4);
TASK_PP(16'h19C3,4);
TASK_PP(16'h19C4,4);
TASK_PP(16'h19C5,4);
TASK_PP(16'h19C6,4);
TASK_PP(16'h19C7,4);
TASK_PP(16'h19C8,4);
TASK_PP(16'h19C9,4);
TASK_PP(16'h19CA,4);
TASK_PP(16'h19CB,4);
TASK_PP(16'h19CC,4);
TASK_PP(16'h19CD,4);
TASK_PP(16'h19CE,4);
TASK_PP(16'h19CF,4);
TASK_PP(16'h19D0,4);
TASK_PP(16'h19D1,4);
TASK_PP(16'h19D2,4);
TASK_PP(16'h19D3,4);
TASK_PP(16'h19D4,4);
TASK_PP(16'h19D5,4);
TASK_PP(16'h19D6,4);
TASK_PP(16'h19D7,4);
TASK_PP(16'h19D8,4);
TASK_PP(16'h19D9,4);
TASK_PP(16'h19DA,4);
TASK_PP(16'h19DB,4);
TASK_PP(16'h19DC,4);
TASK_PP(16'h19DD,4);
TASK_PP(16'h19DE,4);
TASK_PP(16'h19DF,4);
TASK_PP(16'h19E0,4);
TASK_PP(16'h19E1,4);
TASK_PP(16'h19E2,4);
TASK_PP(16'h19E3,4);
TASK_PP(16'h19E4,4);
TASK_PP(16'h19E5,4);
TASK_PP(16'h19E6,4);
TASK_PP(16'h19E7,4);
TASK_PP(16'h19E8,4);
TASK_PP(16'h19E9,4);
TASK_PP(16'h19EA,4);
TASK_PP(16'h19EB,4);
TASK_PP(16'h19EC,4);
TASK_PP(16'h19ED,4);
TASK_PP(16'h19EE,4);
TASK_PP(16'h19EF,4);
TASK_PP(16'h19F0,4);
TASK_PP(16'h19F1,4);
TASK_PP(16'h19F2,4);
TASK_PP(16'h19F3,4);
TASK_PP(16'h19F4,4);
TASK_PP(16'h19F5,4);
TASK_PP(16'h19F6,4);
TASK_PP(16'h19F7,4);
TASK_PP(16'h19F8,4);
TASK_PP(16'h19F9,4);
TASK_PP(16'h19FA,4);
TASK_PP(16'h19FB,4);
TASK_PP(16'h19FC,4);
TASK_PP(16'h19FD,4);
TASK_PP(16'h19FE,4);
TASK_PP(16'h19FF,4);
TASK_PP(16'h1A00,4);
TASK_PP(16'h1A01,4);
TASK_PP(16'h1A02,4);
TASK_PP(16'h1A03,4);
TASK_PP(16'h1A04,4);
TASK_PP(16'h1A05,4);
TASK_PP(16'h1A06,4);
TASK_PP(16'h1A07,4);
TASK_PP(16'h1A08,4);
TASK_PP(16'h1A09,4);
TASK_PP(16'h1A0A,4);
TASK_PP(16'h1A0B,4);
TASK_PP(16'h1A0C,4);
TASK_PP(16'h1A0D,4);
TASK_PP(16'h1A0E,4);
TASK_PP(16'h1A0F,4);
TASK_PP(16'h1A10,4);
TASK_PP(16'h1A11,4);
TASK_PP(16'h1A12,4);
TASK_PP(16'h1A13,4);
TASK_PP(16'h1A14,4);
TASK_PP(16'h1A15,4);
TASK_PP(16'h1A16,4);
TASK_PP(16'h1A17,4);
TASK_PP(16'h1A18,4);
TASK_PP(16'h1A19,4);
TASK_PP(16'h1A1A,4);
TASK_PP(16'h1A1B,4);
TASK_PP(16'h1A1C,4);
TASK_PP(16'h1A1D,4);
TASK_PP(16'h1A1E,4);
TASK_PP(16'h1A1F,4);
TASK_PP(16'h1A20,4);
TASK_PP(16'h1A21,4);
TASK_PP(16'h1A22,4);
TASK_PP(16'h1A23,4);
TASK_PP(16'h1A24,4);
TASK_PP(16'h1A25,4);
TASK_PP(16'h1A26,4);
TASK_PP(16'h1A27,4);
TASK_PP(16'h1A28,4);
TASK_PP(16'h1A29,4);
TASK_PP(16'h1A2A,4);
TASK_PP(16'h1A2B,4);
TASK_PP(16'h1A2C,4);
TASK_PP(16'h1A2D,4);
TASK_PP(16'h1A2E,4);
TASK_PP(16'h1A2F,4);
TASK_PP(16'h1A30,4);
TASK_PP(16'h1A31,4);
TASK_PP(16'h1A32,4);
TASK_PP(16'h1A33,4);
TASK_PP(16'h1A34,4);
TASK_PP(16'h1A35,4);
TASK_PP(16'h1A36,4);
TASK_PP(16'h1A37,4);
TASK_PP(16'h1A38,4);
TASK_PP(16'h1A39,4);
TASK_PP(16'h1A3A,4);
TASK_PP(16'h1A3B,4);
TASK_PP(16'h1A3C,4);
TASK_PP(16'h1A3D,4);
TASK_PP(16'h1A3E,4);
TASK_PP(16'h1A3F,4);
TASK_PP(16'h1A40,4);
TASK_PP(16'h1A41,4);
TASK_PP(16'h1A42,4);
TASK_PP(16'h1A43,4);
TASK_PP(16'h1A44,4);
TASK_PP(16'h1A45,4);
TASK_PP(16'h1A46,4);
TASK_PP(16'h1A47,4);
TASK_PP(16'h1A48,4);
TASK_PP(16'h1A49,4);
TASK_PP(16'h1A4A,4);
TASK_PP(16'h1A4B,4);
TASK_PP(16'h1A4C,4);
TASK_PP(16'h1A4D,4);
TASK_PP(16'h1A4E,4);
TASK_PP(16'h1A4F,4);
TASK_PP(16'h1A50,4);
TASK_PP(16'h1A51,4);
TASK_PP(16'h1A52,4);
TASK_PP(16'h1A53,4);
TASK_PP(16'h1A54,4);
TASK_PP(16'h1A55,4);
TASK_PP(16'h1A56,4);
TASK_PP(16'h1A57,4);
TASK_PP(16'h1A58,4);
TASK_PP(16'h1A59,4);
TASK_PP(16'h1A5A,4);
TASK_PP(16'h1A5B,4);
TASK_PP(16'h1A5C,4);
TASK_PP(16'h1A5D,4);
TASK_PP(16'h1A5E,4);
TASK_PP(16'h1A5F,4);
TASK_PP(16'h1A60,4);
TASK_PP(16'h1A61,4);
TASK_PP(16'h1A62,4);
TASK_PP(16'h1A63,4);
TASK_PP(16'h1A64,4);
TASK_PP(16'h1A65,4);
TASK_PP(16'h1A66,4);
TASK_PP(16'h1A67,4);
TASK_PP(16'h1A68,4);
TASK_PP(16'h1A69,4);
TASK_PP(16'h1A6A,4);
TASK_PP(16'h1A6B,4);
TASK_PP(16'h1A6C,4);
TASK_PP(16'h1A6D,4);
TASK_PP(16'h1A6E,4);
TASK_PP(16'h1A6F,4);
TASK_PP(16'h1A70,4);
TASK_PP(16'h1A71,4);
TASK_PP(16'h1A72,4);
TASK_PP(16'h1A73,4);
TASK_PP(16'h1A74,4);
TASK_PP(16'h1A75,4);
TASK_PP(16'h1A76,4);
TASK_PP(16'h1A77,4);
TASK_PP(16'h1A78,4);
TASK_PP(16'h1A79,4);
TASK_PP(16'h1A7A,4);
TASK_PP(16'h1A7B,4);
TASK_PP(16'h1A7C,4);
TASK_PP(16'h1A7D,4);
TASK_PP(16'h1A7E,4);
TASK_PP(16'h1A7F,4);
TASK_PP(16'h1A80,4);
TASK_PP(16'h1A81,4);
TASK_PP(16'h1A82,4);
TASK_PP(16'h1A83,4);
TASK_PP(16'h1A84,4);
TASK_PP(16'h1A85,4);
TASK_PP(16'h1A86,4);
TASK_PP(16'h1A87,4);
TASK_PP(16'h1A88,4);
TASK_PP(16'h1A89,4);
TASK_PP(16'h1A8A,4);
TASK_PP(16'h1A8B,4);
TASK_PP(16'h1A8C,4);
TASK_PP(16'h1A8D,4);
TASK_PP(16'h1A8E,4);
TASK_PP(16'h1A8F,4);
TASK_PP(16'h1A90,4);
TASK_PP(16'h1A91,4);
TASK_PP(16'h1A92,4);
TASK_PP(16'h1A93,4);
TASK_PP(16'h1A94,4);
TASK_PP(16'h1A95,4);
TASK_PP(16'h1A96,4);
TASK_PP(16'h1A97,4);
TASK_PP(16'h1A98,4);
TASK_PP(16'h1A99,4);
TASK_PP(16'h1A9A,4);
TASK_PP(16'h1A9B,4);
TASK_PP(16'h1A9C,4);
TASK_PP(16'h1A9D,4);
TASK_PP(16'h1A9E,4);
TASK_PP(16'h1A9F,4);
TASK_PP(16'h1AA0,4);
TASK_PP(16'h1AA1,4);
TASK_PP(16'h1AA2,4);
TASK_PP(16'h1AA3,4);
TASK_PP(16'h1AA4,4);
TASK_PP(16'h1AA5,4);
TASK_PP(16'h1AA6,4);
TASK_PP(16'h1AA7,4);
TASK_PP(16'h1AA8,4);
TASK_PP(16'h1AA9,4);
TASK_PP(16'h1AAA,4);
TASK_PP(16'h1AAB,4);
TASK_PP(16'h1AAC,4);
TASK_PP(16'h1AAD,4);
TASK_PP(16'h1AAE,4);
TASK_PP(16'h1AAF,4);
TASK_PP(16'h1AB0,4);
TASK_PP(16'h1AB1,4);
TASK_PP(16'h1AB2,4);
TASK_PP(16'h1AB3,4);
TASK_PP(16'h1AB4,4);
TASK_PP(16'h1AB5,4);
TASK_PP(16'h1AB6,4);
TASK_PP(16'h1AB7,4);
TASK_PP(16'h1AB8,4);
TASK_PP(16'h1AB9,4);
TASK_PP(16'h1ABA,4);
TASK_PP(16'h1ABB,4);
TASK_PP(16'h1ABC,4);
TASK_PP(16'h1ABD,4);
TASK_PP(16'h1ABE,4);
TASK_PP(16'h1ABF,4);
TASK_PP(16'h1AC0,4);
TASK_PP(16'h1AC1,4);
TASK_PP(16'h1AC2,4);
TASK_PP(16'h1AC3,4);
TASK_PP(16'h1AC4,4);
TASK_PP(16'h1AC5,4);
TASK_PP(16'h1AC6,4);
TASK_PP(16'h1AC7,4);
TASK_PP(16'h1AC8,4);
TASK_PP(16'h1AC9,4);
TASK_PP(16'h1ACA,4);
TASK_PP(16'h1ACB,4);
TASK_PP(16'h1ACC,4);
TASK_PP(16'h1ACD,4);
TASK_PP(16'h1ACE,4);
TASK_PP(16'h1ACF,4);
TASK_PP(16'h1AD0,4);
TASK_PP(16'h1AD1,4);
TASK_PP(16'h1AD2,4);
TASK_PP(16'h1AD3,4);
TASK_PP(16'h1AD4,4);
TASK_PP(16'h1AD5,4);
TASK_PP(16'h1AD6,4);
TASK_PP(16'h1AD7,4);
TASK_PP(16'h1AD8,4);
TASK_PP(16'h1AD9,4);
TASK_PP(16'h1ADA,4);
TASK_PP(16'h1ADB,4);
TASK_PP(16'h1ADC,4);
TASK_PP(16'h1ADD,4);
TASK_PP(16'h1ADE,4);
TASK_PP(16'h1ADF,4);
TASK_PP(16'h1AE0,4);
TASK_PP(16'h1AE1,4);
TASK_PP(16'h1AE2,4);
TASK_PP(16'h1AE3,4);
TASK_PP(16'h1AE4,4);
TASK_PP(16'h1AE5,4);
TASK_PP(16'h1AE6,4);
TASK_PP(16'h1AE7,4);
TASK_PP(16'h1AE8,4);
TASK_PP(16'h1AE9,4);
TASK_PP(16'h1AEA,4);
TASK_PP(16'h1AEB,4);
TASK_PP(16'h1AEC,4);
TASK_PP(16'h1AED,4);
TASK_PP(16'h1AEE,4);
TASK_PP(16'h1AEF,4);
TASK_PP(16'h1AF0,4);
TASK_PP(16'h1AF1,4);
TASK_PP(16'h1AF2,4);
TASK_PP(16'h1AF3,4);
TASK_PP(16'h1AF4,4);
TASK_PP(16'h1AF5,4);
TASK_PP(16'h1AF6,4);
TASK_PP(16'h1AF7,4);
TASK_PP(16'h1AF8,4);
TASK_PP(16'h1AF9,4);
TASK_PP(16'h1AFA,4);
TASK_PP(16'h1AFB,4);
TASK_PP(16'h1AFC,4);
TASK_PP(16'h1AFD,4);
TASK_PP(16'h1AFE,4);
TASK_PP(16'h1AFF,4);
TASK_PP(16'h1B00,4);
TASK_PP(16'h1B01,4);
TASK_PP(16'h1B02,4);
TASK_PP(16'h1B03,4);
TASK_PP(16'h1B04,4);
TASK_PP(16'h1B05,4);
TASK_PP(16'h1B06,4);
TASK_PP(16'h1B07,4);
TASK_PP(16'h1B08,4);
TASK_PP(16'h1B09,4);
TASK_PP(16'h1B0A,4);
TASK_PP(16'h1B0B,4);
TASK_PP(16'h1B0C,4);
TASK_PP(16'h1B0D,4);
TASK_PP(16'h1B0E,4);
TASK_PP(16'h1B0F,4);
TASK_PP(16'h1B10,4);
TASK_PP(16'h1B11,4);
TASK_PP(16'h1B12,4);
TASK_PP(16'h1B13,4);
TASK_PP(16'h1B14,4);
TASK_PP(16'h1B15,4);
TASK_PP(16'h1B16,4);
TASK_PP(16'h1B17,4);
TASK_PP(16'h1B18,4);
TASK_PP(16'h1B19,4);
TASK_PP(16'h1B1A,4);
TASK_PP(16'h1B1B,4);
TASK_PP(16'h1B1C,4);
TASK_PP(16'h1B1D,4);
TASK_PP(16'h1B1E,4);
TASK_PP(16'h1B1F,4);
TASK_PP(16'h1B20,4);
TASK_PP(16'h1B21,4);
TASK_PP(16'h1B22,4);
TASK_PP(16'h1B23,4);
TASK_PP(16'h1B24,4);
TASK_PP(16'h1B25,4);
TASK_PP(16'h1B26,4);
TASK_PP(16'h1B27,4);
TASK_PP(16'h1B28,4);
TASK_PP(16'h1B29,4);
TASK_PP(16'h1B2A,4);
TASK_PP(16'h1B2B,4);
TASK_PP(16'h1B2C,4);
TASK_PP(16'h1B2D,4);
TASK_PP(16'h1B2E,4);
TASK_PP(16'h1B2F,4);
TASK_PP(16'h1B30,4);
TASK_PP(16'h1B31,4);
TASK_PP(16'h1B32,4);
TASK_PP(16'h1B33,4);
TASK_PP(16'h1B34,4);
TASK_PP(16'h1B35,4);
TASK_PP(16'h1B36,4);
TASK_PP(16'h1B37,4);
TASK_PP(16'h1B38,4);
TASK_PP(16'h1B39,4);
TASK_PP(16'h1B3A,4);
TASK_PP(16'h1B3B,4);
TASK_PP(16'h1B3C,4);
TASK_PP(16'h1B3D,4);
TASK_PP(16'h1B3E,4);
TASK_PP(16'h1B3F,4);
TASK_PP(16'h1B40,4);
TASK_PP(16'h1B41,4);
TASK_PP(16'h1B42,4);
TASK_PP(16'h1B43,4);
TASK_PP(16'h1B44,4);
TASK_PP(16'h1B45,4);
TASK_PP(16'h1B46,4);
TASK_PP(16'h1B47,4);
TASK_PP(16'h1B48,4);
TASK_PP(16'h1B49,4);
TASK_PP(16'h1B4A,4);
TASK_PP(16'h1B4B,4);
TASK_PP(16'h1B4C,4);
TASK_PP(16'h1B4D,4);
TASK_PP(16'h1B4E,4);
TASK_PP(16'h1B4F,4);
TASK_PP(16'h1B50,4);
TASK_PP(16'h1B51,4);
TASK_PP(16'h1B52,4);
TASK_PP(16'h1B53,4);
TASK_PP(16'h1B54,4);
TASK_PP(16'h1B55,4);
TASK_PP(16'h1B56,4);
TASK_PP(16'h1B57,4);
TASK_PP(16'h1B58,4);
TASK_PP(16'h1B59,4);
TASK_PP(16'h1B5A,4);
TASK_PP(16'h1B5B,4);
TASK_PP(16'h1B5C,4);
TASK_PP(16'h1B5D,4);
TASK_PP(16'h1B5E,4);
TASK_PP(16'h1B5F,4);
TASK_PP(16'h1B60,4);
TASK_PP(16'h1B61,4);
TASK_PP(16'h1B62,4);
TASK_PP(16'h1B63,4);
TASK_PP(16'h1B64,4);
TASK_PP(16'h1B65,4);
TASK_PP(16'h1B66,4);
TASK_PP(16'h1B67,4);
TASK_PP(16'h1B68,4);
TASK_PP(16'h1B69,4);
TASK_PP(16'h1B6A,4);
TASK_PP(16'h1B6B,4);
TASK_PP(16'h1B6C,4);
TASK_PP(16'h1B6D,4);
TASK_PP(16'h1B6E,4);
TASK_PP(16'h1B6F,4);
TASK_PP(16'h1B70,4);
TASK_PP(16'h1B71,4);
TASK_PP(16'h1B72,4);
TASK_PP(16'h1B73,4);
TASK_PP(16'h1B74,4);
TASK_PP(16'h1B75,4);
TASK_PP(16'h1B76,4);
TASK_PP(16'h1B77,4);
TASK_PP(16'h1B78,4);
TASK_PP(16'h1B79,4);
TASK_PP(16'h1B7A,4);
TASK_PP(16'h1B7B,4);
TASK_PP(16'h1B7C,4);
TASK_PP(16'h1B7D,4);
TASK_PP(16'h1B7E,4);
TASK_PP(16'h1B7F,4);
TASK_PP(16'h1B80,4);
TASK_PP(16'h1B81,4);
TASK_PP(16'h1B82,4);
TASK_PP(16'h1B83,4);
TASK_PP(16'h1B84,4);
TASK_PP(16'h1B85,4);
TASK_PP(16'h1B86,4);
TASK_PP(16'h1B87,4);
TASK_PP(16'h1B88,4);
TASK_PP(16'h1B89,4);
TASK_PP(16'h1B8A,4);
TASK_PP(16'h1B8B,4);
TASK_PP(16'h1B8C,4);
TASK_PP(16'h1B8D,4);
TASK_PP(16'h1B8E,4);
TASK_PP(16'h1B8F,4);
TASK_PP(16'h1B90,4);
TASK_PP(16'h1B91,4);
TASK_PP(16'h1B92,4);
TASK_PP(16'h1B93,4);
TASK_PP(16'h1B94,4);
TASK_PP(16'h1B95,4);
TASK_PP(16'h1B96,4);
TASK_PP(16'h1B97,4);
TASK_PP(16'h1B98,4);
TASK_PP(16'h1B99,4);
TASK_PP(16'h1B9A,4);
TASK_PP(16'h1B9B,4);
TASK_PP(16'h1B9C,4);
TASK_PP(16'h1B9D,4);
TASK_PP(16'h1B9E,4);
TASK_PP(16'h1B9F,4);
TASK_PP(16'h1BA0,4);
TASK_PP(16'h1BA1,4);
TASK_PP(16'h1BA2,4);
TASK_PP(16'h1BA3,4);
TASK_PP(16'h1BA4,4);
TASK_PP(16'h1BA5,4);
TASK_PP(16'h1BA6,4);
TASK_PP(16'h1BA7,4);
TASK_PP(16'h1BA8,4);
TASK_PP(16'h1BA9,4);
TASK_PP(16'h1BAA,4);
TASK_PP(16'h1BAB,4);
TASK_PP(16'h1BAC,4);
TASK_PP(16'h1BAD,4);
TASK_PP(16'h1BAE,4);
TASK_PP(16'h1BAF,4);
TASK_PP(16'h1BB0,4);
TASK_PP(16'h1BB1,4);
TASK_PP(16'h1BB2,4);
TASK_PP(16'h1BB3,4);
TASK_PP(16'h1BB4,4);
TASK_PP(16'h1BB5,4);
TASK_PP(16'h1BB6,4);
TASK_PP(16'h1BB7,4);
TASK_PP(16'h1BB8,4);
TASK_PP(16'h1BB9,4);
TASK_PP(16'h1BBA,4);
TASK_PP(16'h1BBB,4);
TASK_PP(16'h1BBC,4);
TASK_PP(16'h1BBD,4);
TASK_PP(16'h1BBE,4);
TASK_PP(16'h1BBF,4);
TASK_PP(16'h1BC0,4);
TASK_PP(16'h1BC1,4);
TASK_PP(16'h1BC2,4);
TASK_PP(16'h1BC3,4);
TASK_PP(16'h1BC4,4);
TASK_PP(16'h1BC5,4);
TASK_PP(16'h1BC6,4);
TASK_PP(16'h1BC7,4);
TASK_PP(16'h1BC8,4);
TASK_PP(16'h1BC9,4);
TASK_PP(16'h1BCA,4);
TASK_PP(16'h1BCB,4);
TASK_PP(16'h1BCC,4);
TASK_PP(16'h1BCD,4);
TASK_PP(16'h1BCE,4);
TASK_PP(16'h1BCF,4);
TASK_PP(16'h1BD0,4);
TASK_PP(16'h1BD1,4);
TASK_PP(16'h1BD2,4);
TASK_PP(16'h1BD3,4);
TASK_PP(16'h1BD4,4);
TASK_PP(16'h1BD5,4);
TASK_PP(16'h1BD6,4);
TASK_PP(16'h1BD7,4);
TASK_PP(16'h1BD8,4);
TASK_PP(16'h1BD9,4);
TASK_PP(16'h1BDA,4);
TASK_PP(16'h1BDB,4);
TASK_PP(16'h1BDC,4);
TASK_PP(16'h1BDD,4);
TASK_PP(16'h1BDE,4);
TASK_PP(16'h1BDF,4);
TASK_PP(16'h1BE0,4);
TASK_PP(16'h1BE1,4);
TASK_PP(16'h1BE2,4);
TASK_PP(16'h1BE3,4);
TASK_PP(16'h1BE4,4);
TASK_PP(16'h1BE5,4);
TASK_PP(16'h1BE6,4);
TASK_PP(16'h1BE7,4);
TASK_PP(16'h1BE8,4);
TASK_PP(16'h1BE9,4);
TASK_PP(16'h1BEA,4);
TASK_PP(16'h1BEB,4);
TASK_PP(16'h1BEC,4);
TASK_PP(16'h1BED,4);
TASK_PP(16'h1BEE,4);
TASK_PP(16'h1BEF,4);
TASK_PP(16'h1BF0,4);
TASK_PP(16'h1BF1,4);
TASK_PP(16'h1BF2,4);
TASK_PP(16'h1BF3,4);
TASK_PP(16'h1BF4,4);
TASK_PP(16'h1BF5,4);
TASK_PP(16'h1BF6,4);
TASK_PP(16'h1BF7,4);
TASK_PP(16'h1BF8,4);
TASK_PP(16'h1BF9,4);
TASK_PP(16'h1BFA,4);
TASK_PP(16'h1BFB,4);
TASK_PP(16'h1BFC,4);
TASK_PP(16'h1BFD,4);
TASK_PP(16'h1BFE,4);
TASK_PP(16'h1BFF,4);
TASK_PP(16'h1C00,4);
TASK_PP(16'h1C01,4);
TASK_PP(16'h1C02,4);
TASK_PP(16'h1C03,4);
TASK_PP(16'h1C04,4);
TASK_PP(16'h1C05,4);
TASK_PP(16'h1C06,4);
TASK_PP(16'h1C07,4);
TASK_PP(16'h1C08,4);
TASK_PP(16'h1C09,4);
TASK_PP(16'h1C0A,4);
TASK_PP(16'h1C0B,4);
TASK_PP(16'h1C0C,4);
TASK_PP(16'h1C0D,4);
TASK_PP(16'h1C0E,4);
TASK_PP(16'h1C0F,4);
TASK_PP(16'h1C10,4);
TASK_PP(16'h1C11,4);
TASK_PP(16'h1C12,4);
TASK_PP(16'h1C13,4);
TASK_PP(16'h1C14,4);
TASK_PP(16'h1C15,4);
TASK_PP(16'h1C16,4);
TASK_PP(16'h1C17,4);
TASK_PP(16'h1C18,4);
TASK_PP(16'h1C19,4);
TASK_PP(16'h1C1A,4);
TASK_PP(16'h1C1B,4);
TASK_PP(16'h1C1C,4);
TASK_PP(16'h1C1D,4);
TASK_PP(16'h1C1E,4);
TASK_PP(16'h1C1F,4);
TASK_PP(16'h1C20,4);
TASK_PP(16'h1C21,4);
TASK_PP(16'h1C22,4);
TASK_PP(16'h1C23,4);
TASK_PP(16'h1C24,4);
TASK_PP(16'h1C25,4);
TASK_PP(16'h1C26,4);
TASK_PP(16'h1C27,4);
TASK_PP(16'h1C28,4);
TASK_PP(16'h1C29,4);
TASK_PP(16'h1C2A,4);
TASK_PP(16'h1C2B,4);
TASK_PP(16'h1C2C,4);
TASK_PP(16'h1C2D,4);
TASK_PP(16'h1C2E,4);
TASK_PP(16'h1C2F,4);
TASK_PP(16'h1C30,4);
TASK_PP(16'h1C31,4);
TASK_PP(16'h1C32,4);
TASK_PP(16'h1C33,4);
TASK_PP(16'h1C34,4);
TASK_PP(16'h1C35,4);
TASK_PP(16'h1C36,4);
TASK_PP(16'h1C37,4);
TASK_PP(16'h1C38,4);
TASK_PP(16'h1C39,4);
TASK_PP(16'h1C3A,4);
TASK_PP(16'h1C3B,4);
TASK_PP(16'h1C3C,4);
TASK_PP(16'h1C3D,4);
TASK_PP(16'h1C3E,4);
TASK_PP(16'h1C3F,4);
TASK_PP(16'h1C40,4);
TASK_PP(16'h1C41,4);
TASK_PP(16'h1C42,4);
TASK_PP(16'h1C43,4);
TASK_PP(16'h1C44,4);
TASK_PP(16'h1C45,4);
TASK_PP(16'h1C46,4);
TASK_PP(16'h1C47,4);
TASK_PP(16'h1C48,4);
TASK_PP(16'h1C49,4);
TASK_PP(16'h1C4A,4);
TASK_PP(16'h1C4B,4);
TASK_PP(16'h1C4C,4);
TASK_PP(16'h1C4D,4);
TASK_PP(16'h1C4E,4);
TASK_PP(16'h1C4F,4);
TASK_PP(16'h1C50,4);
TASK_PP(16'h1C51,4);
TASK_PP(16'h1C52,4);
TASK_PP(16'h1C53,4);
TASK_PP(16'h1C54,4);
TASK_PP(16'h1C55,4);
TASK_PP(16'h1C56,4);
TASK_PP(16'h1C57,4);
TASK_PP(16'h1C58,4);
TASK_PP(16'h1C59,4);
TASK_PP(16'h1C5A,4);
TASK_PP(16'h1C5B,4);
TASK_PP(16'h1C5C,4);
TASK_PP(16'h1C5D,4);
TASK_PP(16'h1C5E,4);
TASK_PP(16'h1C5F,4);
TASK_PP(16'h1C60,4);
TASK_PP(16'h1C61,4);
TASK_PP(16'h1C62,4);
TASK_PP(16'h1C63,4);
TASK_PP(16'h1C64,4);
TASK_PP(16'h1C65,4);
TASK_PP(16'h1C66,4);
TASK_PP(16'h1C67,4);
TASK_PP(16'h1C68,4);
TASK_PP(16'h1C69,4);
TASK_PP(16'h1C6A,4);
TASK_PP(16'h1C6B,4);
TASK_PP(16'h1C6C,4);
TASK_PP(16'h1C6D,4);
TASK_PP(16'h1C6E,4);
TASK_PP(16'h1C6F,4);
TASK_PP(16'h1C70,4);
TASK_PP(16'h1C71,4);
TASK_PP(16'h1C72,4);
TASK_PP(16'h1C73,4);
TASK_PP(16'h1C74,4);
TASK_PP(16'h1C75,4);
TASK_PP(16'h1C76,4);
TASK_PP(16'h1C77,4);
TASK_PP(16'h1C78,4);
TASK_PP(16'h1C79,4);
TASK_PP(16'h1C7A,4);
TASK_PP(16'h1C7B,4);
TASK_PP(16'h1C7C,4);
TASK_PP(16'h1C7D,4);
TASK_PP(16'h1C7E,4);
TASK_PP(16'h1C7F,4);
TASK_PP(16'h1C80,4);
TASK_PP(16'h1C81,4);
TASK_PP(16'h1C82,4);
TASK_PP(16'h1C83,4);
TASK_PP(16'h1C84,4);
TASK_PP(16'h1C85,4);
TASK_PP(16'h1C86,4);
TASK_PP(16'h1C87,4);
TASK_PP(16'h1C88,4);
TASK_PP(16'h1C89,4);
TASK_PP(16'h1C8A,4);
TASK_PP(16'h1C8B,4);
TASK_PP(16'h1C8C,4);
TASK_PP(16'h1C8D,4);
TASK_PP(16'h1C8E,4);
TASK_PP(16'h1C8F,4);
TASK_PP(16'h1C90,4);
TASK_PP(16'h1C91,4);
TASK_PP(16'h1C92,4);
TASK_PP(16'h1C93,4);
TASK_PP(16'h1C94,4);
TASK_PP(16'h1C95,4);
TASK_PP(16'h1C96,4);
TASK_PP(16'h1C97,4);
TASK_PP(16'h1C98,4);
TASK_PP(16'h1C99,4);
TASK_PP(16'h1C9A,4);
TASK_PP(16'h1C9B,4);
TASK_PP(16'h1C9C,4);
TASK_PP(16'h1C9D,4);
TASK_PP(16'h1C9E,4);
TASK_PP(16'h1C9F,4);
TASK_PP(16'h1CA0,4);
TASK_PP(16'h1CA1,4);
TASK_PP(16'h1CA2,4);
TASK_PP(16'h1CA3,4);
TASK_PP(16'h1CA4,4);
TASK_PP(16'h1CA5,4);
TASK_PP(16'h1CA6,4);
TASK_PP(16'h1CA7,4);
TASK_PP(16'h1CA8,4);
TASK_PP(16'h1CA9,4);
TASK_PP(16'h1CAA,4);
TASK_PP(16'h1CAB,4);
TASK_PP(16'h1CAC,4);
TASK_PP(16'h1CAD,4);
TASK_PP(16'h1CAE,4);
TASK_PP(16'h1CAF,4);
TASK_PP(16'h1CB0,4);
TASK_PP(16'h1CB1,4);
TASK_PP(16'h1CB2,4);
TASK_PP(16'h1CB3,4);
TASK_PP(16'h1CB4,4);
TASK_PP(16'h1CB5,4);
TASK_PP(16'h1CB6,4);
TASK_PP(16'h1CB7,4);
TASK_PP(16'h1CB8,4);
TASK_PP(16'h1CB9,4);
TASK_PP(16'h1CBA,4);
TASK_PP(16'h1CBB,4);
TASK_PP(16'h1CBC,4);
TASK_PP(16'h1CBD,4);
TASK_PP(16'h1CBE,4);
TASK_PP(16'h1CBF,4);
TASK_PP(16'h1CC0,4);
TASK_PP(16'h1CC1,4);
TASK_PP(16'h1CC2,4);
TASK_PP(16'h1CC3,4);
TASK_PP(16'h1CC4,4);
TASK_PP(16'h1CC5,4);
TASK_PP(16'h1CC6,4);
TASK_PP(16'h1CC7,4);
TASK_PP(16'h1CC8,4);
TASK_PP(16'h1CC9,4);
TASK_PP(16'h1CCA,4);
TASK_PP(16'h1CCB,4);
TASK_PP(16'h1CCC,4);
TASK_PP(16'h1CCD,4);
TASK_PP(16'h1CCE,4);
TASK_PP(16'h1CCF,4);
TASK_PP(16'h1CD0,4);
TASK_PP(16'h1CD1,4);
TASK_PP(16'h1CD2,4);
TASK_PP(16'h1CD3,4);
TASK_PP(16'h1CD4,4);
TASK_PP(16'h1CD5,4);
TASK_PP(16'h1CD6,4);
TASK_PP(16'h1CD7,4);
TASK_PP(16'h1CD8,4);
TASK_PP(16'h1CD9,4);
TASK_PP(16'h1CDA,4);
TASK_PP(16'h1CDB,4);
TASK_PP(16'h1CDC,4);
TASK_PP(16'h1CDD,4);
TASK_PP(16'h1CDE,4);
TASK_PP(16'h1CDF,4);
TASK_PP(16'h1CE0,4);
TASK_PP(16'h1CE1,4);
TASK_PP(16'h1CE2,4);
TASK_PP(16'h1CE3,4);
TASK_PP(16'h1CE4,4);
TASK_PP(16'h1CE5,4);
TASK_PP(16'h1CE6,4);
TASK_PP(16'h1CE7,4);
TASK_PP(16'h1CE8,4);
TASK_PP(16'h1CE9,4);
TASK_PP(16'h1CEA,4);
TASK_PP(16'h1CEB,4);
TASK_PP(16'h1CEC,4);
TASK_PP(16'h1CED,4);
TASK_PP(16'h1CEE,4);
TASK_PP(16'h1CEF,4);
TASK_PP(16'h1CF0,4);
TASK_PP(16'h1CF1,4);
TASK_PP(16'h1CF2,4);
TASK_PP(16'h1CF3,4);
TASK_PP(16'h1CF4,4);
TASK_PP(16'h1CF5,4);
TASK_PP(16'h1CF6,4);
TASK_PP(16'h1CF7,4);
TASK_PP(16'h1CF8,4);
TASK_PP(16'h1CF9,4);
TASK_PP(16'h1CFA,4);
TASK_PP(16'h1CFB,4);
TASK_PP(16'h1CFC,4);
TASK_PP(16'h1CFD,4);
TASK_PP(16'h1CFE,4);
TASK_PP(16'h1CFF,4);
TASK_PP(16'h1D00,4);
TASK_PP(16'h1D01,4);
TASK_PP(16'h1D02,4);
TASK_PP(16'h1D03,4);
TASK_PP(16'h1D04,4);
TASK_PP(16'h1D05,4);
TASK_PP(16'h1D06,4);
TASK_PP(16'h1D07,4);
TASK_PP(16'h1D08,4);
TASK_PP(16'h1D09,4);
TASK_PP(16'h1D0A,4);
TASK_PP(16'h1D0B,4);
TASK_PP(16'h1D0C,4);
TASK_PP(16'h1D0D,4);
TASK_PP(16'h1D0E,4);
TASK_PP(16'h1D0F,4);
TASK_PP(16'h1D10,4);
TASK_PP(16'h1D11,4);
TASK_PP(16'h1D12,4);
TASK_PP(16'h1D13,4);
TASK_PP(16'h1D14,4);
TASK_PP(16'h1D15,4);
TASK_PP(16'h1D16,4);
TASK_PP(16'h1D17,4);
TASK_PP(16'h1D18,4);
TASK_PP(16'h1D19,4);
TASK_PP(16'h1D1A,4);
TASK_PP(16'h1D1B,4);
TASK_PP(16'h1D1C,4);
TASK_PP(16'h1D1D,4);
TASK_PP(16'h1D1E,4);
TASK_PP(16'h1D1F,4);
TASK_PP(16'h1D20,4);
TASK_PP(16'h1D21,4);
TASK_PP(16'h1D22,4);
TASK_PP(16'h1D23,4);
TASK_PP(16'h1D24,4);
TASK_PP(16'h1D25,4);
TASK_PP(16'h1D26,4);
TASK_PP(16'h1D27,4);
TASK_PP(16'h1D28,4);
TASK_PP(16'h1D29,4);
TASK_PP(16'h1D2A,4);
TASK_PP(16'h1D2B,4);
TASK_PP(16'h1D2C,4);
TASK_PP(16'h1D2D,4);
TASK_PP(16'h1D2E,4);
TASK_PP(16'h1D2F,4);
TASK_PP(16'h1D30,4);
TASK_PP(16'h1D31,4);
TASK_PP(16'h1D32,4);
TASK_PP(16'h1D33,4);
TASK_PP(16'h1D34,4);
TASK_PP(16'h1D35,4);
TASK_PP(16'h1D36,4);
TASK_PP(16'h1D37,4);
TASK_PP(16'h1D38,4);
TASK_PP(16'h1D39,4);
TASK_PP(16'h1D3A,4);
TASK_PP(16'h1D3B,4);
TASK_PP(16'h1D3C,4);
TASK_PP(16'h1D3D,4);
TASK_PP(16'h1D3E,4);
TASK_PP(16'h1D3F,4);
TASK_PP(16'h1D40,4);
TASK_PP(16'h1D41,4);
TASK_PP(16'h1D42,4);
TASK_PP(16'h1D43,4);
TASK_PP(16'h1D44,4);
TASK_PP(16'h1D45,4);
TASK_PP(16'h1D46,4);
TASK_PP(16'h1D47,4);
TASK_PP(16'h1D48,4);
TASK_PP(16'h1D49,4);
TASK_PP(16'h1D4A,4);
TASK_PP(16'h1D4B,4);
TASK_PP(16'h1D4C,4);
TASK_PP(16'h1D4D,4);
TASK_PP(16'h1D4E,4);
TASK_PP(16'h1D4F,4);
TASK_PP(16'h1D50,4);
TASK_PP(16'h1D51,4);
TASK_PP(16'h1D52,4);
TASK_PP(16'h1D53,4);
TASK_PP(16'h1D54,4);
TASK_PP(16'h1D55,4);
TASK_PP(16'h1D56,4);
TASK_PP(16'h1D57,4);
TASK_PP(16'h1D58,4);
TASK_PP(16'h1D59,4);
TASK_PP(16'h1D5A,4);
TASK_PP(16'h1D5B,4);
TASK_PP(16'h1D5C,4);
TASK_PP(16'h1D5D,4);
TASK_PP(16'h1D5E,4);
TASK_PP(16'h1D5F,4);
TASK_PP(16'h1D60,4);
TASK_PP(16'h1D61,4);
TASK_PP(16'h1D62,4);
TASK_PP(16'h1D63,4);
TASK_PP(16'h1D64,4);
TASK_PP(16'h1D65,4);
TASK_PP(16'h1D66,4);
TASK_PP(16'h1D67,4);
TASK_PP(16'h1D68,4);
TASK_PP(16'h1D69,4);
TASK_PP(16'h1D6A,4);
TASK_PP(16'h1D6B,4);
TASK_PP(16'h1D6C,4);
TASK_PP(16'h1D6D,4);
TASK_PP(16'h1D6E,4);
TASK_PP(16'h1D6F,4);
TASK_PP(16'h1D70,4);
TASK_PP(16'h1D71,4);
TASK_PP(16'h1D72,4);
TASK_PP(16'h1D73,4);
TASK_PP(16'h1D74,4);
TASK_PP(16'h1D75,4);
TASK_PP(16'h1D76,4);
TASK_PP(16'h1D77,4);
TASK_PP(16'h1D78,4);
TASK_PP(16'h1D79,4);
TASK_PP(16'h1D7A,4);
TASK_PP(16'h1D7B,4);
TASK_PP(16'h1D7C,4);
TASK_PP(16'h1D7D,4);
TASK_PP(16'h1D7E,4);
TASK_PP(16'h1D7F,4);
TASK_PP(16'h1D80,4);
TASK_PP(16'h1D81,4);
TASK_PP(16'h1D82,4);
TASK_PP(16'h1D83,4);
TASK_PP(16'h1D84,4);
TASK_PP(16'h1D85,4);
TASK_PP(16'h1D86,4);
TASK_PP(16'h1D87,4);
TASK_PP(16'h1D88,4);
TASK_PP(16'h1D89,4);
TASK_PP(16'h1D8A,4);
TASK_PP(16'h1D8B,4);
TASK_PP(16'h1D8C,4);
TASK_PP(16'h1D8D,4);
TASK_PP(16'h1D8E,4);
TASK_PP(16'h1D8F,4);
TASK_PP(16'h1D90,4);
TASK_PP(16'h1D91,4);
TASK_PP(16'h1D92,4);
TASK_PP(16'h1D93,4);
TASK_PP(16'h1D94,4);
TASK_PP(16'h1D95,4);
TASK_PP(16'h1D96,4);
TASK_PP(16'h1D97,4);
TASK_PP(16'h1D98,4);
TASK_PP(16'h1D99,4);
TASK_PP(16'h1D9A,4);
TASK_PP(16'h1D9B,4);
TASK_PP(16'h1D9C,4);
TASK_PP(16'h1D9D,4);
TASK_PP(16'h1D9E,4);
TASK_PP(16'h1D9F,4);
TASK_PP(16'h1DA0,4);
TASK_PP(16'h1DA1,4);
TASK_PP(16'h1DA2,4);
TASK_PP(16'h1DA3,4);
TASK_PP(16'h1DA4,4);
TASK_PP(16'h1DA5,4);
TASK_PP(16'h1DA6,4);
TASK_PP(16'h1DA7,4);
TASK_PP(16'h1DA8,4);
TASK_PP(16'h1DA9,4);
TASK_PP(16'h1DAA,4);
TASK_PP(16'h1DAB,4);
TASK_PP(16'h1DAC,4);
TASK_PP(16'h1DAD,4);
TASK_PP(16'h1DAE,4);
TASK_PP(16'h1DAF,4);
TASK_PP(16'h1DB0,4);
TASK_PP(16'h1DB1,4);
TASK_PP(16'h1DB2,4);
TASK_PP(16'h1DB3,4);
TASK_PP(16'h1DB4,4);
TASK_PP(16'h1DB5,4);
TASK_PP(16'h1DB6,4);
TASK_PP(16'h1DB7,4);
TASK_PP(16'h1DB8,4);
TASK_PP(16'h1DB9,4);
TASK_PP(16'h1DBA,4);
TASK_PP(16'h1DBB,4);
TASK_PP(16'h1DBC,4);
TASK_PP(16'h1DBD,4);
TASK_PP(16'h1DBE,4);
TASK_PP(16'h1DBF,4);
TASK_PP(16'h1DC0,4);
TASK_PP(16'h1DC1,4);
TASK_PP(16'h1DC2,4);
TASK_PP(16'h1DC3,4);
TASK_PP(16'h1DC4,4);
TASK_PP(16'h1DC5,4);
TASK_PP(16'h1DC6,4);
TASK_PP(16'h1DC7,4);
TASK_PP(16'h1DC8,4);
TASK_PP(16'h1DC9,4);
TASK_PP(16'h1DCA,4);
TASK_PP(16'h1DCB,4);
TASK_PP(16'h1DCC,4);
TASK_PP(16'h1DCD,4);
TASK_PP(16'h1DCE,4);
TASK_PP(16'h1DCF,4);
TASK_PP(16'h1DD0,4);
TASK_PP(16'h1DD1,4);
TASK_PP(16'h1DD2,4);
TASK_PP(16'h1DD3,4);
TASK_PP(16'h1DD4,4);
TASK_PP(16'h1DD5,4);
TASK_PP(16'h1DD6,4);
TASK_PP(16'h1DD7,4);
TASK_PP(16'h1DD8,4);
TASK_PP(16'h1DD9,4);
TASK_PP(16'h1DDA,4);
TASK_PP(16'h1DDB,4);
TASK_PP(16'h1DDC,4);
TASK_PP(16'h1DDD,4);
TASK_PP(16'h1DDE,4);
TASK_PP(16'h1DDF,4);
TASK_PP(16'h1DE0,4);
TASK_PP(16'h1DE1,4);
TASK_PP(16'h1DE2,4);
TASK_PP(16'h1DE3,4);
TASK_PP(16'h1DE4,4);
TASK_PP(16'h1DE5,4);
TASK_PP(16'h1DE6,4);
TASK_PP(16'h1DE7,4);
TASK_PP(16'h1DE8,4);
TASK_PP(16'h1DE9,4);
TASK_PP(16'h1DEA,4);
TASK_PP(16'h1DEB,4);
TASK_PP(16'h1DEC,4);
TASK_PP(16'h1DED,4);
TASK_PP(16'h1DEE,4);
TASK_PP(16'h1DEF,4);
TASK_PP(16'h1DF0,4);
TASK_PP(16'h1DF1,4);
TASK_PP(16'h1DF2,4);
TASK_PP(16'h1DF3,4);
TASK_PP(16'h1DF4,4);
TASK_PP(16'h1DF5,4);
TASK_PP(16'h1DF6,4);
TASK_PP(16'h1DF7,4);
TASK_PP(16'h1DF8,4);
TASK_PP(16'h1DF9,4);
TASK_PP(16'h1DFA,4);
TASK_PP(16'h1DFB,4);
TASK_PP(16'h1DFC,4);
TASK_PP(16'h1DFD,4);
TASK_PP(16'h1DFE,4);
TASK_PP(16'h1DFF,4);
TASK_PP(16'h1E00,4);
TASK_PP(16'h1E01,4);
TASK_PP(16'h1E02,4);
TASK_PP(16'h1E03,4);
TASK_PP(16'h1E04,4);
TASK_PP(16'h1E05,4);
TASK_PP(16'h1E06,4);
TASK_PP(16'h1E07,4);
TASK_PP(16'h1E08,4);
TASK_PP(16'h1E09,4);
TASK_PP(16'h1E0A,4);
TASK_PP(16'h1E0B,4);
TASK_PP(16'h1E0C,4);
TASK_PP(16'h1E0D,4);
TASK_PP(16'h1E0E,4);
TASK_PP(16'h1E0F,4);
TASK_PP(16'h1E10,4);
TASK_PP(16'h1E11,4);
TASK_PP(16'h1E12,4);
TASK_PP(16'h1E13,4);
TASK_PP(16'h1E14,4);
TASK_PP(16'h1E15,4);
TASK_PP(16'h1E16,4);
TASK_PP(16'h1E17,4);
TASK_PP(16'h1E18,4);
TASK_PP(16'h1E19,4);
TASK_PP(16'h1E1A,4);
TASK_PP(16'h1E1B,4);
TASK_PP(16'h1E1C,4);
TASK_PP(16'h1E1D,4);
TASK_PP(16'h1E1E,4);
TASK_PP(16'h1E1F,4);
TASK_PP(16'h1E20,4);
TASK_PP(16'h1E21,4);
TASK_PP(16'h1E22,4);
TASK_PP(16'h1E23,4);
TASK_PP(16'h1E24,4);
TASK_PP(16'h1E25,4);
TASK_PP(16'h1E26,4);
TASK_PP(16'h1E27,4);
TASK_PP(16'h1E28,4);
TASK_PP(16'h1E29,4);
TASK_PP(16'h1E2A,4);
TASK_PP(16'h1E2B,4);
TASK_PP(16'h1E2C,4);
TASK_PP(16'h1E2D,4);
TASK_PP(16'h1E2E,4);
TASK_PP(16'h1E2F,4);
TASK_PP(16'h1E30,4);
TASK_PP(16'h1E31,4);
TASK_PP(16'h1E32,4);
TASK_PP(16'h1E33,4);
TASK_PP(16'h1E34,4);
TASK_PP(16'h1E35,4);
TASK_PP(16'h1E36,4);
TASK_PP(16'h1E37,4);
TASK_PP(16'h1E38,4);
TASK_PP(16'h1E39,4);
TASK_PP(16'h1E3A,4);
TASK_PP(16'h1E3B,4);
TASK_PP(16'h1E3C,4);
TASK_PP(16'h1E3D,4);
TASK_PP(16'h1E3E,4);
TASK_PP(16'h1E3F,4);
TASK_PP(16'h1E40,4);
TASK_PP(16'h1E41,4);
TASK_PP(16'h1E42,4);
TASK_PP(16'h1E43,4);
TASK_PP(16'h1E44,4);
TASK_PP(16'h1E45,4);
TASK_PP(16'h1E46,4);
TASK_PP(16'h1E47,4);
TASK_PP(16'h1E48,4);
TASK_PP(16'h1E49,4);
TASK_PP(16'h1E4A,4);
TASK_PP(16'h1E4B,4);
TASK_PP(16'h1E4C,4);
TASK_PP(16'h1E4D,4);
TASK_PP(16'h1E4E,4);
TASK_PP(16'h1E4F,4);
TASK_PP(16'h1E50,4);
TASK_PP(16'h1E51,4);
TASK_PP(16'h1E52,4);
TASK_PP(16'h1E53,4);
TASK_PP(16'h1E54,4);
TASK_PP(16'h1E55,4);
TASK_PP(16'h1E56,4);
TASK_PP(16'h1E57,4);
TASK_PP(16'h1E58,4);
TASK_PP(16'h1E59,4);
TASK_PP(16'h1E5A,4);
TASK_PP(16'h1E5B,4);
TASK_PP(16'h1E5C,4);
TASK_PP(16'h1E5D,4);
TASK_PP(16'h1E5E,4);
TASK_PP(16'h1E5F,4);
TASK_PP(16'h1E60,4);
TASK_PP(16'h1E61,4);
TASK_PP(16'h1E62,4);
TASK_PP(16'h1E63,4);
TASK_PP(16'h1E64,4);
TASK_PP(16'h1E65,4);
TASK_PP(16'h1E66,4);
TASK_PP(16'h1E67,4);
TASK_PP(16'h1E68,4);
TASK_PP(16'h1E69,4);
TASK_PP(16'h1E6A,4);
TASK_PP(16'h1E6B,4);
TASK_PP(16'h1E6C,4);
TASK_PP(16'h1E6D,4);
TASK_PP(16'h1E6E,4);
TASK_PP(16'h1E6F,4);
TASK_PP(16'h1E70,4);
TASK_PP(16'h1E71,4);
TASK_PP(16'h1E72,4);
TASK_PP(16'h1E73,4);
TASK_PP(16'h1E74,4);
TASK_PP(16'h1E75,4);
TASK_PP(16'h1E76,4);
TASK_PP(16'h1E77,4);
TASK_PP(16'h1E78,4);
TASK_PP(16'h1E79,4);
TASK_PP(16'h1E7A,4);
TASK_PP(16'h1E7B,4);
TASK_PP(16'h1E7C,4);
TASK_PP(16'h1E7D,4);
TASK_PP(16'h1E7E,4);
TASK_PP(16'h1E7F,4);
TASK_PP(16'h1E80,4);
TASK_PP(16'h1E81,4);
TASK_PP(16'h1E82,4);
TASK_PP(16'h1E83,4);
TASK_PP(16'h1E84,4);
TASK_PP(16'h1E85,4);
TASK_PP(16'h1E86,4);
TASK_PP(16'h1E87,4);
TASK_PP(16'h1E88,4);
TASK_PP(16'h1E89,4);
TASK_PP(16'h1E8A,4);
TASK_PP(16'h1E8B,4);
TASK_PP(16'h1E8C,4);
TASK_PP(16'h1E8D,4);
TASK_PP(16'h1E8E,4);
TASK_PP(16'h1E8F,4);
TASK_PP(16'h1E90,4);
TASK_PP(16'h1E91,4);
TASK_PP(16'h1E92,4);
TASK_PP(16'h1E93,4);
TASK_PP(16'h1E94,4);
TASK_PP(16'h1E95,4);
TASK_PP(16'h1E96,4);
TASK_PP(16'h1E97,4);
TASK_PP(16'h1E98,4);
TASK_PP(16'h1E99,4);
TASK_PP(16'h1E9A,4);
TASK_PP(16'h1E9B,4);
TASK_PP(16'h1E9C,4);
TASK_PP(16'h1E9D,4);
TASK_PP(16'h1E9E,4);
TASK_PP(16'h1E9F,4);
TASK_PP(16'h1EA0,4);
TASK_PP(16'h1EA1,4);
TASK_PP(16'h1EA2,4);
TASK_PP(16'h1EA3,4);
TASK_PP(16'h1EA4,4);
TASK_PP(16'h1EA5,4);
TASK_PP(16'h1EA6,4);
TASK_PP(16'h1EA7,4);
TASK_PP(16'h1EA8,4);
TASK_PP(16'h1EA9,4);
TASK_PP(16'h1EAA,4);
TASK_PP(16'h1EAB,4);
TASK_PP(16'h1EAC,4);
TASK_PP(16'h1EAD,4);
TASK_PP(16'h1EAE,4);
TASK_PP(16'h1EAF,4);
TASK_PP(16'h1EB0,4);
TASK_PP(16'h1EB1,4);
TASK_PP(16'h1EB2,4);
TASK_PP(16'h1EB3,4);
TASK_PP(16'h1EB4,4);
TASK_PP(16'h1EB5,4);
TASK_PP(16'h1EB6,4);
TASK_PP(16'h1EB7,4);
TASK_PP(16'h1EB8,4);
TASK_PP(16'h1EB9,4);
TASK_PP(16'h1EBA,4);
TASK_PP(16'h1EBB,4);
TASK_PP(16'h1EBC,4);
TASK_PP(16'h1EBD,4);
TASK_PP(16'h1EBE,4);
TASK_PP(16'h1EBF,4);
TASK_PP(16'h1EC0,4);
TASK_PP(16'h1EC1,4);
TASK_PP(16'h1EC2,4);
TASK_PP(16'h1EC3,4);
TASK_PP(16'h1EC4,4);
TASK_PP(16'h1EC5,4);
TASK_PP(16'h1EC6,4);
TASK_PP(16'h1EC7,4);
TASK_PP(16'h1EC8,4);
TASK_PP(16'h1EC9,4);
TASK_PP(16'h1ECA,4);
TASK_PP(16'h1ECB,4);
TASK_PP(16'h1ECC,4);
TASK_PP(16'h1ECD,4);
TASK_PP(16'h1ECE,4);
TASK_PP(16'h1ECF,4);
TASK_PP(16'h1ED0,4);
TASK_PP(16'h1ED1,4);
TASK_PP(16'h1ED2,4);
TASK_PP(16'h1ED3,4);
TASK_PP(16'h1ED4,4);
TASK_PP(16'h1ED5,4);
TASK_PP(16'h1ED6,4);
TASK_PP(16'h1ED7,4);
TASK_PP(16'h1ED8,4);
TASK_PP(16'h1ED9,4);
TASK_PP(16'h1EDA,4);
TASK_PP(16'h1EDB,4);
TASK_PP(16'h1EDC,4);
TASK_PP(16'h1EDD,4);
TASK_PP(16'h1EDE,4);
TASK_PP(16'h1EDF,4);
TASK_PP(16'h1EE0,4);
TASK_PP(16'h1EE1,4);
TASK_PP(16'h1EE2,4);
TASK_PP(16'h1EE3,4);
TASK_PP(16'h1EE4,4);
TASK_PP(16'h1EE5,4);
TASK_PP(16'h1EE6,4);
TASK_PP(16'h1EE7,4);
TASK_PP(16'h1EE8,4);
TASK_PP(16'h1EE9,4);
TASK_PP(16'h1EEA,4);
TASK_PP(16'h1EEB,4);
TASK_PP(16'h1EEC,4);
TASK_PP(16'h1EED,4);
TASK_PP(16'h1EEE,4);
TASK_PP(16'h1EEF,4);
TASK_PP(16'h1EF0,4);
TASK_PP(16'h1EF1,4);
TASK_PP(16'h1EF2,4);
TASK_PP(16'h1EF3,4);
TASK_PP(16'h1EF4,4);
TASK_PP(16'h1EF5,4);
TASK_PP(16'h1EF6,4);
TASK_PP(16'h1EF7,4);
TASK_PP(16'h1EF8,4);
TASK_PP(16'h1EF9,4);
TASK_PP(16'h1EFA,4);
TASK_PP(16'h1EFB,4);
TASK_PP(16'h1EFC,4);
TASK_PP(16'h1EFD,4);
TASK_PP(16'h1EFE,4);
TASK_PP(16'h1EFF,4);
TASK_PP(16'h1F00,4);
TASK_PP(16'h1F01,4);
TASK_PP(16'h1F02,4);
TASK_PP(16'h1F03,4);
TASK_PP(16'h1F04,4);
TASK_PP(16'h1F05,4);
TASK_PP(16'h1F06,4);
TASK_PP(16'h1F07,4);
TASK_PP(16'h1F08,4);
TASK_PP(16'h1F09,4);
TASK_PP(16'h1F0A,4);
TASK_PP(16'h1F0B,4);
TASK_PP(16'h1F0C,4);
TASK_PP(16'h1F0D,4);
TASK_PP(16'h1F0E,4);
TASK_PP(16'h1F0F,4);
TASK_PP(16'h1F10,4);
TASK_PP(16'h1F11,4);
TASK_PP(16'h1F12,4);
TASK_PP(16'h1F13,4);
TASK_PP(16'h1F14,4);
TASK_PP(16'h1F15,4);
TASK_PP(16'h1F16,4);
TASK_PP(16'h1F17,4);
TASK_PP(16'h1F18,4);
TASK_PP(16'h1F19,4);
TASK_PP(16'h1F1A,4);
TASK_PP(16'h1F1B,4);
TASK_PP(16'h1F1C,4);
TASK_PP(16'h1F1D,4);
TASK_PP(16'h1F1E,4);
TASK_PP(16'h1F1F,4);
TASK_PP(16'h1F20,4);
TASK_PP(16'h1F21,4);
TASK_PP(16'h1F22,4);
TASK_PP(16'h1F23,4);
TASK_PP(16'h1F24,4);
TASK_PP(16'h1F25,4);
TASK_PP(16'h1F26,4);
TASK_PP(16'h1F27,4);
TASK_PP(16'h1F28,4);
TASK_PP(16'h1F29,4);
TASK_PP(16'h1F2A,4);
TASK_PP(16'h1F2B,4);
TASK_PP(16'h1F2C,4);
TASK_PP(16'h1F2D,4);
TASK_PP(16'h1F2E,4);
TASK_PP(16'h1F2F,4);
TASK_PP(16'h1F30,4);
TASK_PP(16'h1F31,4);
TASK_PP(16'h1F32,4);
TASK_PP(16'h1F33,4);
TASK_PP(16'h1F34,4);
TASK_PP(16'h1F35,4);
TASK_PP(16'h1F36,4);
TASK_PP(16'h1F37,4);
TASK_PP(16'h1F38,4);
TASK_PP(16'h1F39,4);
TASK_PP(16'h1F3A,4);
TASK_PP(16'h1F3B,4);
TASK_PP(16'h1F3C,4);
TASK_PP(16'h1F3D,4);
TASK_PP(16'h1F3E,4);
TASK_PP(16'h1F3F,4);
TASK_PP(16'h1F40,4);
TASK_PP(16'h1F41,4);
TASK_PP(16'h1F42,4);
TASK_PP(16'h1F43,4);
TASK_PP(16'h1F44,4);
TASK_PP(16'h1F45,4);
TASK_PP(16'h1F46,4);
TASK_PP(16'h1F47,4);
TASK_PP(16'h1F48,4);
TASK_PP(16'h1F49,4);
TASK_PP(16'h1F4A,4);
TASK_PP(16'h1F4B,4);
TASK_PP(16'h1F4C,4);
TASK_PP(16'h1F4D,4);
TASK_PP(16'h1F4E,4);
TASK_PP(16'h1F4F,4);
TASK_PP(16'h1F50,4);
TASK_PP(16'h1F51,4);
TASK_PP(16'h1F52,4);
TASK_PP(16'h1F53,4);
TASK_PP(16'h1F54,4);
TASK_PP(16'h1F55,4);
TASK_PP(16'h1F56,4);
TASK_PP(16'h1F57,4);
TASK_PP(16'h1F58,4);
TASK_PP(16'h1F59,4);
TASK_PP(16'h1F5A,4);
TASK_PP(16'h1F5B,4);
TASK_PP(16'h1F5C,4);
TASK_PP(16'h1F5D,4);
TASK_PP(16'h1F5E,4);
TASK_PP(16'h1F5F,4);
TASK_PP(16'h1F60,4);
TASK_PP(16'h1F61,4);
TASK_PP(16'h1F62,4);
TASK_PP(16'h1F63,4);
TASK_PP(16'h1F64,4);
TASK_PP(16'h1F65,4);
TASK_PP(16'h1F66,4);
TASK_PP(16'h1F67,4);
TASK_PP(16'h1F68,4);
TASK_PP(16'h1F69,4);
TASK_PP(16'h1F6A,4);
TASK_PP(16'h1F6B,4);
TASK_PP(16'h1F6C,4);
TASK_PP(16'h1F6D,4);
TASK_PP(16'h1F6E,4);
TASK_PP(16'h1F6F,4);
TASK_PP(16'h1F70,4);
TASK_PP(16'h1F71,4);
TASK_PP(16'h1F72,4);
TASK_PP(16'h1F73,4);
TASK_PP(16'h1F74,4);
TASK_PP(16'h1F75,4);
TASK_PP(16'h1F76,4);
TASK_PP(16'h1F77,4);
TASK_PP(16'h1F78,4);
TASK_PP(16'h1F79,4);
TASK_PP(16'h1F7A,4);
TASK_PP(16'h1F7B,4);
TASK_PP(16'h1F7C,4);
TASK_PP(16'h1F7D,4);
TASK_PP(16'h1F7E,4);
TASK_PP(16'h1F7F,4);
TASK_PP(16'h1F80,4);
TASK_PP(16'h1F81,4);
TASK_PP(16'h1F82,4);
TASK_PP(16'h1F83,4);
TASK_PP(16'h1F84,4);
TASK_PP(16'h1F85,4);
TASK_PP(16'h1F86,4);
TASK_PP(16'h1F87,4);
TASK_PP(16'h1F88,4);
TASK_PP(16'h1F89,4);
TASK_PP(16'h1F8A,4);
TASK_PP(16'h1F8B,4);
TASK_PP(16'h1F8C,4);
TASK_PP(16'h1F8D,4);
TASK_PP(16'h1F8E,4);
TASK_PP(16'h1F8F,4);
TASK_PP(16'h1F90,4);
TASK_PP(16'h1F91,4);
TASK_PP(16'h1F92,4);
TASK_PP(16'h1F93,4);
TASK_PP(16'h1F94,4);
TASK_PP(16'h1F95,4);
TASK_PP(16'h1F96,4);
TASK_PP(16'h1F97,4);
TASK_PP(16'h1F98,4);
TASK_PP(16'h1F99,4);
TASK_PP(16'h1F9A,4);
TASK_PP(16'h1F9B,4);
TASK_PP(16'h1F9C,4);
TASK_PP(16'h1F9D,4);
TASK_PP(16'h1F9E,4);
TASK_PP(16'h1F9F,4);
TASK_PP(16'h1FA0,4);
TASK_PP(16'h1FA1,4);
TASK_PP(16'h1FA2,4);
TASK_PP(16'h1FA3,4);
TASK_PP(16'h1FA4,4);
TASK_PP(16'h1FA5,4);
TASK_PP(16'h1FA6,4);
TASK_PP(16'h1FA7,4);
TASK_PP(16'h1FA8,4);
TASK_PP(16'h1FA9,4);
TASK_PP(16'h1FAA,4);
TASK_PP(16'h1FAB,4);
TASK_PP(16'h1FAC,4);
TASK_PP(16'h1FAD,4);
TASK_PP(16'h1FAE,4);
TASK_PP(16'h1FAF,4);
TASK_PP(16'h1FB0,4);
TASK_PP(16'h1FB1,4);
TASK_PP(16'h1FB2,4);
TASK_PP(16'h1FB3,4);
TASK_PP(16'h1FB4,4);
TASK_PP(16'h1FB5,4);
TASK_PP(16'h1FB6,4);
TASK_PP(16'h1FB7,4);
TASK_PP(16'h1FB8,4);
TASK_PP(16'h1FB9,4);
TASK_PP(16'h1FBA,4);
TASK_PP(16'h1FBB,4);
TASK_PP(16'h1FBC,4);
TASK_PP(16'h1FBD,4);
TASK_PP(16'h1FBE,4);
TASK_PP(16'h1FBF,4);
TASK_PP(16'h1FC0,4);
TASK_PP(16'h1FC1,4);
TASK_PP(16'h1FC2,4);
TASK_PP(16'h1FC3,4);
TASK_PP(16'h1FC4,4);
TASK_PP(16'h1FC5,4);
TASK_PP(16'h1FC6,4);
TASK_PP(16'h1FC7,4);
TASK_PP(16'h1FC8,4);
TASK_PP(16'h1FC9,4);
TASK_PP(16'h1FCA,4);
TASK_PP(16'h1FCB,4);
TASK_PP(16'h1FCC,4);
TASK_PP(16'h1FCD,4);
TASK_PP(16'h1FCE,4);
TASK_PP(16'h1FCF,4);
TASK_PP(16'h1FD0,4);
TASK_PP(16'h1FD1,4);
TASK_PP(16'h1FD2,4);
TASK_PP(16'h1FD3,4);
TASK_PP(16'h1FD4,4);
TASK_PP(16'h1FD5,4);
TASK_PP(16'h1FD6,4);
TASK_PP(16'h1FD7,4);
TASK_PP(16'h1FD8,4);
TASK_PP(16'h1FD9,4);
TASK_PP(16'h1FDA,4);
TASK_PP(16'h1FDB,4);
TASK_PP(16'h1FDC,4);
TASK_PP(16'h1FDD,4);
TASK_PP(16'h1FDE,4);
TASK_PP(16'h1FDF,4);
TASK_PP(16'h1FE0,4);
TASK_PP(16'h1FE1,4);
TASK_PP(16'h1FE2,4);
TASK_PP(16'h1FE3,4);
TASK_PP(16'h1FE4,4);
TASK_PP(16'h1FE5,4);
TASK_PP(16'h1FE6,4);
TASK_PP(16'h1FE7,4);
TASK_PP(16'h1FE8,4);
TASK_PP(16'h1FE9,4);
TASK_PP(16'h1FEA,4);
TASK_PP(16'h1FEB,4);
TASK_PP(16'h1FEC,4);
TASK_PP(16'h1FED,4);
TASK_PP(16'h1FEE,4);
TASK_PP(16'h1FEF,4);
TASK_PP(16'h1FF0,4);
TASK_PP(16'h1FF1,4);
TASK_PP(16'h1FF2,4);
TASK_PP(16'h1FF3,4);
TASK_PP(16'h1FF4,4);
TASK_PP(16'h1FF5,4);
TASK_PP(16'h1FF6,4);
TASK_PP(16'h1FF7,4);
TASK_PP(16'h1FF8,4);
TASK_PP(16'h1FF9,4);
TASK_PP(16'h1FFA,4);
TASK_PP(16'h1FFB,4);
TASK_PP(16'h1FFC,4);
TASK_PP(16'h1FFD,4);
TASK_PP(16'h1FFE,4);
TASK_PP(16'h1FFF,4);
TASK_PP(16'h2000,4);
TASK_PP(16'h2001,4);
TASK_PP(16'h2002,4);
TASK_PP(16'h2003,4);
TASK_PP(16'h2004,4);
TASK_PP(16'h2005,4);
TASK_PP(16'h2006,4);
TASK_PP(16'h2007,4);
TASK_PP(16'h2008,4);
TASK_PP(16'h2009,4);
TASK_PP(16'h200A,4);
TASK_PP(16'h200B,4);
TASK_PP(16'h200C,4);
TASK_PP(16'h200D,4);
TASK_PP(16'h200E,4);
TASK_PP(16'h200F,4);
TASK_PP(16'h2010,4);
TASK_PP(16'h2011,4);
TASK_PP(16'h2012,4);
TASK_PP(16'h2013,4);
TASK_PP(16'h2014,4);
TASK_PP(16'h2015,4);
TASK_PP(16'h2016,4);
TASK_PP(16'h2017,4);
TASK_PP(16'h2018,4);
TASK_PP(16'h2019,4);
TASK_PP(16'h201A,4);
TASK_PP(16'h201B,4);
TASK_PP(16'h201C,4);
TASK_PP(16'h201D,4);
TASK_PP(16'h201E,4);
TASK_PP(16'h201F,4);
TASK_PP(16'h2020,4);
TASK_PP(16'h2021,4);
TASK_PP(16'h2022,4);
TASK_PP(16'h2023,4);
TASK_PP(16'h2024,4);
TASK_PP(16'h2025,4);
TASK_PP(16'h2026,4);
TASK_PP(16'h2027,4);
TASK_PP(16'h2028,4);
TASK_PP(16'h2029,4);
TASK_PP(16'h202A,4);
TASK_PP(16'h202B,4);
TASK_PP(16'h202C,4);
TASK_PP(16'h202D,4);
TASK_PP(16'h202E,4);
TASK_PP(16'h202F,4);
TASK_PP(16'h2030,4);
TASK_PP(16'h2031,4);
TASK_PP(16'h2032,4);
TASK_PP(16'h2033,4);
TASK_PP(16'h2034,4);
TASK_PP(16'h2035,4);
TASK_PP(16'h2036,4);
TASK_PP(16'h2037,4);
TASK_PP(16'h2038,4);
TASK_PP(16'h2039,4);
TASK_PP(16'h203A,4);
TASK_PP(16'h203B,4);
TASK_PP(16'h203C,4);
TASK_PP(16'h203D,4);
TASK_PP(16'h203E,4);
TASK_PP(16'h203F,4);
TASK_PP(16'h2040,4);
TASK_PP(16'h2041,4);
TASK_PP(16'h2042,4);
TASK_PP(16'h2043,4);
TASK_PP(16'h2044,4);
TASK_PP(16'h2045,4);
TASK_PP(16'h2046,4);
TASK_PP(16'h2047,4);
TASK_PP(16'h2048,4);
TASK_PP(16'h2049,4);
TASK_PP(16'h204A,4);
TASK_PP(16'h204B,4);
TASK_PP(16'h204C,4);
TASK_PP(16'h204D,4);
TASK_PP(16'h204E,4);
TASK_PP(16'h204F,4);
TASK_PP(16'h2050,4);
TASK_PP(16'h2051,4);
TASK_PP(16'h2052,4);
TASK_PP(16'h2053,4);
TASK_PP(16'h2054,4);
TASK_PP(16'h2055,4);
TASK_PP(16'h2056,4);
TASK_PP(16'h2057,4);
TASK_PP(16'h2058,4);
TASK_PP(16'h2059,4);
TASK_PP(16'h205A,4);
TASK_PP(16'h205B,4);
TASK_PP(16'h205C,4);
TASK_PP(16'h205D,4);
TASK_PP(16'h205E,4);
TASK_PP(16'h205F,4);
TASK_PP(16'h2060,4);
TASK_PP(16'h2061,4);
TASK_PP(16'h2062,4);
TASK_PP(16'h2063,4);
TASK_PP(16'h2064,4);
TASK_PP(16'h2065,4);
TASK_PP(16'h2066,4);
TASK_PP(16'h2067,4);
TASK_PP(16'h2068,4);
TASK_PP(16'h2069,4);
TASK_PP(16'h206A,4);
TASK_PP(16'h206B,4);
TASK_PP(16'h206C,4);
TASK_PP(16'h206D,4);
TASK_PP(16'h206E,4);
TASK_PP(16'h206F,4);
TASK_PP(16'h2070,4);
TASK_PP(16'h2071,4);
TASK_PP(16'h2072,4);
TASK_PP(16'h2073,4);
TASK_PP(16'h2074,4);
TASK_PP(16'h2075,4);
TASK_PP(16'h2076,4);
TASK_PP(16'h2077,4);
TASK_PP(16'h2078,4);
TASK_PP(16'h2079,4);
TASK_PP(16'h207A,4);
TASK_PP(16'h207B,4);
TASK_PP(16'h207C,4);
TASK_PP(16'h207D,4);
TASK_PP(16'h207E,4);
TASK_PP(16'h207F,4);
TASK_PP(16'h2080,4);
TASK_PP(16'h2081,4);
TASK_PP(16'h2082,4);
TASK_PP(16'h2083,4);
TASK_PP(16'h2084,4);
TASK_PP(16'h2085,4);
TASK_PP(16'h2086,4);
TASK_PP(16'h2087,4);
TASK_PP(16'h2088,4);
TASK_PP(16'h2089,4);
TASK_PP(16'h208A,4);
TASK_PP(16'h208B,4);
TASK_PP(16'h208C,4);
TASK_PP(16'h208D,4);
TASK_PP(16'h208E,4);
TASK_PP(16'h208F,4);
TASK_PP(16'h2090,4);
TASK_PP(16'h2091,4);
TASK_PP(16'h2092,4);
TASK_PP(16'h2093,4);
TASK_PP(16'h2094,4);
TASK_PP(16'h2095,4);
TASK_PP(16'h2096,4);
TASK_PP(16'h2097,4);
TASK_PP(16'h2098,4);
TASK_PP(16'h2099,4);
TASK_PP(16'h209A,4);
TASK_PP(16'h209B,4);
TASK_PP(16'h209C,4);
TASK_PP(16'h209D,4);
TASK_PP(16'h209E,4);
TASK_PP(16'h209F,4);
TASK_PP(16'h20A0,4);
TASK_PP(16'h20A1,4);
TASK_PP(16'h20A2,4);
TASK_PP(16'h20A3,4);
TASK_PP(16'h20A4,4);
TASK_PP(16'h20A5,4);
TASK_PP(16'h20A6,4);
TASK_PP(16'h20A7,4);
TASK_PP(16'h20A8,4);
TASK_PP(16'h20A9,4);
TASK_PP(16'h20AA,4);
TASK_PP(16'h20AB,4);
TASK_PP(16'h20AC,4);
TASK_PP(16'h20AD,4);
TASK_PP(16'h20AE,4);
TASK_PP(16'h20AF,4);
TASK_PP(16'h20B0,4);
TASK_PP(16'h20B1,4);
TASK_PP(16'h20B2,4);
TASK_PP(16'h20B3,4);
TASK_PP(16'h20B4,4);
TASK_PP(16'h20B5,4);
TASK_PP(16'h20B6,4);
TASK_PP(16'h20B7,4);
TASK_PP(16'h20B8,4);
TASK_PP(16'h20B9,4);
TASK_PP(16'h20BA,4);
TASK_PP(16'h20BB,4);
TASK_PP(16'h20BC,4);
TASK_PP(16'h20BD,4);
TASK_PP(16'h20BE,4);
TASK_PP(16'h20BF,4);
TASK_PP(16'h20C0,4);
TASK_PP(16'h20C1,4);
TASK_PP(16'h20C2,4);
TASK_PP(16'h20C3,4);
TASK_PP(16'h20C4,4);
TASK_PP(16'h20C5,4);
TASK_PP(16'h20C6,4);
TASK_PP(16'h20C7,4);
TASK_PP(16'h20C8,4);
TASK_PP(16'h20C9,4);
TASK_PP(16'h20CA,4);
TASK_PP(16'h20CB,4);
TASK_PP(16'h20CC,4);
TASK_PP(16'h20CD,4);
TASK_PP(16'h20CE,4);
TASK_PP(16'h20CF,4);
TASK_PP(16'h20D0,4);
TASK_PP(16'h20D1,4);
TASK_PP(16'h20D2,4);
TASK_PP(16'h20D3,4);
TASK_PP(16'h20D4,4);
TASK_PP(16'h20D5,4);
TASK_PP(16'h20D6,4);
TASK_PP(16'h20D7,4);
TASK_PP(16'h20D8,4);
TASK_PP(16'h20D9,4);
TASK_PP(16'h20DA,4);
TASK_PP(16'h20DB,4);
TASK_PP(16'h20DC,4);
TASK_PP(16'h20DD,4);
TASK_PP(16'h20DE,4);
TASK_PP(16'h20DF,4);
TASK_PP(16'h20E0,4);
TASK_PP(16'h20E1,4);
TASK_PP(16'h20E2,4);
TASK_PP(16'h20E3,4);
TASK_PP(16'h20E4,4);
TASK_PP(16'h20E5,4);
TASK_PP(16'h20E6,4);
TASK_PP(16'h20E7,4);
TASK_PP(16'h20E8,4);
TASK_PP(16'h20E9,4);
TASK_PP(16'h20EA,4);
TASK_PP(16'h20EB,4);
TASK_PP(16'h20EC,4);
TASK_PP(16'h20ED,4);
TASK_PP(16'h20EE,4);
TASK_PP(16'h20EF,4);
TASK_PP(16'h20F0,4);
TASK_PP(16'h20F1,4);
TASK_PP(16'h20F2,4);
TASK_PP(16'h20F3,4);
TASK_PP(16'h20F4,4);
TASK_PP(16'h20F5,4);
TASK_PP(16'h20F6,4);
TASK_PP(16'h20F7,4);
TASK_PP(16'h20F8,4);
TASK_PP(16'h20F9,4);
TASK_PP(16'h20FA,4);
TASK_PP(16'h20FB,4);
TASK_PP(16'h20FC,4);
TASK_PP(16'h20FD,4);
TASK_PP(16'h20FE,4);
TASK_PP(16'h20FF,4);
TASK_PP(16'h2100,4);
TASK_PP(16'h2101,4);
TASK_PP(16'h2102,4);
TASK_PP(16'h2103,4);
TASK_PP(16'h2104,4);
TASK_PP(16'h2105,4);
TASK_PP(16'h2106,4);
TASK_PP(16'h2107,4);
TASK_PP(16'h2108,4);
TASK_PP(16'h2109,4);
TASK_PP(16'h210A,4);
TASK_PP(16'h210B,4);
TASK_PP(16'h210C,4);
TASK_PP(16'h210D,4);
TASK_PP(16'h210E,4);
TASK_PP(16'h210F,4);
TASK_PP(16'h2110,4);
TASK_PP(16'h2111,4);
TASK_PP(16'h2112,4);
TASK_PP(16'h2113,4);
TASK_PP(16'h2114,4);
TASK_PP(16'h2115,4);
TASK_PP(16'h2116,4);
TASK_PP(16'h2117,4);
TASK_PP(16'h2118,4);
TASK_PP(16'h2119,4);
TASK_PP(16'h211A,4);
TASK_PP(16'h211B,4);
TASK_PP(16'h211C,4);
TASK_PP(16'h211D,4);
TASK_PP(16'h211E,4);
TASK_PP(16'h211F,4);
TASK_PP(16'h2120,4);
TASK_PP(16'h2121,4);
TASK_PP(16'h2122,4);
TASK_PP(16'h2123,4);
TASK_PP(16'h2124,4);
TASK_PP(16'h2125,4);
TASK_PP(16'h2126,4);
TASK_PP(16'h2127,4);
TASK_PP(16'h2128,4);
TASK_PP(16'h2129,4);
TASK_PP(16'h212A,4);
TASK_PP(16'h212B,4);
TASK_PP(16'h212C,4);
TASK_PP(16'h212D,4);
TASK_PP(16'h212E,4);
TASK_PP(16'h212F,4);
TASK_PP(16'h2130,4);
TASK_PP(16'h2131,4);
TASK_PP(16'h2132,4);
TASK_PP(16'h2133,4);
TASK_PP(16'h2134,4);
TASK_PP(16'h2135,4);
TASK_PP(16'h2136,4);
TASK_PP(16'h2137,4);
TASK_PP(16'h2138,4);
TASK_PP(16'h2139,4);
TASK_PP(16'h213A,4);
TASK_PP(16'h213B,4);
TASK_PP(16'h213C,4);
TASK_PP(16'h213D,4);
TASK_PP(16'h213E,4);
TASK_PP(16'h213F,4);
TASK_PP(16'h2140,4);
TASK_PP(16'h2141,4);
TASK_PP(16'h2142,4);
TASK_PP(16'h2143,4);
TASK_PP(16'h2144,4);
TASK_PP(16'h2145,4);
TASK_PP(16'h2146,4);
TASK_PP(16'h2147,4);
TASK_PP(16'h2148,4);
TASK_PP(16'h2149,4);
TASK_PP(16'h214A,4);
TASK_PP(16'h214B,4);
TASK_PP(16'h214C,4);
TASK_PP(16'h214D,4);
TASK_PP(16'h214E,4);
TASK_PP(16'h214F,4);
TASK_PP(16'h2150,4);
TASK_PP(16'h2151,4);
TASK_PP(16'h2152,4);
TASK_PP(16'h2153,4);
TASK_PP(16'h2154,4);
TASK_PP(16'h2155,4);
TASK_PP(16'h2156,4);
TASK_PP(16'h2157,4);
TASK_PP(16'h2158,4);
TASK_PP(16'h2159,4);
TASK_PP(16'h215A,4);
TASK_PP(16'h215B,4);
TASK_PP(16'h215C,4);
TASK_PP(16'h215D,4);
TASK_PP(16'h215E,4);
TASK_PP(16'h215F,4);
TASK_PP(16'h2160,4);
TASK_PP(16'h2161,4);
TASK_PP(16'h2162,4);
TASK_PP(16'h2163,4);
TASK_PP(16'h2164,4);
TASK_PP(16'h2165,4);
TASK_PP(16'h2166,4);
TASK_PP(16'h2167,4);
TASK_PP(16'h2168,4);
TASK_PP(16'h2169,4);
TASK_PP(16'h216A,4);
TASK_PP(16'h216B,4);
TASK_PP(16'h216C,4);
TASK_PP(16'h216D,4);
TASK_PP(16'h216E,4);
TASK_PP(16'h216F,4);
TASK_PP(16'h2170,4);
TASK_PP(16'h2171,4);
TASK_PP(16'h2172,4);
TASK_PP(16'h2173,4);
TASK_PP(16'h2174,4);
TASK_PP(16'h2175,4);
TASK_PP(16'h2176,4);
TASK_PP(16'h2177,4);
TASK_PP(16'h2178,4);
TASK_PP(16'h2179,4);
TASK_PP(16'h217A,4);
TASK_PP(16'h217B,4);
TASK_PP(16'h217C,4);
TASK_PP(16'h217D,4);
TASK_PP(16'h217E,4);
TASK_PP(16'h217F,4);
TASK_PP(16'h2180,4);
TASK_PP(16'h2181,4);
TASK_PP(16'h2182,4);
TASK_PP(16'h2183,4);
TASK_PP(16'h2184,4);
TASK_PP(16'h2185,4);
TASK_PP(16'h2186,4);
TASK_PP(16'h2187,4);
TASK_PP(16'h2188,4);
TASK_PP(16'h2189,4);
TASK_PP(16'h218A,4);
TASK_PP(16'h218B,4);
TASK_PP(16'h218C,4);
TASK_PP(16'h218D,4);
TASK_PP(16'h218E,4);
TASK_PP(16'h218F,4);
TASK_PP(16'h2190,4);
TASK_PP(16'h2191,4);
TASK_PP(16'h2192,4);
TASK_PP(16'h2193,4);
TASK_PP(16'h2194,4);
TASK_PP(16'h2195,4);
TASK_PP(16'h2196,4);
TASK_PP(16'h2197,4);
TASK_PP(16'h2198,4);
TASK_PP(16'h2199,4);
TASK_PP(16'h219A,4);
TASK_PP(16'h219B,4);
TASK_PP(16'h219C,4);
TASK_PP(16'h219D,4);
TASK_PP(16'h219E,4);
TASK_PP(16'h219F,4);
TASK_PP(16'h21A0,4);
TASK_PP(16'h21A1,4);
TASK_PP(16'h21A2,4);
TASK_PP(16'h21A3,4);
TASK_PP(16'h21A4,4);
TASK_PP(16'h21A5,4);
TASK_PP(16'h21A6,4);
TASK_PP(16'h21A7,4);
TASK_PP(16'h21A8,4);
TASK_PP(16'h21A9,4);
TASK_PP(16'h21AA,4);
TASK_PP(16'h21AB,4);
TASK_PP(16'h21AC,4);
TASK_PP(16'h21AD,4);
TASK_PP(16'h21AE,4);
TASK_PP(16'h21AF,4);
TASK_PP(16'h21B0,4);
TASK_PP(16'h21B1,4);
TASK_PP(16'h21B2,4);
TASK_PP(16'h21B3,4);
TASK_PP(16'h21B4,4);
TASK_PP(16'h21B5,4);
TASK_PP(16'h21B6,4);
TASK_PP(16'h21B7,4);
TASK_PP(16'h21B8,4);
TASK_PP(16'h21B9,4);
TASK_PP(16'h21BA,4);
TASK_PP(16'h21BB,4);
TASK_PP(16'h21BC,4);
TASK_PP(16'h21BD,4);
TASK_PP(16'h21BE,4);
TASK_PP(16'h21BF,4);
TASK_PP(16'h21C0,4);
TASK_PP(16'h21C1,4);
TASK_PP(16'h21C2,4);
TASK_PP(16'h21C3,4);
TASK_PP(16'h21C4,4);
TASK_PP(16'h21C5,4);
TASK_PP(16'h21C6,4);
TASK_PP(16'h21C7,4);
TASK_PP(16'h21C8,4);
TASK_PP(16'h21C9,4);
TASK_PP(16'h21CA,4);
TASK_PP(16'h21CB,4);
TASK_PP(16'h21CC,4);
TASK_PP(16'h21CD,4);
TASK_PP(16'h21CE,4);
TASK_PP(16'h21CF,4);
TASK_PP(16'h21D0,4);
TASK_PP(16'h21D1,4);
TASK_PP(16'h21D2,4);
TASK_PP(16'h21D3,4);
TASK_PP(16'h21D4,4);
TASK_PP(16'h21D5,4);
TASK_PP(16'h21D6,4);
TASK_PP(16'h21D7,4);
TASK_PP(16'h21D8,4);
TASK_PP(16'h21D9,4);
TASK_PP(16'h21DA,4);
TASK_PP(16'h21DB,4);
TASK_PP(16'h21DC,4);
TASK_PP(16'h21DD,4);
TASK_PP(16'h21DE,4);
TASK_PP(16'h21DF,4);
TASK_PP(16'h21E0,4);
TASK_PP(16'h21E1,4);
TASK_PP(16'h21E2,4);
TASK_PP(16'h21E3,4);
TASK_PP(16'h21E4,4);
TASK_PP(16'h21E5,4);
TASK_PP(16'h21E6,4);
TASK_PP(16'h21E7,4);
TASK_PP(16'h21E8,4);
TASK_PP(16'h21E9,4);
TASK_PP(16'h21EA,4);
TASK_PP(16'h21EB,4);
TASK_PP(16'h21EC,4);
TASK_PP(16'h21ED,4);
TASK_PP(16'h21EE,4);
TASK_PP(16'h21EF,4);
TASK_PP(16'h21F0,4);
TASK_PP(16'h21F1,4);
TASK_PP(16'h21F2,4);
TASK_PP(16'h21F3,4);
TASK_PP(16'h21F4,4);
TASK_PP(16'h21F5,4);
TASK_PP(16'h21F6,4);
TASK_PP(16'h21F7,4);
TASK_PP(16'h21F8,4);
TASK_PP(16'h21F9,4);
TASK_PP(16'h21FA,4);
TASK_PP(16'h21FB,4);
TASK_PP(16'h21FC,4);
TASK_PP(16'h21FD,4);
TASK_PP(16'h21FE,4);
TASK_PP(16'h21FF,4);
TASK_PP(16'h2200,4);
TASK_PP(16'h2201,4);
TASK_PP(16'h2202,4);
TASK_PP(16'h2203,4);
TASK_PP(16'h2204,4);
TASK_PP(16'h2205,4);
TASK_PP(16'h2206,4);
TASK_PP(16'h2207,4);
TASK_PP(16'h2208,4);
TASK_PP(16'h2209,4);
TASK_PP(16'h220A,4);
TASK_PP(16'h220B,4);
TASK_PP(16'h220C,4);
TASK_PP(16'h220D,4);
TASK_PP(16'h220E,4);
TASK_PP(16'h220F,4);
TASK_PP(16'h2210,4);
TASK_PP(16'h2211,4);
TASK_PP(16'h2212,4);
TASK_PP(16'h2213,4);
TASK_PP(16'h2214,4);
TASK_PP(16'h2215,4);
TASK_PP(16'h2216,4);
TASK_PP(16'h2217,4);
TASK_PP(16'h2218,4);
TASK_PP(16'h2219,4);
TASK_PP(16'h221A,4);
TASK_PP(16'h221B,4);
TASK_PP(16'h221C,4);
TASK_PP(16'h221D,4);
TASK_PP(16'h221E,4);
TASK_PP(16'h221F,4);
TASK_PP(16'h2220,4);
TASK_PP(16'h2221,4);
TASK_PP(16'h2222,4);
TASK_PP(16'h2223,4);
TASK_PP(16'h2224,4);
TASK_PP(16'h2225,4);
TASK_PP(16'h2226,4);
TASK_PP(16'h2227,4);
TASK_PP(16'h2228,4);
TASK_PP(16'h2229,4);
TASK_PP(16'h222A,4);
TASK_PP(16'h222B,4);
TASK_PP(16'h222C,4);
TASK_PP(16'h222D,4);
TASK_PP(16'h222E,4);
TASK_PP(16'h222F,4);
TASK_PP(16'h2230,4);
TASK_PP(16'h2231,4);
TASK_PP(16'h2232,4);
TASK_PP(16'h2233,4);
TASK_PP(16'h2234,4);
TASK_PP(16'h2235,4);
TASK_PP(16'h2236,4);
TASK_PP(16'h2237,4);
TASK_PP(16'h2238,4);
TASK_PP(16'h2239,4);
TASK_PP(16'h223A,4);
TASK_PP(16'h223B,4);
TASK_PP(16'h223C,4);
TASK_PP(16'h223D,4);
TASK_PP(16'h223E,4);
TASK_PP(16'h223F,4);
TASK_PP(16'h2240,4);
TASK_PP(16'h2241,4);
TASK_PP(16'h2242,4);
TASK_PP(16'h2243,4);
TASK_PP(16'h2244,4);
TASK_PP(16'h2245,4);
TASK_PP(16'h2246,4);
TASK_PP(16'h2247,4);
TASK_PP(16'h2248,4);
TASK_PP(16'h2249,4);
TASK_PP(16'h224A,4);
TASK_PP(16'h224B,4);
TASK_PP(16'h224C,4);
TASK_PP(16'h224D,4);
TASK_PP(16'h224E,4);
TASK_PP(16'h224F,4);
TASK_PP(16'h2250,4);
TASK_PP(16'h2251,4);
TASK_PP(16'h2252,4);
TASK_PP(16'h2253,4);
TASK_PP(16'h2254,4);
TASK_PP(16'h2255,4);
TASK_PP(16'h2256,4);
TASK_PP(16'h2257,4);
TASK_PP(16'h2258,4);
TASK_PP(16'h2259,4);
TASK_PP(16'h225A,4);
TASK_PP(16'h225B,4);
TASK_PP(16'h225C,4);
TASK_PP(16'h225D,4);
TASK_PP(16'h225E,4);
TASK_PP(16'h225F,4);
TASK_PP(16'h2260,4);
TASK_PP(16'h2261,4);
TASK_PP(16'h2262,4);
TASK_PP(16'h2263,4);
TASK_PP(16'h2264,4);
TASK_PP(16'h2265,4);
TASK_PP(16'h2266,4);
TASK_PP(16'h2267,4);
TASK_PP(16'h2268,4);
TASK_PP(16'h2269,4);
TASK_PP(16'h226A,4);
TASK_PP(16'h226B,4);
TASK_PP(16'h226C,4);
TASK_PP(16'h226D,4);
TASK_PP(16'h226E,4);
TASK_PP(16'h226F,4);
TASK_PP(16'h2270,4);
TASK_PP(16'h2271,4);
TASK_PP(16'h2272,4);
TASK_PP(16'h2273,4);
TASK_PP(16'h2274,4);
TASK_PP(16'h2275,4);
TASK_PP(16'h2276,4);
TASK_PP(16'h2277,4);
TASK_PP(16'h2278,4);
TASK_PP(16'h2279,4);
TASK_PP(16'h227A,4);
TASK_PP(16'h227B,4);
TASK_PP(16'h227C,4);
TASK_PP(16'h227D,4);
TASK_PP(16'h227E,4);
TASK_PP(16'h227F,4);
TASK_PP(16'h2280,4);
TASK_PP(16'h2281,4);
TASK_PP(16'h2282,4);
TASK_PP(16'h2283,4);
TASK_PP(16'h2284,4);
TASK_PP(16'h2285,4);
TASK_PP(16'h2286,4);
TASK_PP(16'h2287,4);
TASK_PP(16'h2288,4);
TASK_PP(16'h2289,4);
TASK_PP(16'h228A,4);
TASK_PP(16'h228B,4);
TASK_PP(16'h228C,4);
TASK_PP(16'h228D,4);
TASK_PP(16'h228E,4);
TASK_PP(16'h228F,4);
TASK_PP(16'h2290,4);
TASK_PP(16'h2291,4);
TASK_PP(16'h2292,4);
TASK_PP(16'h2293,4);
TASK_PP(16'h2294,4);
TASK_PP(16'h2295,4);
TASK_PP(16'h2296,4);
TASK_PP(16'h2297,4);
TASK_PP(16'h2298,4);
TASK_PP(16'h2299,4);
TASK_PP(16'h229A,4);
TASK_PP(16'h229B,4);
TASK_PP(16'h229C,4);
TASK_PP(16'h229D,4);
TASK_PP(16'h229E,4);
TASK_PP(16'h229F,4);
TASK_PP(16'h22A0,4);
TASK_PP(16'h22A1,4);
TASK_PP(16'h22A2,4);
TASK_PP(16'h22A3,4);
TASK_PP(16'h22A4,4);
TASK_PP(16'h22A5,4);
TASK_PP(16'h22A6,4);
TASK_PP(16'h22A7,4);
TASK_PP(16'h22A8,4);
TASK_PP(16'h22A9,4);
TASK_PP(16'h22AA,4);
TASK_PP(16'h22AB,4);
TASK_PP(16'h22AC,4);
TASK_PP(16'h22AD,4);
TASK_PP(16'h22AE,4);
TASK_PP(16'h22AF,4);
TASK_PP(16'h22B0,4);
TASK_PP(16'h22B1,4);
TASK_PP(16'h22B2,4);
TASK_PP(16'h22B3,4);
TASK_PP(16'h22B4,4);
TASK_PP(16'h22B5,4);
TASK_PP(16'h22B6,4);
TASK_PP(16'h22B7,4);
TASK_PP(16'h22B8,4);
TASK_PP(16'h22B9,4);
TASK_PP(16'h22BA,4);
TASK_PP(16'h22BB,4);
TASK_PP(16'h22BC,4);
TASK_PP(16'h22BD,4);
TASK_PP(16'h22BE,4);
TASK_PP(16'h22BF,4);
TASK_PP(16'h22C0,4);
TASK_PP(16'h22C1,4);
TASK_PP(16'h22C2,4);
TASK_PP(16'h22C3,4);
TASK_PP(16'h22C4,4);
TASK_PP(16'h22C5,4);
TASK_PP(16'h22C6,4);
TASK_PP(16'h22C7,4);
TASK_PP(16'h22C8,4);
TASK_PP(16'h22C9,4);
TASK_PP(16'h22CA,4);
TASK_PP(16'h22CB,4);
TASK_PP(16'h22CC,4);
TASK_PP(16'h22CD,4);
TASK_PP(16'h22CE,4);
TASK_PP(16'h22CF,4);
TASK_PP(16'h22D0,4);
TASK_PP(16'h22D1,4);
TASK_PP(16'h22D2,4);
TASK_PP(16'h22D3,4);
TASK_PP(16'h22D4,4);
TASK_PP(16'h22D5,4);
TASK_PP(16'h22D6,4);
TASK_PP(16'h22D7,4);
TASK_PP(16'h22D8,4);
TASK_PP(16'h22D9,4);
TASK_PP(16'h22DA,4);
TASK_PP(16'h22DB,4);
TASK_PP(16'h22DC,4);
TASK_PP(16'h22DD,4);
TASK_PP(16'h22DE,4);
TASK_PP(16'h22DF,4);
TASK_PP(16'h22E0,4);
TASK_PP(16'h22E1,4);
TASK_PP(16'h22E2,4);
TASK_PP(16'h22E3,4);
TASK_PP(16'h22E4,4);
TASK_PP(16'h22E5,4);
TASK_PP(16'h22E6,4);
TASK_PP(16'h22E7,4);
TASK_PP(16'h22E8,4);
TASK_PP(16'h22E9,4);
TASK_PP(16'h22EA,4);
TASK_PP(16'h22EB,4);
TASK_PP(16'h22EC,4);
TASK_PP(16'h22ED,4);
TASK_PP(16'h22EE,4);
TASK_PP(16'h22EF,4);
TASK_PP(16'h22F0,4);
TASK_PP(16'h22F1,4);
TASK_PP(16'h22F2,4);
TASK_PP(16'h22F3,4);
TASK_PP(16'h22F4,4);
TASK_PP(16'h22F5,4);
TASK_PP(16'h22F6,4);
TASK_PP(16'h22F7,4);
TASK_PP(16'h22F8,4);
TASK_PP(16'h22F9,4);
TASK_PP(16'h22FA,4);
TASK_PP(16'h22FB,4);
TASK_PP(16'h22FC,4);
TASK_PP(16'h22FD,4);
TASK_PP(16'h22FE,4);
TASK_PP(16'h22FF,4);
TASK_PP(16'h2300,4);
TASK_PP(16'h2301,4);
TASK_PP(16'h2302,4);
TASK_PP(16'h2303,4);
TASK_PP(16'h2304,4);
TASK_PP(16'h2305,4);
TASK_PP(16'h2306,4);
TASK_PP(16'h2307,4);
TASK_PP(16'h2308,4);
TASK_PP(16'h2309,4);
TASK_PP(16'h230A,4);
TASK_PP(16'h230B,4);
TASK_PP(16'h230C,4);
TASK_PP(16'h230D,4);
TASK_PP(16'h230E,4);
TASK_PP(16'h230F,4);
TASK_PP(16'h2310,4);
TASK_PP(16'h2311,4);
TASK_PP(16'h2312,4);
TASK_PP(16'h2313,4);
TASK_PP(16'h2314,4);
TASK_PP(16'h2315,4);
TASK_PP(16'h2316,4);
TASK_PP(16'h2317,4);
TASK_PP(16'h2318,4);
TASK_PP(16'h2319,4);
TASK_PP(16'h231A,4);
TASK_PP(16'h231B,4);
TASK_PP(16'h231C,4);
TASK_PP(16'h231D,4);
TASK_PP(16'h231E,4);
TASK_PP(16'h231F,4);
TASK_PP(16'h2320,4);
TASK_PP(16'h2321,4);
TASK_PP(16'h2322,4);
TASK_PP(16'h2323,4);
TASK_PP(16'h2324,4);
TASK_PP(16'h2325,4);
TASK_PP(16'h2326,4);
TASK_PP(16'h2327,4);
TASK_PP(16'h2328,4);
TASK_PP(16'h2329,4);
TASK_PP(16'h232A,4);
TASK_PP(16'h232B,4);
TASK_PP(16'h232C,4);
TASK_PP(16'h232D,4);
TASK_PP(16'h232E,4);
TASK_PP(16'h232F,4);
TASK_PP(16'h2330,4);
TASK_PP(16'h2331,4);
TASK_PP(16'h2332,4);
TASK_PP(16'h2333,4);
TASK_PP(16'h2334,4);
TASK_PP(16'h2335,4);
TASK_PP(16'h2336,4);
TASK_PP(16'h2337,4);
TASK_PP(16'h2338,4);
TASK_PP(16'h2339,4);
TASK_PP(16'h233A,4);
TASK_PP(16'h233B,4);
TASK_PP(16'h233C,4);
TASK_PP(16'h233D,4);
TASK_PP(16'h233E,4);
TASK_PP(16'h233F,4);
TASK_PP(16'h2340,4);
TASK_PP(16'h2341,4);
TASK_PP(16'h2342,4);
TASK_PP(16'h2343,4);
TASK_PP(16'h2344,4);
TASK_PP(16'h2345,4);
TASK_PP(16'h2346,4);
TASK_PP(16'h2347,4);
TASK_PP(16'h2348,4);
TASK_PP(16'h2349,4);
TASK_PP(16'h234A,4);
TASK_PP(16'h234B,4);
TASK_PP(16'h234C,4);
TASK_PP(16'h234D,4);
TASK_PP(16'h234E,4);
TASK_PP(16'h234F,4);
TASK_PP(16'h2350,4);
TASK_PP(16'h2351,4);
TASK_PP(16'h2352,4);
TASK_PP(16'h2353,4);
TASK_PP(16'h2354,4);
TASK_PP(16'h2355,4);
TASK_PP(16'h2356,4);
TASK_PP(16'h2357,4);
TASK_PP(16'h2358,4);
TASK_PP(16'h2359,4);
TASK_PP(16'h235A,4);
TASK_PP(16'h235B,4);
TASK_PP(16'h235C,4);
TASK_PP(16'h235D,4);
TASK_PP(16'h235E,4);
TASK_PP(16'h235F,4);
TASK_PP(16'h2360,4);
TASK_PP(16'h2361,4);
TASK_PP(16'h2362,4);
TASK_PP(16'h2363,4);
TASK_PP(16'h2364,4);
TASK_PP(16'h2365,4);
TASK_PP(16'h2366,4);
TASK_PP(16'h2367,4);
TASK_PP(16'h2368,4);
TASK_PP(16'h2369,4);
TASK_PP(16'h236A,4);
TASK_PP(16'h236B,4);
TASK_PP(16'h236C,4);
TASK_PP(16'h236D,4);
TASK_PP(16'h236E,4);
TASK_PP(16'h236F,4);
TASK_PP(16'h2370,4);
TASK_PP(16'h2371,4);
TASK_PP(16'h2372,4);
TASK_PP(16'h2373,4);
TASK_PP(16'h2374,4);
TASK_PP(16'h2375,4);
TASK_PP(16'h2376,4);
TASK_PP(16'h2377,4);
TASK_PP(16'h2378,4);
TASK_PP(16'h2379,4);
TASK_PP(16'h237A,4);
TASK_PP(16'h237B,4);
TASK_PP(16'h237C,4);
TASK_PP(16'h237D,4);
TASK_PP(16'h237E,4);
TASK_PP(16'h237F,4);
TASK_PP(16'h2380,4);
TASK_PP(16'h2381,4);
TASK_PP(16'h2382,4);
TASK_PP(16'h2383,4);
TASK_PP(16'h2384,4);
TASK_PP(16'h2385,4);
TASK_PP(16'h2386,4);
TASK_PP(16'h2387,4);
TASK_PP(16'h2388,4);
TASK_PP(16'h2389,4);
TASK_PP(16'h238A,4);
TASK_PP(16'h238B,4);
TASK_PP(16'h238C,4);
TASK_PP(16'h238D,4);
TASK_PP(16'h238E,4);
TASK_PP(16'h238F,4);
TASK_PP(16'h2390,4);
TASK_PP(16'h2391,4);
TASK_PP(16'h2392,4);
TASK_PP(16'h2393,4);
TASK_PP(16'h2394,4);
TASK_PP(16'h2395,4);
TASK_PP(16'h2396,4);
TASK_PP(16'h2397,4);
TASK_PP(16'h2398,4);
TASK_PP(16'h2399,4);
TASK_PP(16'h239A,4);
TASK_PP(16'h239B,4);
TASK_PP(16'h239C,4);
TASK_PP(16'h239D,4);
TASK_PP(16'h239E,4);
TASK_PP(16'h239F,4);
TASK_PP(16'h23A0,4);
TASK_PP(16'h23A1,4);
TASK_PP(16'h23A2,4);
TASK_PP(16'h23A3,4);
TASK_PP(16'h23A4,4);
TASK_PP(16'h23A5,4);
TASK_PP(16'h23A6,4);
TASK_PP(16'h23A7,4);
TASK_PP(16'h23A8,4);
TASK_PP(16'h23A9,4);
TASK_PP(16'h23AA,4);
TASK_PP(16'h23AB,4);
TASK_PP(16'h23AC,4);
TASK_PP(16'h23AD,4);
TASK_PP(16'h23AE,4);
TASK_PP(16'h23AF,4);
TASK_PP(16'h23B0,4);
TASK_PP(16'h23B1,4);
TASK_PP(16'h23B2,4);
TASK_PP(16'h23B3,4);
TASK_PP(16'h23B4,4);
TASK_PP(16'h23B5,4);
TASK_PP(16'h23B6,4);
TASK_PP(16'h23B7,4);
TASK_PP(16'h23B8,4);
TASK_PP(16'h23B9,4);
TASK_PP(16'h23BA,4);
TASK_PP(16'h23BB,4);
TASK_PP(16'h23BC,4);
TASK_PP(16'h23BD,4);
TASK_PP(16'h23BE,4);
TASK_PP(16'h23BF,4);
TASK_PP(16'h23C0,4);
TASK_PP(16'h23C1,4);
TASK_PP(16'h23C2,4);
TASK_PP(16'h23C3,4);
TASK_PP(16'h23C4,4);
TASK_PP(16'h23C5,4);
TASK_PP(16'h23C6,4);
TASK_PP(16'h23C7,4);
TASK_PP(16'h23C8,4);
TASK_PP(16'h23C9,4);
TASK_PP(16'h23CA,4);
TASK_PP(16'h23CB,4);
TASK_PP(16'h23CC,4);
TASK_PP(16'h23CD,4);
TASK_PP(16'h23CE,4);
TASK_PP(16'h23CF,4);
TASK_PP(16'h23D0,4);
TASK_PP(16'h23D1,4);
TASK_PP(16'h23D2,4);
TASK_PP(16'h23D3,4);
TASK_PP(16'h23D4,4);
TASK_PP(16'h23D5,4);
TASK_PP(16'h23D6,4);
TASK_PP(16'h23D7,4);
TASK_PP(16'h23D8,4);
TASK_PP(16'h23D9,4);
TASK_PP(16'h23DA,4);
TASK_PP(16'h23DB,4);
TASK_PP(16'h23DC,4);
TASK_PP(16'h23DD,4);
TASK_PP(16'h23DE,4);
TASK_PP(16'h23DF,4);
TASK_PP(16'h23E0,4);
TASK_PP(16'h23E1,4);
TASK_PP(16'h23E2,4);
TASK_PP(16'h23E3,4);
TASK_PP(16'h23E4,4);
TASK_PP(16'h23E5,4);
TASK_PP(16'h23E6,4);
TASK_PP(16'h23E7,4);
TASK_PP(16'h23E8,4);
TASK_PP(16'h23E9,4);
TASK_PP(16'h23EA,4);
TASK_PP(16'h23EB,4);
TASK_PP(16'h23EC,4);
TASK_PP(16'h23ED,4);
TASK_PP(16'h23EE,4);
TASK_PP(16'h23EF,4);
TASK_PP(16'h23F0,4);
TASK_PP(16'h23F1,4);
TASK_PP(16'h23F2,4);
TASK_PP(16'h23F3,4);
TASK_PP(16'h23F4,4);
TASK_PP(16'h23F5,4);
TASK_PP(16'h23F6,4);
TASK_PP(16'h23F7,4);
TASK_PP(16'h23F8,4);
TASK_PP(16'h23F9,4);
TASK_PP(16'h23FA,4);
TASK_PP(16'h23FB,4);
TASK_PP(16'h23FC,4);
TASK_PP(16'h23FD,4);
TASK_PP(16'h23FE,4);
TASK_PP(16'h23FF,4);
TASK_PP(16'h2400,4);
TASK_PP(16'h2401,4);
TASK_PP(16'h2402,4);
TASK_PP(16'h2403,4);
TASK_PP(16'h2404,4);
TASK_PP(16'h2405,4);
TASK_PP(16'h2406,4);
TASK_PP(16'h2407,4);
TASK_PP(16'h2408,4);
TASK_PP(16'h2409,4);
TASK_PP(16'h240A,4);
TASK_PP(16'h240B,4);
TASK_PP(16'h240C,4);
TASK_PP(16'h240D,4);
TASK_PP(16'h240E,4);
TASK_PP(16'h240F,4);
TASK_PP(16'h2410,4);
TASK_PP(16'h2411,4);
TASK_PP(16'h2412,4);
TASK_PP(16'h2413,4);
TASK_PP(16'h2414,4);
TASK_PP(16'h2415,4);
TASK_PP(16'h2416,4);
TASK_PP(16'h2417,4);
TASK_PP(16'h2418,4);
TASK_PP(16'h2419,4);
TASK_PP(16'h241A,4);
TASK_PP(16'h241B,4);
TASK_PP(16'h241C,4);
TASK_PP(16'h241D,4);
TASK_PP(16'h241E,4);
TASK_PP(16'h241F,4);
TASK_PP(16'h2420,4);
TASK_PP(16'h2421,4);
TASK_PP(16'h2422,4);
TASK_PP(16'h2423,4);
TASK_PP(16'h2424,4);
TASK_PP(16'h2425,4);
TASK_PP(16'h2426,4);
TASK_PP(16'h2427,4);
TASK_PP(16'h2428,4);
TASK_PP(16'h2429,4);
TASK_PP(16'h242A,4);
TASK_PP(16'h242B,4);
TASK_PP(16'h242C,4);
TASK_PP(16'h242D,4);
TASK_PP(16'h242E,4);
TASK_PP(16'h242F,4);
TASK_PP(16'h2430,4);
TASK_PP(16'h2431,4);
TASK_PP(16'h2432,4);
TASK_PP(16'h2433,4);
TASK_PP(16'h2434,4);
TASK_PP(16'h2435,4);
TASK_PP(16'h2436,4);
TASK_PP(16'h2437,4);
TASK_PP(16'h2438,4);
TASK_PP(16'h2439,4);
TASK_PP(16'h243A,4);
TASK_PP(16'h243B,4);
TASK_PP(16'h243C,4);
TASK_PP(16'h243D,4);
TASK_PP(16'h243E,4);
TASK_PP(16'h243F,4);
TASK_PP(16'h2440,4);
TASK_PP(16'h2441,4);
TASK_PP(16'h2442,4);
TASK_PP(16'h2443,4);
TASK_PP(16'h2444,4);
TASK_PP(16'h2445,4);
TASK_PP(16'h2446,4);
TASK_PP(16'h2447,4);
TASK_PP(16'h2448,4);
TASK_PP(16'h2449,4);
TASK_PP(16'h244A,4);
TASK_PP(16'h244B,4);
TASK_PP(16'h244C,4);
TASK_PP(16'h244D,4);
TASK_PP(16'h244E,4);
TASK_PP(16'h244F,4);
TASK_PP(16'h2450,4);
TASK_PP(16'h2451,4);
TASK_PP(16'h2452,4);
TASK_PP(16'h2453,4);
TASK_PP(16'h2454,4);
TASK_PP(16'h2455,4);
TASK_PP(16'h2456,4);
TASK_PP(16'h2457,4);
TASK_PP(16'h2458,4);
TASK_PP(16'h2459,4);
TASK_PP(16'h245A,4);
TASK_PP(16'h245B,4);
TASK_PP(16'h245C,4);
TASK_PP(16'h245D,4);
TASK_PP(16'h245E,4);
TASK_PP(16'h245F,4);
TASK_PP(16'h2460,4);
TASK_PP(16'h2461,4);
TASK_PP(16'h2462,4);
TASK_PP(16'h2463,4);
TASK_PP(16'h2464,4);
TASK_PP(16'h2465,4);
TASK_PP(16'h2466,4);
TASK_PP(16'h2467,4);
TASK_PP(16'h2468,4);
TASK_PP(16'h2469,4);
TASK_PP(16'h246A,4);
TASK_PP(16'h246B,4);
TASK_PP(16'h246C,4);
TASK_PP(16'h246D,4);
TASK_PP(16'h246E,4);
TASK_PP(16'h246F,4);
TASK_PP(16'h2470,4);
TASK_PP(16'h2471,4);
TASK_PP(16'h2472,4);
TASK_PP(16'h2473,4);
TASK_PP(16'h2474,4);
TASK_PP(16'h2475,4);
TASK_PP(16'h2476,4);
TASK_PP(16'h2477,4);
TASK_PP(16'h2478,4);
TASK_PP(16'h2479,4);
TASK_PP(16'h247A,4);
TASK_PP(16'h247B,4);
TASK_PP(16'h247C,4);
TASK_PP(16'h247D,4);
TASK_PP(16'h247E,4);
TASK_PP(16'h247F,4);
TASK_PP(16'h2480,4);
TASK_PP(16'h2481,4);
TASK_PP(16'h2482,4);
TASK_PP(16'h2483,4);
TASK_PP(16'h2484,4);
TASK_PP(16'h2485,4);
TASK_PP(16'h2486,4);
TASK_PP(16'h2487,4);
TASK_PP(16'h2488,4);
TASK_PP(16'h2489,4);
TASK_PP(16'h248A,4);
TASK_PP(16'h248B,4);
TASK_PP(16'h248C,4);
TASK_PP(16'h248D,4);
TASK_PP(16'h248E,4);
TASK_PP(16'h248F,4);
TASK_PP(16'h2490,4);
TASK_PP(16'h2491,4);
TASK_PP(16'h2492,4);
TASK_PP(16'h2493,4);
TASK_PP(16'h2494,4);
TASK_PP(16'h2495,4);
TASK_PP(16'h2496,4);
TASK_PP(16'h2497,4);
TASK_PP(16'h2498,4);
TASK_PP(16'h2499,4);
TASK_PP(16'h249A,4);
TASK_PP(16'h249B,4);
TASK_PP(16'h249C,4);
TASK_PP(16'h249D,4);
TASK_PP(16'h249E,4);
TASK_PP(16'h249F,4);
TASK_PP(16'h24A0,4);
TASK_PP(16'h24A1,4);
TASK_PP(16'h24A2,4);
TASK_PP(16'h24A3,4);
TASK_PP(16'h24A4,4);
TASK_PP(16'h24A5,4);
TASK_PP(16'h24A6,4);
TASK_PP(16'h24A7,4);
TASK_PP(16'h24A8,4);
TASK_PP(16'h24A9,4);
TASK_PP(16'h24AA,4);
TASK_PP(16'h24AB,4);
TASK_PP(16'h24AC,4);
TASK_PP(16'h24AD,4);
TASK_PP(16'h24AE,4);
TASK_PP(16'h24AF,4);
TASK_PP(16'h24B0,4);
TASK_PP(16'h24B1,4);
TASK_PP(16'h24B2,4);
TASK_PP(16'h24B3,4);
TASK_PP(16'h24B4,4);
TASK_PP(16'h24B5,4);
TASK_PP(16'h24B6,4);
TASK_PP(16'h24B7,4);
TASK_PP(16'h24B8,4);
TASK_PP(16'h24B9,4);
TASK_PP(16'h24BA,4);
TASK_PP(16'h24BB,4);
TASK_PP(16'h24BC,4);
TASK_PP(16'h24BD,4);
TASK_PP(16'h24BE,4);
TASK_PP(16'h24BF,4);
TASK_PP(16'h24C0,4);
TASK_PP(16'h24C1,4);
TASK_PP(16'h24C2,4);
TASK_PP(16'h24C3,4);
TASK_PP(16'h24C4,4);
TASK_PP(16'h24C5,4);
TASK_PP(16'h24C6,4);
TASK_PP(16'h24C7,4);
TASK_PP(16'h24C8,4);
TASK_PP(16'h24C9,4);
TASK_PP(16'h24CA,4);
TASK_PP(16'h24CB,4);
TASK_PP(16'h24CC,4);
TASK_PP(16'h24CD,4);
TASK_PP(16'h24CE,4);
TASK_PP(16'h24CF,4);
TASK_PP(16'h24D0,4);
TASK_PP(16'h24D1,4);
TASK_PP(16'h24D2,4);
TASK_PP(16'h24D3,4);
TASK_PP(16'h24D4,4);
TASK_PP(16'h24D5,4);
TASK_PP(16'h24D6,4);
TASK_PP(16'h24D7,4);
TASK_PP(16'h24D8,4);
TASK_PP(16'h24D9,4);
TASK_PP(16'h24DA,4);
TASK_PP(16'h24DB,4);
TASK_PP(16'h24DC,4);
TASK_PP(16'h24DD,4);
TASK_PP(16'h24DE,4);
TASK_PP(16'h24DF,4);
TASK_PP(16'h24E0,4);
TASK_PP(16'h24E1,4);
TASK_PP(16'h24E2,4);
TASK_PP(16'h24E3,4);
TASK_PP(16'h24E4,4);
TASK_PP(16'h24E5,4);
TASK_PP(16'h24E6,4);
TASK_PP(16'h24E7,4);
TASK_PP(16'h24E8,4);
TASK_PP(16'h24E9,4);
TASK_PP(16'h24EA,4);
TASK_PP(16'h24EB,4);
TASK_PP(16'h24EC,4);
TASK_PP(16'h24ED,4);
TASK_PP(16'h24EE,4);
TASK_PP(16'h24EF,4);
TASK_PP(16'h24F0,4);
TASK_PP(16'h24F1,4);
TASK_PP(16'h24F2,4);
TASK_PP(16'h24F3,4);
TASK_PP(16'h24F4,4);
TASK_PP(16'h24F5,4);
TASK_PP(16'h24F6,4);
TASK_PP(16'h24F7,4);
TASK_PP(16'h24F8,4);
TASK_PP(16'h24F9,4);
TASK_PP(16'h24FA,4);
TASK_PP(16'h24FB,4);
TASK_PP(16'h24FC,4);
TASK_PP(16'h24FD,4);
TASK_PP(16'h24FE,4);
TASK_PP(16'h24FF,4);
TASK_PP(16'h2500,4);
TASK_PP(16'h2501,4);
TASK_PP(16'h2502,4);
TASK_PP(16'h2503,4);
TASK_PP(16'h2504,4);
TASK_PP(16'h2505,4);
TASK_PP(16'h2506,4);
TASK_PP(16'h2507,4);
TASK_PP(16'h2508,4);
TASK_PP(16'h2509,4);
TASK_PP(16'h250A,4);
TASK_PP(16'h250B,4);
TASK_PP(16'h250C,4);
TASK_PP(16'h250D,4);
TASK_PP(16'h250E,4);
TASK_PP(16'h250F,4);
TASK_PP(16'h2510,4);
TASK_PP(16'h2511,4);
TASK_PP(16'h2512,4);
TASK_PP(16'h2513,4);
TASK_PP(16'h2514,4);
TASK_PP(16'h2515,4);
TASK_PP(16'h2516,4);
TASK_PP(16'h2517,4);
TASK_PP(16'h2518,4);
TASK_PP(16'h2519,4);
TASK_PP(16'h251A,4);
TASK_PP(16'h251B,4);
TASK_PP(16'h251C,4);
TASK_PP(16'h251D,4);
TASK_PP(16'h251E,4);
TASK_PP(16'h251F,4);
TASK_PP(16'h2520,4);
TASK_PP(16'h2521,4);
TASK_PP(16'h2522,4);
TASK_PP(16'h2523,4);
TASK_PP(16'h2524,4);
TASK_PP(16'h2525,4);
TASK_PP(16'h2526,4);
TASK_PP(16'h2527,4);
TASK_PP(16'h2528,4);
TASK_PP(16'h2529,4);
TASK_PP(16'h252A,4);
TASK_PP(16'h252B,4);
TASK_PP(16'h252C,4);
TASK_PP(16'h252D,4);
TASK_PP(16'h252E,4);
TASK_PP(16'h252F,4);
TASK_PP(16'h2530,4);
TASK_PP(16'h2531,4);
TASK_PP(16'h2532,4);
TASK_PP(16'h2533,4);
TASK_PP(16'h2534,4);
TASK_PP(16'h2535,4);
TASK_PP(16'h2536,4);
TASK_PP(16'h2537,4);
TASK_PP(16'h2538,4);
TASK_PP(16'h2539,4);
TASK_PP(16'h253A,4);
TASK_PP(16'h253B,4);
TASK_PP(16'h253C,4);
TASK_PP(16'h253D,4);
TASK_PP(16'h253E,4);
TASK_PP(16'h253F,4);
TASK_PP(16'h2540,4);
TASK_PP(16'h2541,4);
TASK_PP(16'h2542,4);
TASK_PP(16'h2543,4);
TASK_PP(16'h2544,4);
TASK_PP(16'h2545,4);
TASK_PP(16'h2546,4);
TASK_PP(16'h2547,4);
TASK_PP(16'h2548,4);
TASK_PP(16'h2549,4);
TASK_PP(16'h254A,4);
TASK_PP(16'h254B,4);
TASK_PP(16'h254C,4);
TASK_PP(16'h254D,4);
TASK_PP(16'h254E,4);
TASK_PP(16'h254F,4);
TASK_PP(16'h2550,4);
TASK_PP(16'h2551,4);
TASK_PP(16'h2552,4);
TASK_PP(16'h2553,4);
TASK_PP(16'h2554,4);
TASK_PP(16'h2555,4);
TASK_PP(16'h2556,4);
TASK_PP(16'h2557,4);
TASK_PP(16'h2558,4);
TASK_PP(16'h2559,4);
TASK_PP(16'h255A,4);
TASK_PP(16'h255B,4);
TASK_PP(16'h255C,4);
TASK_PP(16'h255D,4);
TASK_PP(16'h255E,4);
TASK_PP(16'h255F,4);
TASK_PP(16'h2560,4);
TASK_PP(16'h2561,4);
TASK_PP(16'h2562,4);
TASK_PP(16'h2563,4);
TASK_PP(16'h2564,4);
TASK_PP(16'h2565,4);
TASK_PP(16'h2566,4);
TASK_PP(16'h2567,4);
TASK_PP(16'h2568,4);
TASK_PP(16'h2569,4);
TASK_PP(16'h256A,4);
TASK_PP(16'h256B,4);
TASK_PP(16'h256C,4);
TASK_PP(16'h256D,4);
TASK_PP(16'h256E,4);
TASK_PP(16'h256F,4);
TASK_PP(16'h2570,4);
TASK_PP(16'h2571,4);
TASK_PP(16'h2572,4);
TASK_PP(16'h2573,4);
TASK_PP(16'h2574,4);
TASK_PP(16'h2575,4);
TASK_PP(16'h2576,4);
TASK_PP(16'h2577,4);
TASK_PP(16'h2578,4);
TASK_PP(16'h2579,4);
TASK_PP(16'h257A,4);
TASK_PP(16'h257B,4);
TASK_PP(16'h257C,4);
TASK_PP(16'h257D,4);
TASK_PP(16'h257E,4);
TASK_PP(16'h257F,4);
TASK_PP(16'h2580,4);
TASK_PP(16'h2581,4);
TASK_PP(16'h2582,4);
TASK_PP(16'h2583,4);
TASK_PP(16'h2584,4);
TASK_PP(16'h2585,4);
TASK_PP(16'h2586,4);
TASK_PP(16'h2587,4);
TASK_PP(16'h2588,4);
TASK_PP(16'h2589,4);
TASK_PP(16'h258A,4);
TASK_PP(16'h258B,4);
TASK_PP(16'h258C,4);
TASK_PP(16'h258D,4);
TASK_PP(16'h258E,4);
TASK_PP(16'h258F,4);
TASK_PP(16'h2590,4);
TASK_PP(16'h2591,4);
TASK_PP(16'h2592,4);
TASK_PP(16'h2593,4);
TASK_PP(16'h2594,4);
TASK_PP(16'h2595,4);
TASK_PP(16'h2596,4);
TASK_PP(16'h2597,4);
TASK_PP(16'h2598,4);
TASK_PP(16'h2599,4);
TASK_PP(16'h259A,4);
TASK_PP(16'h259B,4);
TASK_PP(16'h259C,4);
TASK_PP(16'h259D,4);
TASK_PP(16'h259E,4);
TASK_PP(16'h259F,4);
TASK_PP(16'h25A0,4);
TASK_PP(16'h25A1,4);
TASK_PP(16'h25A2,4);
TASK_PP(16'h25A3,4);
TASK_PP(16'h25A4,4);
TASK_PP(16'h25A5,4);
TASK_PP(16'h25A6,4);
TASK_PP(16'h25A7,4);
TASK_PP(16'h25A8,4);
TASK_PP(16'h25A9,4);
TASK_PP(16'h25AA,4);
TASK_PP(16'h25AB,4);
TASK_PP(16'h25AC,4);
TASK_PP(16'h25AD,4);
TASK_PP(16'h25AE,4);
TASK_PP(16'h25AF,4);
TASK_PP(16'h25B0,4);
TASK_PP(16'h25B1,4);
TASK_PP(16'h25B2,4);
TASK_PP(16'h25B3,4);
TASK_PP(16'h25B4,4);
TASK_PP(16'h25B5,4);
TASK_PP(16'h25B6,4);
TASK_PP(16'h25B7,4);
TASK_PP(16'h25B8,4);
TASK_PP(16'h25B9,4);
TASK_PP(16'h25BA,4);
TASK_PP(16'h25BB,4);
TASK_PP(16'h25BC,4);
TASK_PP(16'h25BD,4);
TASK_PP(16'h25BE,4);
TASK_PP(16'h25BF,4);
TASK_PP(16'h25C0,4);
TASK_PP(16'h25C1,4);
TASK_PP(16'h25C2,4);
TASK_PP(16'h25C3,4);
TASK_PP(16'h25C4,4);
TASK_PP(16'h25C5,4);
TASK_PP(16'h25C6,4);
TASK_PP(16'h25C7,4);
TASK_PP(16'h25C8,4);
TASK_PP(16'h25C9,4);
TASK_PP(16'h25CA,4);
TASK_PP(16'h25CB,4);
TASK_PP(16'h25CC,4);
TASK_PP(16'h25CD,4);
TASK_PP(16'h25CE,4);
TASK_PP(16'h25CF,4);
TASK_PP(16'h25D0,4);
TASK_PP(16'h25D1,4);
TASK_PP(16'h25D2,4);
TASK_PP(16'h25D3,4);
TASK_PP(16'h25D4,4);
TASK_PP(16'h25D5,4);
TASK_PP(16'h25D6,4);
TASK_PP(16'h25D7,4);
TASK_PP(16'h25D8,4);
TASK_PP(16'h25D9,4);
TASK_PP(16'h25DA,4);
TASK_PP(16'h25DB,4);
TASK_PP(16'h25DC,4);
TASK_PP(16'h25DD,4);
TASK_PP(16'h25DE,4);
TASK_PP(16'h25DF,4);
TASK_PP(16'h25E0,4);
TASK_PP(16'h25E1,4);
TASK_PP(16'h25E2,4);
TASK_PP(16'h25E3,4);
TASK_PP(16'h25E4,4);
TASK_PP(16'h25E5,4);
TASK_PP(16'h25E6,4);
TASK_PP(16'h25E7,4);
TASK_PP(16'h25E8,4);
TASK_PP(16'h25E9,4);
TASK_PP(16'h25EA,4);
TASK_PP(16'h25EB,4);
TASK_PP(16'h25EC,4);
TASK_PP(16'h25ED,4);
TASK_PP(16'h25EE,4);
TASK_PP(16'h25EF,4);
TASK_PP(16'h25F0,4);
TASK_PP(16'h25F1,4);
TASK_PP(16'h25F2,4);
TASK_PP(16'h25F3,4);
TASK_PP(16'h25F4,4);
TASK_PP(16'h25F5,4);
TASK_PP(16'h25F6,4);
TASK_PP(16'h25F7,4);
TASK_PP(16'h25F8,4);
TASK_PP(16'h25F9,4);
TASK_PP(16'h25FA,4);
TASK_PP(16'h25FB,4);
TASK_PP(16'h25FC,4);
TASK_PP(16'h25FD,4);
TASK_PP(16'h25FE,4);
TASK_PP(16'h25FF,4);
TASK_PP(16'h2600,4);
TASK_PP(16'h2601,4);
TASK_PP(16'h2602,4);
TASK_PP(16'h2603,4);
TASK_PP(16'h2604,4);
TASK_PP(16'h2605,4);
TASK_PP(16'h2606,4);
TASK_PP(16'h2607,4);
TASK_PP(16'h2608,4);
TASK_PP(16'h2609,4);
TASK_PP(16'h260A,4);
TASK_PP(16'h260B,4);
TASK_PP(16'h260C,4);
TASK_PP(16'h260D,4);
TASK_PP(16'h260E,4);
TASK_PP(16'h260F,4);
TASK_PP(16'h2610,4);
TASK_PP(16'h2611,4);
TASK_PP(16'h2612,4);
TASK_PP(16'h2613,4);
TASK_PP(16'h2614,4);
TASK_PP(16'h2615,4);
TASK_PP(16'h2616,4);
TASK_PP(16'h2617,4);
TASK_PP(16'h2618,4);
TASK_PP(16'h2619,4);
TASK_PP(16'h261A,4);
TASK_PP(16'h261B,4);
TASK_PP(16'h261C,4);
TASK_PP(16'h261D,4);
TASK_PP(16'h261E,4);
TASK_PP(16'h261F,4);
TASK_PP(16'h2620,4);
TASK_PP(16'h2621,4);
TASK_PP(16'h2622,4);
TASK_PP(16'h2623,4);
TASK_PP(16'h2624,4);
TASK_PP(16'h2625,4);
TASK_PP(16'h2626,4);
TASK_PP(16'h2627,4);
TASK_PP(16'h2628,4);
TASK_PP(16'h2629,4);
TASK_PP(16'h262A,4);
TASK_PP(16'h262B,4);
TASK_PP(16'h262C,4);
TASK_PP(16'h262D,4);
TASK_PP(16'h262E,4);
TASK_PP(16'h262F,4);
TASK_PP(16'h2630,4);
TASK_PP(16'h2631,4);
TASK_PP(16'h2632,4);
TASK_PP(16'h2633,4);
TASK_PP(16'h2634,4);
TASK_PP(16'h2635,4);
TASK_PP(16'h2636,4);
TASK_PP(16'h2637,4);
TASK_PP(16'h2638,4);
TASK_PP(16'h2639,4);
TASK_PP(16'h263A,4);
TASK_PP(16'h263B,4);
TASK_PP(16'h263C,4);
TASK_PP(16'h263D,4);
TASK_PP(16'h263E,4);
TASK_PP(16'h263F,4);
TASK_PP(16'h2640,4);
TASK_PP(16'h2641,4);
TASK_PP(16'h2642,4);
TASK_PP(16'h2643,4);
TASK_PP(16'h2644,4);
TASK_PP(16'h2645,4);
TASK_PP(16'h2646,4);
TASK_PP(16'h2647,4);
TASK_PP(16'h2648,4);
TASK_PP(16'h2649,4);
TASK_PP(16'h264A,4);
TASK_PP(16'h264B,4);
TASK_PP(16'h264C,4);
TASK_PP(16'h264D,4);
TASK_PP(16'h264E,4);
TASK_PP(16'h264F,4);
TASK_PP(16'h2650,4);
TASK_PP(16'h2651,4);
TASK_PP(16'h2652,4);
TASK_PP(16'h2653,4);
TASK_PP(16'h2654,4);
TASK_PP(16'h2655,4);
TASK_PP(16'h2656,4);
TASK_PP(16'h2657,4);
TASK_PP(16'h2658,4);
TASK_PP(16'h2659,4);
TASK_PP(16'h265A,4);
TASK_PP(16'h265B,4);
TASK_PP(16'h265C,4);
TASK_PP(16'h265D,4);
TASK_PP(16'h265E,4);
TASK_PP(16'h265F,4);
TASK_PP(16'h2660,4);
TASK_PP(16'h2661,4);
TASK_PP(16'h2662,4);
TASK_PP(16'h2663,4);
TASK_PP(16'h2664,4);
TASK_PP(16'h2665,4);
TASK_PP(16'h2666,4);
TASK_PP(16'h2667,4);
TASK_PP(16'h2668,4);
TASK_PP(16'h2669,4);
TASK_PP(16'h266A,4);
TASK_PP(16'h266B,4);
TASK_PP(16'h266C,4);
TASK_PP(16'h266D,4);
TASK_PP(16'h266E,4);
TASK_PP(16'h266F,4);
TASK_PP(16'h2670,4);
TASK_PP(16'h2671,4);
TASK_PP(16'h2672,4);
TASK_PP(16'h2673,4);
TASK_PP(16'h2674,4);
TASK_PP(16'h2675,4);
TASK_PP(16'h2676,4);
TASK_PP(16'h2677,4);
TASK_PP(16'h2678,4);
TASK_PP(16'h2679,4);
TASK_PP(16'h267A,4);
TASK_PP(16'h267B,4);
TASK_PP(16'h267C,4);
TASK_PP(16'h267D,4);
TASK_PP(16'h267E,4);
TASK_PP(16'h267F,4);
TASK_PP(16'h2680,4);
TASK_PP(16'h2681,4);
TASK_PP(16'h2682,4);
TASK_PP(16'h2683,4);
TASK_PP(16'h2684,4);
TASK_PP(16'h2685,4);
TASK_PP(16'h2686,4);
TASK_PP(16'h2687,4);
TASK_PP(16'h2688,4);
TASK_PP(16'h2689,4);
TASK_PP(16'h268A,4);
TASK_PP(16'h268B,4);
TASK_PP(16'h268C,4);
TASK_PP(16'h268D,4);
TASK_PP(16'h268E,4);
TASK_PP(16'h268F,4);
TASK_PP(16'h2690,4);
TASK_PP(16'h2691,4);
TASK_PP(16'h2692,4);
TASK_PP(16'h2693,4);
TASK_PP(16'h2694,4);
TASK_PP(16'h2695,4);
TASK_PP(16'h2696,4);
TASK_PP(16'h2697,4);
TASK_PP(16'h2698,4);
TASK_PP(16'h2699,4);
TASK_PP(16'h269A,4);
TASK_PP(16'h269B,4);
TASK_PP(16'h269C,4);
TASK_PP(16'h269D,4);
TASK_PP(16'h269E,4);
TASK_PP(16'h269F,4);
TASK_PP(16'h26A0,4);
TASK_PP(16'h26A1,4);
TASK_PP(16'h26A2,4);
TASK_PP(16'h26A3,4);
TASK_PP(16'h26A4,4);
TASK_PP(16'h26A5,4);
TASK_PP(16'h26A6,4);
TASK_PP(16'h26A7,4);
TASK_PP(16'h26A8,4);
TASK_PP(16'h26A9,4);
TASK_PP(16'h26AA,4);
TASK_PP(16'h26AB,4);
TASK_PP(16'h26AC,4);
TASK_PP(16'h26AD,4);
TASK_PP(16'h26AE,4);
TASK_PP(16'h26AF,4);
TASK_PP(16'h26B0,4);
TASK_PP(16'h26B1,4);
TASK_PP(16'h26B2,4);
TASK_PP(16'h26B3,4);
TASK_PP(16'h26B4,4);
TASK_PP(16'h26B5,4);
TASK_PP(16'h26B6,4);
TASK_PP(16'h26B7,4);
TASK_PP(16'h26B8,4);
TASK_PP(16'h26B9,4);
TASK_PP(16'h26BA,4);
TASK_PP(16'h26BB,4);
TASK_PP(16'h26BC,4);
TASK_PP(16'h26BD,4);
TASK_PP(16'h26BE,4);
TASK_PP(16'h26BF,4);
TASK_PP(16'h26C0,4);
TASK_PP(16'h26C1,4);
TASK_PP(16'h26C2,4);
TASK_PP(16'h26C3,4);
TASK_PP(16'h26C4,4);
TASK_PP(16'h26C5,4);
TASK_PP(16'h26C6,4);
TASK_PP(16'h26C7,4);
TASK_PP(16'h26C8,4);
TASK_PP(16'h26C9,4);
TASK_PP(16'h26CA,4);
TASK_PP(16'h26CB,4);
TASK_PP(16'h26CC,4);
TASK_PP(16'h26CD,4);
TASK_PP(16'h26CE,4);
TASK_PP(16'h26CF,4);
TASK_PP(16'h26D0,4);
TASK_PP(16'h26D1,4);
TASK_PP(16'h26D2,4);
TASK_PP(16'h26D3,4);
TASK_PP(16'h26D4,4);
TASK_PP(16'h26D5,4);
TASK_PP(16'h26D6,4);
TASK_PP(16'h26D7,4);
TASK_PP(16'h26D8,4);
TASK_PP(16'h26D9,4);
TASK_PP(16'h26DA,4);
TASK_PP(16'h26DB,4);
TASK_PP(16'h26DC,4);
TASK_PP(16'h26DD,4);
TASK_PP(16'h26DE,4);
TASK_PP(16'h26DF,4);
TASK_PP(16'h26E0,4);
TASK_PP(16'h26E1,4);
TASK_PP(16'h26E2,4);
TASK_PP(16'h26E3,4);
TASK_PP(16'h26E4,4);
TASK_PP(16'h26E5,4);
TASK_PP(16'h26E6,4);
TASK_PP(16'h26E7,4);
TASK_PP(16'h26E8,4);
TASK_PP(16'h26E9,4);
TASK_PP(16'h26EA,4);
TASK_PP(16'h26EB,4);
TASK_PP(16'h26EC,4);
TASK_PP(16'h26ED,4);
TASK_PP(16'h26EE,4);
TASK_PP(16'h26EF,4);
TASK_PP(16'h26F0,4);
TASK_PP(16'h26F1,4);
TASK_PP(16'h26F2,4);
TASK_PP(16'h26F3,4);
TASK_PP(16'h26F4,4);
TASK_PP(16'h26F5,4);
TASK_PP(16'h26F6,4);
TASK_PP(16'h26F7,4);
TASK_PP(16'h26F8,4);
TASK_PP(16'h26F9,4);
TASK_PP(16'h26FA,4);
TASK_PP(16'h26FB,4);
TASK_PP(16'h26FC,4);
TASK_PP(16'h26FD,4);
TASK_PP(16'h26FE,4);
TASK_PP(16'h26FF,4);
TASK_PP(16'h2700,4);
TASK_PP(16'h2701,4);
TASK_PP(16'h2702,4);
TASK_PP(16'h2703,4);
TASK_PP(16'h2704,4);
TASK_PP(16'h2705,4);
TASK_PP(16'h2706,4);
TASK_PP(16'h2707,4);
TASK_PP(16'h2708,4);
TASK_PP(16'h2709,4);
TASK_PP(16'h270A,4);
TASK_PP(16'h270B,4);
TASK_PP(16'h270C,4);
TASK_PP(16'h270D,4);
TASK_PP(16'h270E,4);
TASK_PP(16'h270F,4);
TASK_PP(16'h2710,4);
TASK_PP(16'h2711,4);
TASK_PP(16'h2712,4);
TASK_PP(16'h2713,4);
TASK_PP(16'h2714,4);
TASK_PP(16'h2715,4);
TASK_PP(16'h2716,4);
TASK_PP(16'h2717,4);
TASK_PP(16'h2718,4);
TASK_PP(16'h2719,4);
TASK_PP(16'h271A,4);
TASK_PP(16'h271B,4);
TASK_PP(16'h271C,4);
TASK_PP(16'h271D,4);
TASK_PP(16'h271E,4);
TASK_PP(16'h271F,4);
TASK_PP(16'h2720,4);
TASK_PP(16'h2721,4);
TASK_PP(16'h2722,4);
TASK_PP(16'h2723,4);
TASK_PP(16'h2724,4);
TASK_PP(16'h2725,4);
TASK_PP(16'h2726,4);
TASK_PP(16'h2727,4);
TASK_PP(16'h2728,4);
TASK_PP(16'h2729,4);
TASK_PP(16'h272A,4);
TASK_PP(16'h272B,4);
TASK_PP(16'h272C,4);
TASK_PP(16'h272D,4);
TASK_PP(16'h272E,4);
TASK_PP(16'h272F,4);
TASK_PP(16'h2730,4);
TASK_PP(16'h2731,4);
TASK_PP(16'h2732,4);
TASK_PP(16'h2733,4);
TASK_PP(16'h2734,4);
TASK_PP(16'h2735,4);
TASK_PP(16'h2736,4);
TASK_PP(16'h2737,4);
TASK_PP(16'h2738,4);
TASK_PP(16'h2739,4);
TASK_PP(16'h273A,4);
TASK_PP(16'h273B,4);
TASK_PP(16'h273C,4);
TASK_PP(16'h273D,4);
TASK_PP(16'h273E,4);
TASK_PP(16'h273F,4);
TASK_PP(16'h2740,4);
TASK_PP(16'h2741,4);
TASK_PP(16'h2742,4);
TASK_PP(16'h2743,4);
TASK_PP(16'h2744,4);
TASK_PP(16'h2745,4);
TASK_PP(16'h2746,4);
TASK_PP(16'h2747,4);
TASK_PP(16'h2748,4);
TASK_PP(16'h2749,4);
TASK_PP(16'h274A,4);
TASK_PP(16'h274B,4);
TASK_PP(16'h274C,4);
TASK_PP(16'h274D,4);
TASK_PP(16'h274E,4);
TASK_PP(16'h274F,4);
TASK_PP(16'h2750,4);
TASK_PP(16'h2751,4);
TASK_PP(16'h2752,4);
TASK_PP(16'h2753,4);
TASK_PP(16'h2754,4);
TASK_PP(16'h2755,4);
TASK_PP(16'h2756,4);
TASK_PP(16'h2757,4);
TASK_PP(16'h2758,4);
TASK_PP(16'h2759,4);
TASK_PP(16'h275A,4);
TASK_PP(16'h275B,4);
TASK_PP(16'h275C,4);
TASK_PP(16'h275D,4);
TASK_PP(16'h275E,4);
TASK_PP(16'h275F,4);
TASK_PP(16'h2760,4);
TASK_PP(16'h2761,4);
TASK_PP(16'h2762,4);
TASK_PP(16'h2763,4);
TASK_PP(16'h2764,4);
TASK_PP(16'h2765,4);
TASK_PP(16'h2766,4);
TASK_PP(16'h2767,4);
TASK_PP(16'h2768,4);
TASK_PP(16'h2769,4);
TASK_PP(16'h276A,4);
TASK_PP(16'h276B,4);
TASK_PP(16'h276C,4);
TASK_PP(16'h276D,4);
TASK_PP(16'h276E,4);
TASK_PP(16'h276F,4);
TASK_PP(16'h2770,4);
TASK_PP(16'h2771,4);
TASK_PP(16'h2772,4);
TASK_PP(16'h2773,4);
TASK_PP(16'h2774,4);
TASK_PP(16'h2775,4);
TASK_PP(16'h2776,4);
TASK_PP(16'h2777,4);
TASK_PP(16'h2778,4);
TASK_PP(16'h2779,4);
TASK_PP(16'h277A,4);
TASK_PP(16'h277B,4);
TASK_PP(16'h277C,4);
TASK_PP(16'h277D,4);
TASK_PP(16'h277E,4);
TASK_PP(16'h277F,4);
TASK_PP(16'h2780,4);
TASK_PP(16'h2781,4);
TASK_PP(16'h2782,4);
TASK_PP(16'h2783,4);
TASK_PP(16'h2784,4);
TASK_PP(16'h2785,4);
TASK_PP(16'h2786,4);
TASK_PP(16'h2787,4);
TASK_PP(16'h2788,4);
TASK_PP(16'h2789,4);
TASK_PP(16'h278A,4);
TASK_PP(16'h278B,4);
TASK_PP(16'h278C,4);
TASK_PP(16'h278D,4);
TASK_PP(16'h278E,4);
TASK_PP(16'h278F,4);
TASK_PP(16'h2790,4);
TASK_PP(16'h2791,4);
TASK_PP(16'h2792,4);
TASK_PP(16'h2793,4);
TASK_PP(16'h2794,4);
TASK_PP(16'h2795,4);
TASK_PP(16'h2796,4);
TASK_PP(16'h2797,4);
TASK_PP(16'h2798,4);
TASK_PP(16'h2799,4);
TASK_PP(16'h279A,4);
TASK_PP(16'h279B,4);
TASK_PP(16'h279C,4);
TASK_PP(16'h279D,4);
TASK_PP(16'h279E,4);
TASK_PP(16'h279F,4);
TASK_PP(16'h27A0,4);
TASK_PP(16'h27A1,4);
TASK_PP(16'h27A2,4);
TASK_PP(16'h27A3,4);
TASK_PP(16'h27A4,4);
TASK_PP(16'h27A5,4);
TASK_PP(16'h27A6,4);
TASK_PP(16'h27A7,4);
TASK_PP(16'h27A8,4);
TASK_PP(16'h27A9,4);
TASK_PP(16'h27AA,4);
TASK_PP(16'h27AB,4);
TASK_PP(16'h27AC,4);
TASK_PP(16'h27AD,4);
TASK_PP(16'h27AE,4);
TASK_PP(16'h27AF,4);
TASK_PP(16'h27B0,4);
TASK_PP(16'h27B1,4);
TASK_PP(16'h27B2,4);
TASK_PP(16'h27B3,4);
TASK_PP(16'h27B4,4);
TASK_PP(16'h27B5,4);
TASK_PP(16'h27B6,4);
TASK_PP(16'h27B7,4);
TASK_PP(16'h27B8,4);
TASK_PP(16'h27B9,4);
TASK_PP(16'h27BA,4);
TASK_PP(16'h27BB,4);
TASK_PP(16'h27BC,4);
TASK_PP(16'h27BD,4);
TASK_PP(16'h27BE,4);
TASK_PP(16'h27BF,4);
TASK_PP(16'h27C0,4);
TASK_PP(16'h27C1,4);
TASK_PP(16'h27C2,4);
TASK_PP(16'h27C3,4);
TASK_PP(16'h27C4,4);
TASK_PP(16'h27C5,4);
TASK_PP(16'h27C6,4);
TASK_PP(16'h27C7,4);
TASK_PP(16'h27C8,4);
TASK_PP(16'h27C9,4);
TASK_PP(16'h27CA,4);
TASK_PP(16'h27CB,4);
TASK_PP(16'h27CC,4);
TASK_PP(16'h27CD,4);
TASK_PP(16'h27CE,4);
TASK_PP(16'h27CF,4);
TASK_PP(16'h27D0,4);
TASK_PP(16'h27D1,4);
TASK_PP(16'h27D2,4);
TASK_PP(16'h27D3,4);
TASK_PP(16'h27D4,4);
TASK_PP(16'h27D5,4);
TASK_PP(16'h27D6,4);
TASK_PP(16'h27D7,4);
TASK_PP(16'h27D8,4);
TASK_PP(16'h27D9,4);
TASK_PP(16'h27DA,4);
TASK_PP(16'h27DB,4);
TASK_PP(16'h27DC,4);
TASK_PP(16'h27DD,4);
TASK_PP(16'h27DE,4);
TASK_PP(16'h27DF,4);
TASK_PP(16'h27E0,4);
TASK_PP(16'h27E1,4);
TASK_PP(16'h27E2,4);
TASK_PP(16'h27E3,4);
TASK_PP(16'h27E4,4);
TASK_PP(16'h27E5,4);
TASK_PP(16'h27E6,4);
TASK_PP(16'h27E7,4);
TASK_PP(16'h27E8,4);
TASK_PP(16'h27E9,4);
TASK_PP(16'h27EA,4);
TASK_PP(16'h27EB,4);
TASK_PP(16'h27EC,4);
TASK_PP(16'h27ED,4);
TASK_PP(16'h27EE,4);
TASK_PP(16'h27EF,4);
TASK_PP(16'h27F0,4);
TASK_PP(16'h27F1,4);
TASK_PP(16'h27F2,4);
TASK_PP(16'h27F3,4);
TASK_PP(16'h27F4,4);
TASK_PP(16'h27F5,4);
TASK_PP(16'h27F6,4);
TASK_PP(16'h27F7,4);
TASK_PP(16'h27F8,4);
TASK_PP(16'h27F9,4);
TASK_PP(16'h27FA,4);
TASK_PP(16'h27FB,4);
TASK_PP(16'h27FC,4);
TASK_PP(16'h27FD,4);
TASK_PP(16'h27FE,4);
TASK_PP(16'h27FF,4);
TASK_PP(16'h2800,4);
TASK_PP(16'h2801,4);
TASK_PP(16'h2802,4);
TASK_PP(16'h2803,4);
TASK_PP(16'h2804,4);
TASK_PP(16'h2805,4);
TASK_PP(16'h2806,4);
TASK_PP(16'h2807,4);
TASK_PP(16'h2808,4);
TASK_PP(16'h2809,4);
TASK_PP(16'h280A,4);
TASK_PP(16'h280B,4);
TASK_PP(16'h280C,4);
TASK_PP(16'h280D,4);
TASK_PP(16'h280E,4);
TASK_PP(16'h280F,4);
TASK_PP(16'h2810,4);
TASK_PP(16'h2811,4);
TASK_PP(16'h2812,4);
TASK_PP(16'h2813,4);
TASK_PP(16'h2814,4);
TASK_PP(16'h2815,4);
TASK_PP(16'h2816,4);
TASK_PP(16'h2817,4);
TASK_PP(16'h2818,4);
TASK_PP(16'h2819,4);
TASK_PP(16'h281A,4);
TASK_PP(16'h281B,4);
TASK_PP(16'h281C,4);
TASK_PP(16'h281D,4);
TASK_PP(16'h281E,4);
TASK_PP(16'h281F,4);
TASK_PP(16'h2820,4);
TASK_PP(16'h2821,4);
TASK_PP(16'h2822,4);
TASK_PP(16'h2823,4);
TASK_PP(16'h2824,4);
TASK_PP(16'h2825,4);
TASK_PP(16'h2826,4);
TASK_PP(16'h2827,4);
TASK_PP(16'h2828,4);
TASK_PP(16'h2829,4);
TASK_PP(16'h282A,4);
TASK_PP(16'h282B,4);
TASK_PP(16'h282C,4);
TASK_PP(16'h282D,4);
TASK_PP(16'h282E,4);
TASK_PP(16'h282F,4);
TASK_PP(16'h2830,4);
TASK_PP(16'h2831,4);
TASK_PP(16'h2832,4);
TASK_PP(16'h2833,4);
TASK_PP(16'h2834,4);
TASK_PP(16'h2835,4);
TASK_PP(16'h2836,4);
TASK_PP(16'h2837,4);
TASK_PP(16'h2838,4);
TASK_PP(16'h2839,4);
TASK_PP(16'h283A,4);
TASK_PP(16'h283B,4);
TASK_PP(16'h283C,4);
TASK_PP(16'h283D,4);
TASK_PP(16'h283E,4);
TASK_PP(16'h283F,4);
TASK_PP(16'h2840,4);
TASK_PP(16'h2841,4);
TASK_PP(16'h2842,4);
TASK_PP(16'h2843,4);
TASK_PP(16'h2844,4);
TASK_PP(16'h2845,4);
TASK_PP(16'h2846,4);
TASK_PP(16'h2847,4);
TASK_PP(16'h2848,4);
TASK_PP(16'h2849,4);
TASK_PP(16'h284A,4);
TASK_PP(16'h284B,4);
TASK_PP(16'h284C,4);
TASK_PP(16'h284D,4);
TASK_PP(16'h284E,4);
TASK_PP(16'h284F,4);
TASK_PP(16'h2850,4);
TASK_PP(16'h2851,4);
TASK_PP(16'h2852,4);
TASK_PP(16'h2853,4);
TASK_PP(16'h2854,4);
TASK_PP(16'h2855,4);
TASK_PP(16'h2856,4);
TASK_PP(16'h2857,4);
TASK_PP(16'h2858,4);
TASK_PP(16'h2859,4);
TASK_PP(16'h285A,4);
TASK_PP(16'h285B,4);
TASK_PP(16'h285C,4);
TASK_PP(16'h285D,4);
TASK_PP(16'h285E,4);
TASK_PP(16'h285F,4);
TASK_PP(16'h2860,4);
TASK_PP(16'h2861,4);
TASK_PP(16'h2862,4);
TASK_PP(16'h2863,4);
TASK_PP(16'h2864,4);
TASK_PP(16'h2865,4);
TASK_PP(16'h2866,4);
TASK_PP(16'h2867,4);
TASK_PP(16'h2868,4);
TASK_PP(16'h2869,4);
TASK_PP(16'h286A,4);
TASK_PP(16'h286B,4);
TASK_PP(16'h286C,4);
TASK_PP(16'h286D,4);
TASK_PP(16'h286E,4);
TASK_PP(16'h286F,4);
TASK_PP(16'h2870,4);
TASK_PP(16'h2871,4);
TASK_PP(16'h2872,4);
TASK_PP(16'h2873,4);
TASK_PP(16'h2874,4);
TASK_PP(16'h2875,4);
TASK_PP(16'h2876,4);
TASK_PP(16'h2877,4);
TASK_PP(16'h2878,4);
TASK_PP(16'h2879,4);
TASK_PP(16'h287A,4);
TASK_PP(16'h287B,4);
TASK_PP(16'h287C,4);
TASK_PP(16'h287D,4);
TASK_PP(16'h287E,4);
TASK_PP(16'h287F,4);
TASK_PP(16'h2880,4);
TASK_PP(16'h2881,4);
TASK_PP(16'h2882,4);
TASK_PP(16'h2883,4);
TASK_PP(16'h2884,4);
TASK_PP(16'h2885,4);
TASK_PP(16'h2886,4);
TASK_PP(16'h2887,4);
TASK_PP(16'h2888,4);
TASK_PP(16'h2889,4);
TASK_PP(16'h288A,4);
TASK_PP(16'h288B,4);
TASK_PP(16'h288C,4);
TASK_PP(16'h288D,4);
TASK_PP(16'h288E,4);
TASK_PP(16'h288F,4);
TASK_PP(16'h2890,4);
TASK_PP(16'h2891,4);
TASK_PP(16'h2892,4);
TASK_PP(16'h2893,4);
TASK_PP(16'h2894,4);
TASK_PP(16'h2895,4);
TASK_PP(16'h2896,4);
TASK_PP(16'h2897,4);
TASK_PP(16'h2898,4);
TASK_PP(16'h2899,4);
TASK_PP(16'h289A,4);
TASK_PP(16'h289B,4);
TASK_PP(16'h289C,4);
TASK_PP(16'h289D,4);
TASK_PP(16'h289E,4);
TASK_PP(16'h289F,4);
TASK_PP(16'h28A0,4);
TASK_PP(16'h28A1,4);
TASK_PP(16'h28A2,4);
TASK_PP(16'h28A3,4);
TASK_PP(16'h28A4,4);
TASK_PP(16'h28A5,4);
TASK_PP(16'h28A6,4);
TASK_PP(16'h28A7,4);
TASK_PP(16'h28A8,4);
TASK_PP(16'h28A9,4);
TASK_PP(16'h28AA,4);
TASK_PP(16'h28AB,4);
TASK_PP(16'h28AC,4);
TASK_PP(16'h28AD,4);
TASK_PP(16'h28AE,4);
TASK_PP(16'h28AF,4);
TASK_PP(16'h28B0,4);
TASK_PP(16'h28B1,4);
TASK_PP(16'h28B2,4);
TASK_PP(16'h28B3,4);
TASK_PP(16'h28B4,4);
TASK_PP(16'h28B5,4);
TASK_PP(16'h28B6,4);
TASK_PP(16'h28B7,4);
TASK_PP(16'h28B8,4);
TASK_PP(16'h28B9,4);
TASK_PP(16'h28BA,4);
TASK_PP(16'h28BB,4);
TASK_PP(16'h28BC,4);
TASK_PP(16'h28BD,4);
TASK_PP(16'h28BE,4);
TASK_PP(16'h28BF,4);
TASK_PP(16'h28C0,4);
TASK_PP(16'h28C1,4);
TASK_PP(16'h28C2,4);
TASK_PP(16'h28C3,4);
TASK_PP(16'h28C4,4);
TASK_PP(16'h28C5,4);
TASK_PP(16'h28C6,4);
TASK_PP(16'h28C7,4);
TASK_PP(16'h28C8,4);
TASK_PP(16'h28C9,4);
TASK_PP(16'h28CA,4);
TASK_PP(16'h28CB,4);
TASK_PP(16'h28CC,4);
TASK_PP(16'h28CD,4);
TASK_PP(16'h28CE,4);
TASK_PP(16'h28CF,4);
TASK_PP(16'h28D0,4);
TASK_PP(16'h28D1,4);
TASK_PP(16'h28D2,4);
TASK_PP(16'h28D3,4);
TASK_PP(16'h28D4,4);
TASK_PP(16'h28D5,4);
TASK_PP(16'h28D6,4);
TASK_PP(16'h28D7,4);
TASK_PP(16'h28D8,4);
TASK_PP(16'h28D9,4);
TASK_PP(16'h28DA,4);
TASK_PP(16'h28DB,4);
TASK_PP(16'h28DC,4);
TASK_PP(16'h28DD,4);
TASK_PP(16'h28DE,4);
TASK_PP(16'h28DF,4);
TASK_PP(16'h28E0,4);
TASK_PP(16'h28E1,4);
TASK_PP(16'h28E2,4);
TASK_PP(16'h28E3,4);
TASK_PP(16'h28E4,4);
TASK_PP(16'h28E5,4);
TASK_PP(16'h28E6,4);
TASK_PP(16'h28E7,4);
TASK_PP(16'h28E8,4);
TASK_PP(16'h28E9,4);
TASK_PP(16'h28EA,4);
TASK_PP(16'h28EB,4);
TASK_PP(16'h28EC,4);
TASK_PP(16'h28ED,4);
TASK_PP(16'h28EE,4);
TASK_PP(16'h28EF,4);
TASK_PP(16'h28F0,4);
TASK_PP(16'h28F1,4);
TASK_PP(16'h28F2,4);
TASK_PP(16'h28F3,4);
TASK_PP(16'h28F4,4);
TASK_PP(16'h28F5,4);
TASK_PP(16'h28F6,4);
TASK_PP(16'h28F7,4);
TASK_PP(16'h28F8,4);
TASK_PP(16'h28F9,4);
TASK_PP(16'h28FA,4);
TASK_PP(16'h28FB,4);
TASK_PP(16'h28FC,4);
TASK_PP(16'h28FD,4);
TASK_PP(16'h28FE,4);
TASK_PP(16'h28FF,4);
TASK_PP(16'h2900,4);
TASK_PP(16'h2901,4);
TASK_PP(16'h2902,4);
TASK_PP(16'h2903,4);
TASK_PP(16'h2904,4);
TASK_PP(16'h2905,4);
TASK_PP(16'h2906,4);
TASK_PP(16'h2907,4);
TASK_PP(16'h2908,4);
TASK_PP(16'h2909,4);
TASK_PP(16'h290A,4);
TASK_PP(16'h290B,4);
TASK_PP(16'h290C,4);
TASK_PP(16'h290D,4);
TASK_PP(16'h290E,4);
TASK_PP(16'h290F,4);
TASK_PP(16'h2910,4);
TASK_PP(16'h2911,4);
TASK_PP(16'h2912,4);
TASK_PP(16'h2913,4);
TASK_PP(16'h2914,4);
TASK_PP(16'h2915,4);
TASK_PP(16'h2916,4);
TASK_PP(16'h2917,4);
TASK_PP(16'h2918,4);
TASK_PP(16'h2919,4);
TASK_PP(16'h291A,4);
TASK_PP(16'h291B,4);
TASK_PP(16'h291C,4);
TASK_PP(16'h291D,4);
TASK_PP(16'h291E,4);
TASK_PP(16'h291F,4);
TASK_PP(16'h2920,4);
TASK_PP(16'h2921,4);
TASK_PP(16'h2922,4);
TASK_PP(16'h2923,4);
TASK_PP(16'h2924,4);
TASK_PP(16'h2925,4);
TASK_PP(16'h2926,4);
TASK_PP(16'h2927,4);
TASK_PP(16'h2928,4);
TASK_PP(16'h2929,4);
TASK_PP(16'h292A,4);
TASK_PP(16'h292B,4);
TASK_PP(16'h292C,4);
TASK_PP(16'h292D,4);
TASK_PP(16'h292E,4);
TASK_PP(16'h292F,4);
TASK_PP(16'h2930,4);
TASK_PP(16'h2931,4);
TASK_PP(16'h2932,4);
TASK_PP(16'h2933,4);
TASK_PP(16'h2934,4);
TASK_PP(16'h2935,4);
TASK_PP(16'h2936,4);
TASK_PP(16'h2937,4);
TASK_PP(16'h2938,4);
TASK_PP(16'h2939,4);
TASK_PP(16'h293A,4);
TASK_PP(16'h293B,4);
TASK_PP(16'h293C,4);
TASK_PP(16'h293D,4);
TASK_PP(16'h293E,4);
TASK_PP(16'h293F,4);
TASK_PP(16'h2940,4);
TASK_PP(16'h2941,4);
TASK_PP(16'h2942,4);
TASK_PP(16'h2943,4);
TASK_PP(16'h2944,4);
TASK_PP(16'h2945,4);
TASK_PP(16'h2946,4);
TASK_PP(16'h2947,4);
TASK_PP(16'h2948,4);
TASK_PP(16'h2949,4);
TASK_PP(16'h294A,4);
TASK_PP(16'h294B,4);
TASK_PP(16'h294C,4);
TASK_PP(16'h294D,4);
TASK_PP(16'h294E,4);
TASK_PP(16'h294F,4);
TASK_PP(16'h2950,4);
TASK_PP(16'h2951,4);
TASK_PP(16'h2952,4);
TASK_PP(16'h2953,4);
TASK_PP(16'h2954,4);
TASK_PP(16'h2955,4);
TASK_PP(16'h2956,4);
TASK_PP(16'h2957,4);
TASK_PP(16'h2958,4);
TASK_PP(16'h2959,4);
TASK_PP(16'h295A,4);
TASK_PP(16'h295B,4);
TASK_PP(16'h295C,4);
TASK_PP(16'h295D,4);
TASK_PP(16'h295E,4);
TASK_PP(16'h295F,4);
TASK_PP(16'h2960,4);
TASK_PP(16'h2961,4);
TASK_PP(16'h2962,4);
TASK_PP(16'h2963,4);
TASK_PP(16'h2964,4);
TASK_PP(16'h2965,4);
TASK_PP(16'h2966,4);
TASK_PP(16'h2967,4);
TASK_PP(16'h2968,4);
TASK_PP(16'h2969,4);
TASK_PP(16'h296A,4);
TASK_PP(16'h296B,4);
TASK_PP(16'h296C,4);
TASK_PP(16'h296D,4);
TASK_PP(16'h296E,4);
TASK_PP(16'h296F,4);
TASK_PP(16'h2970,4);
TASK_PP(16'h2971,4);
TASK_PP(16'h2972,4);
TASK_PP(16'h2973,4);
TASK_PP(16'h2974,4);
TASK_PP(16'h2975,4);
TASK_PP(16'h2976,4);
TASK_PP(16'h2977,4);
TASK_PP(16'h2978,4);
TASK_PP(16'h2979,4);
TASK_PP(16'h297A,4);
TASK_PP(16'h297B,4);
TASK_PP(16'h297C,4);
TASK_PP(16'h297D,4);
TASK_PP(16'h297E,4);
TASK_PP(16'h297F,4);
TASK_PP(16'h2980,4);
TASK_PP(16'h2981,4);
TASK_PP(16'h2982,4);
TASK_PP(16'h2983,4);
TASK_PP(16'h2984,4);
TASK_PP(16'h2985,4);
TASK_PP(16'h2986,4);
TASK_PP(16'h2987,4);
TASK_PP(16'h2988,4);
TASK_PP(16'h2989,4);
TASK_PP(16'h298A,4);
TASK_PP(16'h298B,4);
TASK_PP(16'h298C,4);
TASK_PP(16'h298D,4);
TASK_PP(16'h298E,4);
TASK_PP(16'h298F,4);
TASK_PP(16'h2990,4);
TASK_PP(16'h2991,4);
TASK_PP(16'h2992,4);
TASK_PP(16'h2993,4);
TASK_PP(16'h2994,4);
TASK_PP(16'h2995,4);
TASK_PP(16'h2996,4);
TASK_PP(16'h2997,4);
TASK_PP(16'h2998,4);
TASK_PP(16'h2999,4);
TASK_PP(16'h299A,4);
TASK_PP(16'h299B,4);
TASK_PP(16'h299C,4);
TASK_PP(16'h299D,4);
TASK_PP(16'h299E,4);
TASK_PP(16'h299F,4);
TASK_PP(16'h29A0,4);
TASK_PP(16'h29A1,4);
TASK_PP(16'h29A2,4);
TASK_PP(16'h29A3,4);
TASK_PP(16'h29A4,4);
TASK_PP(16'h29A5,4);
TASK_PP(16'h29A6,4);
TASK_PP(16'h29A7,4);
TASK_PP(16'h29A8,4);
TASK_PP(16'h29A9,4);
TASK_PP(16'h29AA,4);
TASK_PP(16'h29AB,4);
TASK_PP(16'h29AC,4);
TASK_PP(16'h29AD,4);
TASK_PP(16'h29AE,4);
TASK_PP(16'h29AF,4);
TASK_PP(16'h29B0,4);
TASK_PP(16'h29B1,4);
TASK_PP(16'h29B2,4);
TASK_PP(16'h29B3,4);
TASK_PP(16'h29B4,4);
TASK_PP(16'h29B5,4);
TASK_PP(16'h29B6,4);
TASK_PP(16'h29B7,4);
TASK_PP(16'h29B8,4);
TASK_PP(16'h29B9,4);
TASK_PP(16'h29BA,4);
TASK_PP(16'h29BB,4);
TASK_PP(16'h29BC,4);
TASK_PP(16'h29BD,4);
TASK_PP(16'h29BE,4);
TASK_PP(16'h29BF,4);
TASK_PP(16'h29C0,4);
TASK_PP(16'h29C1,4);
TASK_PP(16'h29C2,4);
TASK_PP(16'h29C3,4);
TASK_PP(16'h29C4,4);
TASK_PP(16'h29C5,4);
TASK_PP(16'h29C6,4);
TASK_PP(16'h29C7,4);
TASK_PP(16'h29C8,4);
TASK_PP(16'h29C9,4);
TASK_PP(16'h29CA,4);
TASK_PP(16'h29CB,4);
TASK_PP(16'h29CC,4);
TASK_PP(16'h29CD,4);
TASK_PP(16'h29CE,4);
TASK_PP(16'h29CF,4);
TASK_PP(16'h29D0,4);
TASK_PP(16'h29D1,4);
TASK_PP(16'h29D2,4);
TASK_PP(16'h29D3,4);
TASK_PP(16'h29D4,4);
TASK_PP(16'h29D5,4);
TASK_PP(16'h29D6,4);
TASK_PP(16'h29D7,4);
TASK_PP(16'h29D8,4);
TASK_PP(16'h29D9,4);
TASK_PP(16'h29DA,4);
TASK_PP(16'h29DB,4);
TASK_PP(16'h29DC,4);
TASK_PP(16'h29DD,4);
TASK_PP(16'h29DE,4);
TASK_PP(16'h29DF,4);
TASK_PP(16'h29E0,4);
TASK_PP(16'h29E1,4);
TASK_PP(16'h29E2,4);
TASK_PP(16'h29E3,4);
TASK_PP(16'h29E4,4);
TASK_PP(16'h29E5,4);
TASK_PP(16'h29E6,4);
TASK_PP(16'h29E7,4);
TASK_PP(16'h29E8,4);
TASK_PP(16'h29E9,4);
TASK_PP(16'h29EA,4);
TASK_PP(16'h29EB,4);
TASK_PP(16'h29EC,4);
TASK_PP(16'h29ED,4);
TASK_PP(16'h29EE,4);
TASK_PP(16'h29EF,4);
TASK_PP(16'h29F0,4);
TASK_PP(16'h29F1,4);
TASK_PP(16'h29F2,4);
TASK_PP(16'h29F3,4);
TASK_PP(16'h29F4,4);
TASK_PP(16'h29F5,4);
TASK_PP(16'h29F6,4);
TASK_PP(16'h29F7,4);
TASK_PP(16'h29F8,4);
TASK_PP(16'h29F9,4);
TASK_PP(16'h29FA,4);
TASK_PP(16'h29FB,4);
TASK_PP(16'h29FC,4);
TASK_PP(16'h29FD,4);
TASK_PP(16'h29FE,4);
TASK_PP(16'h29FF,4);
TASK_PP(16'h2A00,4);
TASK_PP(16'h2A01,4);
TASK_PP(16'h2A02,4);
TASK_PP(16'h2A03,4);
TASK_PP(16'h2A04,4);
TASK_PP(16'h2A05,4);
TASK_PP(16'h2A06,4);
TASK_PP(16'h2A07,4);
TASK_PP(16'h2A08,4);
TASK_PP(16'h2A09,4);
TASK_PP(16'h2A0A,4);
TASK_PP(16'h2A0B,4);
TASK_PP(16'h2A0C,4);
TASK_PP(16'h2A0D,4);
TASK_PP(16'h2A0E,4);
TASK_PP(16'h2A0F,4);
TASK_PP(16'h2A10,4);
TASK_PP(16'h2A11,4);
TASK_PP(16'h2A12,4);
TASK_PP(16'h2A13,4);
TASK_PP(16'h2A14,4);
TASK_PP(16'h2A15,4);
TASK_PP(16'h2A16,4);
TASK_PP(16'h2A17,4);
TASK_PP(16'h2A18,4);
TASK_PP(16'h2A19,4);
TASK_PP(16'h2A1A,4);
TASK_PP(16'h2A1B,4);
TASK_PP(16'h2A1C,4);
TASK_PP(16'h2A1D,4);
TASK_PP(16'h2A1E,4);
TASK_PP(16'h2A1F,4);
TASK_PP(16'h2A20,4);
TASK_PP(16'h2A21,4);
TASK_PP(16'h2A22,4);
TASK_PP(16'h2A23,4);
TASK_PP(16'h2A24,4);
TASK_PP(16'h2A25,4);
TASK_PP(16'h2A26,4);
TASK_PP(16'h2A27,4);
TASK_PP(16'h2A28,4);
TASK_PP(16'h2A29,4);
TASK_PP(16'h2A2A,4);
TASK_PP(16'h2A2B,4);
TASK_PP(16'h2A2C,4);
TASK_PP(16'h2A2D,4);
TASK_PP(16'h2A2E,4);
TASK_PP(16'h2A2F,4);
TASK_PP(16'h2A30,4);
TASK_PP(16'h2A31,4);
TASK_PP(16'h2A32,4);
TASK_PP(16'h2A33,4);
TASK_PP(16'h2A34,4);
TASK_PP(16'h2A35,4);
TASK_PP(16'h2A36,4);
TASK_PP(16'h2A37,4);
TASK_PP(16'h2A38,4);
TASK_PP(16'h2A39,4);
TASK_PP(16'h2A3A,4);
TASK_PP(16'h2A3B,4);
TASK_PP(16'h2A3C,4);
TASK_PP(16'h2A3D,4);
TASK_PP(16'h2A3E,4);
TASK_PP(16'h2A3F,4);
TASK_PP(16'h2A40,4);
TASK_PP(16'h2A41,4);
TASK_PP(16'h2A42,4);
TASK_PP(16'h2A43,4);
TASK_PP(16'h2A44,4);
TASK_PP(16'h2A45,4);
TASK_PP(16'h2A46,4);
TASK_PP(16'h2A47,4);
TASK_PP(16'h2A48,4);
TASK_PP(16'h2A49,4);
TASK_PP(16'h2A4A,4);
TASK_PP(16'h2A4B,4);
TASK_PP(16'h2A4C,4);
TASK_PP(16'h2A4D,4);
TASK_PP(16'h2A4E,4);
TASK_PP(16'h2A4F,4);
TASK_PP(16'h2A50,4);
TASK_PP(16'h2A51,4);
TASK_PP(16'h2A52,4);
TASK_PP(16'h2A53,4);
TASK_PP(16'h2A54,4);
TASK_PP(16'h2A55,4);
TASK_PP(16'h2A56,4);
TASK_PP(16'h2A57,4);
TASK_PP(16'h2A58,4);
TASK_PP(16'h2A59,4);
TASK_PP(16'h2A5A,4);
TASK_PP(16'h2A5B,4);
TASK_PP(16'h2A5C,4);
TASK_PP(16'h2A5D,4);
TASK_PP(16'h2A5E,4);
TASK_PP(16'h2A5F,4);
TASK_PP(16'h2A60,4);
TASK_PP(16'h2A61,4);
TASK_PP(16'h2A62,4);
TASK_PP(16'h2A63,4);
TASK_PP(16'h2A64,4);
TASK_PP(16'h2A65,4);
TASK_PP(16'h2A66,4);
TASK_PP(16'h2A67,4);
TASK_PP(16'h2A68,4);
TASK_PP(16'h2A69,4);
TASK_PP(16'h2A6A,4);
TASK_PP(16'h2A6B,4);
TASK_PP(16'h2A6C,4);
TASK_PP(16'h2A6D,4);
TASK_PP(16'h2A6E,4);
TASK_PP(16'h2A6F,4);
TASK_PP(16'h2A70,4);
TASK_PP(16'h2A71,4);
TASK_PP(16'h2A72,4);
TASK_PP(16'h2A73,4);
TASK_PP(16'h2A74,4);
TASK_PP(16'h2A75,4);
TASK_PP(16'h2A76,4);
TASK_PP(16'h2A77,4);
TASK_PP(16'h2A78,4);
TASK_PP(16'h2A79,4);
TASK_PP(16'h2A7A,4);
TASK_PP(16'h2A7B,4);
TASK_PP(16'h2A7C,4);
TASK_PP(16'h2A7D,4);
TASK_PP(16'h2A7E,4);
TASK_PP(16'h2A7F,4);
TASK_PP(16'h2A80,4);
TASK_PP(16'h2A81,4);
TASK_PP(16'h2A82,4);
TASK_PP(16'h2A83,4);
TASK_PP(16'h2A84,4);
TASK_PP(16'h2A85,4);
TASK_PP(16'h2A86,4);
TASK_PP(16'h2A87,4);
TASK_PP(16'h2A88,4);
TASK_PP(16'h2A89,4);
TASK_PP(16'h2A8A,4);
TASK_PP(16'h2A8B,4);
TASK_PP(16'h2A8C,4);
TASK_PP(16'h2A8D,4);
TASK_PP(16'h2A8E,4);
TASK_PP(16'h2A8F,4);
TASK_PP(16'h2A90,4);
TASK_PP(16'h2A91,4);
TASK_PP(16'h2A92,4);
TASK_PP(16'h2A93,4);
TASK_PP(16'h2A94,4);
TASK_PP(16'h2A95,4);
TASK_PP(16'h2A96,4);
TASK_PP(16'h2A97,4);
TASK_PP(16'h2A98,4);
TASK_PP(16'h2A99,4);
TASK_PP(16'h2A9A,4);
TASK_PP(16'h2A9B,4);
TASK_PP(16'h2A9C,4);
TASK_PP(16'h2A9D,4);
TASK_PP(16'h2A9E,4);
TASK_PP(16'h2A9F,4);
TASK_PP(16'h2AA0,4);
TASK_PP(16'h2AA1,4);
TASK_PP(16'h2AA2,4);
TASK_PP(16'h2AA3,4);
TASK_PP(16'h2AA4,4);
TASK_PP(16'h2AA5,4);
TASK_PP(16'h2AA6,4);
TASK_PP(16'h2AA7,4);
TASK_PP(16'h2AA8,4);
TASK_PP(16'h2AA9,4);
TASK_PP(16'h2AAA,4);
TASK_PP(16'h2AAB,4);
TASK_PP(16'h2AAC,4);
TASK_PP(16'h2AAD,4);
TASK_PP(16'h2AAE,4);
TASK_PP(16'h2AAF,4);
TASK_PP(16'h2AB0,4);
TASK_PP(16'h2AB1,4);
TASK_PP(16'h2AB2,4);
TASK_PP(16'h2AB3,4);
TASK_PP(16'h2AB4,4);
TASK_PP(16'h2AB5,4);
TASK_PP(16'h2AB6,4);
TASK_PP(16'h2AB7,4);
TASK_PP(16'h2AB8,4);
TASK_PP(16'h2AB9,4);
TASK_PP(16'h2ABA,4);
TASK_PP(16'h2ABB,4);
TASK_PP(16'h2ABC,4);
TASK_PP(16'h2ABD,4);
TASK_PP(16'h2ABE,4);
TASK_PP(16'h2ABF,4);
TASK_PP(16'h2AC0,4);
TASK_PP(16'h2AC1,4);
TASK_PP(16'h2AC2,4);
TASK_PP(16'h2AC3,4);
TASK_PP(16'h2AC4,4);
TASK_PP(16'h2AC5,4);
TASK_PP(16'h2AC6,4);
TASK_PP(16'h2AC7,4);
TASK_PP(16'h2AC8,4);
TASK_PP(16'h2AC9,4);
TASK_PP(16'h2ACA,4);
TASK_PP(16'h2ACB,4);
TASK_PP(16'h2ACC,4);
TASK_PP(16'h2ACD,4);
TASK_PP(16'h2ACE,4);
TASK_PP(16'h2ACF,4);
TASK_PP(16'h2AD0,4);
TASK_PP(16'h2AD1,4);
TASK_PP(16'h2AD2,4);
TASK_PP(16'h2AD3,4);
TASK_PP(16'h2AD4,4);
TASK_PP(16'h2AD5,4);
TASK_PP(16'h2AD6,4);
TASK_PP(16'h2AD7,4);
TASK_PP(16'h2AD8,4);
TASK_PP(16'h2AD9,4);
TASK_PP(16'h2ADA,4);
TASK_PP(16'h2ADB,4);
TASK_PP(16'h2ADC,4);
TASK_PP(16'h2ADD,4);
TASK_PP(16'h2ADE,4);
TASK_PP(16'h2ADF,4);
TASK_PP(16'h2AE0,4);
TASK_PP(16'h2AE1,4);
TASK_PP(16'h2AE2,4);
TASK_PP(16'h2AE3,4);
TASK_PP(16'h2AE4,4);
TASK_PP(16'h2AE5,4);
TASK_PP(16'h2AE6,4);
TASK_PP(16'h2AE7,4);
TASK_PP(16'h2AE8,4);
TASK_PP(16'h2AE9,4);
TASK_PP(16'h2AEA,4);
TASK_PP(16'h2AEB,4);
TASK_PP(16'h2AEC,4);
TASK_PP(16'h2AED,4);
TASK_PP(16'h2AEE,4);
TASK_PP(16'h2AEF,4);
TASK_PP(16'h2AF0,4);
TASK_PP(16'h2AF1,4);
TASK_PP(16'h2AF2,4);
TASK_PP(16'h2AF3,4);
TASK_PP(16'h2AF4,4);
TASK_PP(16'h2AF5,4);
TASK_PP(16'h2AF6,4);
TASK_PP(16'h2AF7,4);
TASK_PP(16'h2AF8,4);
TASK_PP(16'h2AF9,4);
TASK_PP(16'h2AFA,4);
TASK_PP(16'h2AFB,4);
TASK_PP(16'h2AFC,4);
TASK_PP(16'h2AFD,4);
TASK_PP(16'h2AFE,4);
TASK_PP(16'h2AFF,4);
TASK_PP(16'h2B00,4);
TASK_PP(16'h2B01,4);
TASK_PP(16'h2B02,4);
TASK_PP(16'h2B03,4);
TASK_PP(16'h2B04,4);
TASK_PP(16'h2B05,4);
TASK_PP(16'h2B06,4);
TASK_PP(16'h2B07,4);
TASK_PP(16'h2B08,4);
TASK_PP(16'h2B09,4);
TASK_PP(16'h2B0A,4);
TASK_PP(16'h2B0B,4);
TASK_PP(16'h2B0C,4);
TASK_PP(16'h2B0D,4);
TASK_PP(16'h2B0E,4);
TASK_PP(16'h2B0F,4);
TASK_PP(16'h2B10,4);
TASK_PP(16'h2B11,4);
TASK_PP(16'h2B12,4);
TASK_PP(16'h2B13,4);
TASK_PP(16'h2B14,4);
TASK_PP(16'h2B15,4);
TASK_PP(16'h2B16,4);
TASK_PP(16'h2B17,4);
TASK_PP(16'h2B18,4);
TASK_PP(16'h2B19,4);
TASK_PP(16'h2B1A,4);
TASK_PP(16'h2B1B,4);
TASK_PP(16'h2B1C,4);
TASK_PP(16'h2B1D,4);
TASK_PP(16'h2B1E,4);
TASK_PP(16'h2B1F,4);
TASK_PP(16'h2B20,4);
TASK_PP(16'h2B21,4);
TASK_PP(16'h2B22,4);
TASK_PP(16'h2B23,4);
TASK_PP(16'h2B24,4);
TASK_PP(16'h2B25,4);
TASK_PP(16'h2B26,4);
TASK_PP(16'h2B27,4);
TASK_PP(16'h2B28,4);
TASK_PP(16'h2B29,4);
TASK_PP(16'h2B2A,4);
TASK_PP(16'h2B2B,4);
TASK_PP(16'h2B2C,4);
TASK_PP(16'h2B2D,4);
TASK_PP(16'h2B2E,4);
TASK_PP(16'h2B2F,4);
TASK_PP(16'h2B30,4);
TASK_PP(16'h2B31,4);
TASK_PP(16'h2B32,4);
TASK_PP(16'h2B33,4);
TASK_PP(16'h2B34,4);
TASK_PP(16'h2B35,4);
TASK_PP(16'h2B36,4);
TASK_PP(16'h2B37,4);
TASK_PP(16'h2B38,4);
TASK_PP(16'h2B39,4);
TASK_PP(16'h2B3A,4);
TASK_PP(16'h2B3B,4);
TASK_PP(16'h2B3C,4);
TASK_PP(16'h2B3D,4);
TASK_PP(16'h2B3E,4);
TASK_PP(16'h2B3F,4);
TASK_PP(16'h2B40,4);
TASK_PP(16'h2B41,4);
TASK_PP(16'h2B42,4);
TASK_PP(16'h2B43,4);
TASK_PP(16'h2B44,4);
TASK_PP(16'h2B45,4);
TASK_PP(16'h2B46,4);
TASK_PP(16'h2B47,4);
TASK_PP(16'h2B48,4);
TASK_PP(16'h2B49,4);
TASK_PP(16'h2B4A,4);
TASK_PP(16'h2B4B,4);
TASK_PP(16'h2B4C,4);
TASK_PP(16'h2B4D,4);
TASK_PP(16'h2B4E,4);
TASK_PP(16'h2B4F,4);
TASK_PP(16'h2B50,4);
TASK_PP(16'h2B51,4);
TASK_PP(16'h2B52,4);
TASK_PP(16'h2B53,4);
TASK_PP(16'h2B54,4);
TASK_PP(16'h2B55,4);
TASK_PP(16'h2B56,4);
TASK_PP(16'h2B57,4);
TASK_PP(16'h2B58,4);
TASK_PP(16'h2B59,4);
TASK_PP(16'h2B5A,4);
TASK_PP(16'h2B5B,4);
TASK_PP(16'h2B5C,4);
TASK_PP(16'h2B5D,4);
TASK_PP(16'h2B5E,4);
TASK_PP(16'h2B5F,4);
TASK_PP(16'h2B60,4);
TASK_PP(16'h2B61,4);
TASK_PP(16'h2B62,4);
TASK_PP(16'h2B63,4);
TASK_PP(16'h2B64,4);
TASK_PP(16'h2B65,4);
TASK_PP(16'h2B66,4);
TASK_PP(16'h2B67,4);
TASK_PP(16'h2B68,4);
TASK_PP(16'h2B69,4);
TASK_PP(16'h2B6A,4);
TASK_PP(16'h2B6B,4);
TASK_PP(16'h2B6C,4);
TASK_PP(16'h2B6D,4);
TASK_PP(16'h2B6E,4);
TASK_PP(16'h2B6F,4);
TASK_PP(16'h2B70,4);
TASK_PP(16'h2B71,4);
TASK_PP(16'h2B72,4);
TASK_PP(16'h2B73,4);
TASK_PP(16'h2B74,4);
TASK_PP(16'h2B75,4);
TASK_PP(16'h2B76,4);
TASK_PP(16'h2B77,4);
TASK_PP(16'h2B78,4);
TASK_PP(16'h2B79,4);
TASK_PP(16'h2B7A,4);
TASK_PP(16'h2B7B,4);
TASK_PP(16'h2B7C,4);
TASK_PP(16'h2B7D,4);
TASK_PP(16'h2B7E,4);
TASK_PP(16'h2B7F,4);
TASK_PP(16'h2B80,4);
TASK_PP(16'h2B81,4);
TASK_PP(16'h2B82,4);
TASK_PP(16'h2B83,4);
TASK_PP(16'h2B84,4);
TASK_PP(16'h2B85,4);
TASK_PP(16'h2B86,4);
TASK_PP(16'h2B87,4);
TASK_PP(16'h2B88,4);
TASK_PP(16'h2B89,4);
TASK_PP(16'h2B8A,4);
TASK_PP(16'h2B8B,4);
TASK_PP(16'h2B8C,4);
TASK_PP(16'h2B8D,4);
TASK_PP(16'h2B8E,4);
TASK_PP(16'h2B8F,4);
TASK_PP(16'h2B90,4);
TASK_PP(16'h2B91,4);
TASK_PP(16'h2B92,4);
TASK_PP(16'h2B93,4);
TASK_PP(16'h2B94,4);
TASK_PP(16'h2B95,4);
TASK_PP(16'h2B96,4);
TASK_PP(16'h2B97,4);
TASK_PP(16'h2B98,4);
TASK_PP(16'h2B99,4);
TASK_PP(16'h2B9A,4);
TASK_PP(16'h2B9B,4);
TASK_PP(16'h2B9C,4);
TASK_PP(16'h2B9D,4);
TASK_PP(16'h2B9E,4);
TASK_PP(16'h2B9F,4);
TASK_PP(16'h2BA0,4);
TASK_PP(16'h2BA1,4);
TASK_PP(16'h2BA2,4);
TASK_PP(16'h2BA3,4);
TASK_PP(16'h2BA4,4);
TASK_PP(16'h2BA5,4);
TASK_PP(16'h2BA6,4);
TASK_PP(16'h2BA7,4);
TASK_PP(16'h2BA8,4);
TASK_PP(16'h2BA9,4);
TASK_PP(16'h2BAA,4);
TASK_PP(16'h2BAB,4);
TASK_PP(16'h2BAC,4);
TASK_PP(16'h2BAD,4);
TASK_PP(16'h2BAE,4);
TASK_PP(16'h2BAF,4);
TASK_PP(16'h2BB0,4);
TASK_PP(16'h2BB1,4);
TASK_PP(16'h2BB2,4);
TASK_PP(16'h2BB3,4);
TASK_PP(16'h2BB4,4);
TASK_PP(16'h2BB5,4);
TASK_PP(16'h2BB6,4);
TASK_PP(16'h2BB7,4);
TASK_PP(16'h2BB8,4);
TASK_PP(16'h2BB9,4);
TASK_PP(16'h2BBA,4);
TASK_PP(16'h2BBB,4);
TASK_PP(16'h2BBC,4);
TASK_PP(16'h2BBD,4);
TASK_PP(16'h2BBE,4);
TASK_PP(16'h2BBF,4);
TASK_PP(16'h2BC0,4);
TASK_PP(16'h2BC1,4);
TASK_PP(16'h2BC2,4);
TASK_PP(16'h2BC3,4);
TASK_PP(16'h2BC4,4);
TASK_PP(16'h2BC5,4);
TASK_PP(16'h2BC6,4);
TASK_PP(16'h2BC7,4);
TASK_PP(16'h2BC8,4);
TASK_PP(16'h2BC9,4);
TASK_PP(16'h2BCA,4);
TASK_PP(16'h2BCB,4);
TASK_PP(16'h2BCC,4);
TASK_PP(16'h2BCD,4);
TASK_PP(16'h2BCE,4);
TASK_PP(16'h2BCF,4);
TASK_PP(16'h2BD0,4);
TASK_PP(16'h2BD1,4);
TASK_PP(16'h2BD2,4);
TASK_PP(16'h2BD3,4);
TASK_PP(16'h2BD4,4);
TASK_PP(16'h2BD5,4);
TASK_PP(16'h2BD6,4);
TASK_PP(16'h2BD7,4);
TASK_PP(16'h2BD8,4);
TASK_PP(16'h2BD9,4);
TASK_PP(16'h2BDA,4);
TASK_PP(16'h2BDB,4);
TASK_PP(16'h2BDC,4);
TASK_PP(16'h2BDD,4);
TASK_PP(16'h2BDE,4);
TASK_PP(16'h2BDF,4);
TASK_PP(16'h2BE0,4);
TASK_PP(16'h2BE1,4);
TASK_PP(16'h2BE2,4);
TASK_PP(16'h2BE3,4);
TASK_PP(16'h2BE4,4);
TASK_PP(16'h2BE5,4);
TASK_PP(16'h2BE6,4);
TASK_PP(16'h2BE7,4);
TASK_PP(16'h2BE8,4);
TASK_PP(16'h2BE9,4);
TASK_PP(16'h2BEA,4);
TASK_PP(16'h2BEB,4);
TASK_PP(16'h2BEC,4);
TASK_PP(16'h2BED,4);
TASK_PP(16'h2BEE,4);
TASK_PP(16'h2BEF,4);
TASK_PP(16'h2BF0,4);
TASK_PP(16'h2BF1,4);
TASK_PP(16'h2BF2,4);
TASK_PP(16'h2BF3,4);
TASK_PP(16'h2BF4,4);
TASK_PP(16'h2BF5,4);
TASK_PP(16'h2BF6,4);
TASK_PP(16'h2BF7,4);
TASK_PP(16'h2BF8,4);
TASK_PP(16'h2BF9,4);
TASK_PP(16'h2BFA,4);
TASK_PP(16'h2BFB,4);
TASK_PP(16'h2BFC,4);
TASK_PP(16'h2BFD,4);
TASK_PP(16'h2BFE,4);
TASK_PP(16'h2BFF,4);
TASK_PP(16'h2C00,4);
TASK_PP(16'h2C01,4);
TASK_PP(16'h2C02,4);
TASK_PP(16'h2C03,4);
TASK_PP(16'h2C04,4);
TASK_PP(16'h2C05,4);
TASK_PP(16'h2C06,4);
TASK_PP(16'h2C07,4);
TASK_PP(16'h2C08,4);
TASK_PP(16'h2C09,4);
TASK_PP(16'h2C0A,4);
TASK_PP(16'h2C0B,4);
TASK_PP(16'h2C0C,4);
TASK_PP(16'h2C0D,4);
TASK_PP(16'h2C0E,4);
TASK_PP(16'h2C0F,4);
TASK_PP(16'h2C10,4);
TASK_PP(16'h2C11,4);
TASK_PP(16'h2C12,4);
TASK_PP(16'h2C13,4);
TASK_PP(16'h2C14,4);
TASK_PP(16'h2C15,4);
TASK_PP(16'h2C16,4);
TASK_PP(16'h2C17,4);
TASK_PP(16'h2C18,4);
TASK_PP(16'h2C19,4);
TASK_PP(16'h2C1A,4);
TASK_PP(16'h2C1B,4);
TASK_PP(16'h2C1C,4);
TASK_PP(16'h2C1D,4);
TASK_PP(16'h2C1E,4);
TASK_PP(16'h2C1F,4);
TASK_PP(16'h2C20,4);
TASK_PP(16'h2C21,4);
TASK_PP(16'h2C22,4);
TASK_PP(16'h2C23,4);
TASK_PP(16'h2C24,4);
TASK_PP(16'h2C25,4);
TASK_PP(16'h2C26,4);
TASK_PP(16'h2C27,4);
TASK_PP(16'h2C28,4);
TASK_PP(16'h2C29,4);
TASK_PP(16'h2C2A,4);
TASK_PP(16'h2C2B,4);
TASK_PP(16'h2C2C,4);
TASK_PP(16'h2C2D,4);
TASK_PP(16'h2C2E,4);
TASK_PP(16'h2C2F,4);
TASK_PP(16'h2C30,4);
TASK_PP(16'h2C31,4);
TASK_PP(16'h2C32,4);
TASK_PP(16'h2C33,4);
TASK_PP(16'h2C34,4);
TASK_PP(16'h2C35,4);
TASK_PP(16'h2C36,4);
TASK_PP(16'h2C37,4);
TASK_PP(16'h2C38,4);
TASK_PP(16'h2C39,4);
TASK_PP(16'h2C3A,4);
TASK_PP(16'h2C3B,4);
TASK_PP(16'h2C3C,4);
TASK_PP(16'h2C3D,4);
TASK_PP(16'h2C3E,4);
TASK_PP(16'h2C3F,4);
TASK_PP(16'h2C40,4);
TASK_PP(16'h2C41,4);
TASK_PP(16'h2C42,4);
TASK_PP(16'h2C43,4);
TASK_PP(16'h2C44,4);
TASK_PP(16'h2C45,4);
TASK_PP(16'h2C46,4);
TASK_PP(16'h2C47,4);
TASK_PP(16'h2C48,4);
TASK_PP(16'h2C49,4);
TASK_PP(16'h2C4A,4);
TASK_PP(16'h2C4B,4);
TASK_PP(16'h2C4C,4);
TASK_PP(16'h2C4D,4);
TASK_PP(16'h2C4E,4);
TASK_PP(16'h2C4F,4);
TASK_PP(16'h2C50,4);
TASK_PP(16'h2C51,4);
TASK_PP(16'h2C52,4);
TASK_PP(16'h2C53,4);
TASK_PP(16'h2C54,4);
TASK_PP(16'h2C55,4);
TASK_PP(16'h2C56,4);
TASK_PP(16'h2C57,4);
TASK_PP(16'h2C58,4);
TASK_PP(16'h2C59,4);
TASK_PP(16'h2C5A,4);
TASK_PP(16'h2C5B,4);
TASK_PP(16'h2C5C,4);
TASK_PP(16'h2C5D,4);
TASK_PP(16'h2C5E,4);
TASK_PP(16'h2C5F,4);
TASK_PP(16'h2C60,4);
TASK_PP(16'h2C61,4);
TASK_PP(16'h2C62,4);
TASK_PP(16'h2C63,4);
TASK_PP(16'h2C64,4);
TASK_PP(16'h2C65,4);
TASK_PP(16'h2C66,4);
TASK_PP(16'h2C67,4);
TASK_PP(16'h2C68,4);
TASK_PP(16'h2C69,4);
TASK_PP(16'h2C6A,4);
TASK_PP(16'h2C6B,4);
TASK_PP(16'h2C6C,4);
TASK_PP(16'h2C6D,4);
TASK_PP(16'h2C6E,4);
TASK_PP(16'h2C6F,4);
TASK_PP(16'h2C70,4);
TASK_PP(16'h2C71,4);
TASK_PP(16'h2C72,4);
TASK_PP(16'h2C73,4);
TASK_PP(16'h2C74,4);
TASK_PP(16'h2C75,4);
TASK_PP(16'h2C76,4);
TASK_PP(16'h2C77,4);
TASK_PP(16'h2C78,4);
TASK_PP(16'h2C79,4);
TASK_PP(16'h2C7A,4);
TASK_PP(16'h2C7B,4);
TASK_PP(16'h2C7C,4);
TASK_PP(16'h2C7D,4);
TASK_PP(16'h2C7E,4);
TASK_PP(16'h2C7F,4);
TASK_PP(16'h2C80,4);
TASK_PP(16'h2C81,4);
TASK_PP(16'h2C82,4);
TASK_PP(16'h2C83,4);
TASK_PP(16'h2C84,4);
TASK_PP(16'h2C85,4);
TASK_PP(16'h2C86,4);
TASK_PP(16'h2C87,4);
TASK_PP(16'h2C88,4);
TASK_PP(16'h2C89,4);
TASK_PP(16'h2C8A,4);
TASK_PP(16'h2C8B,4);
TASK_PP(16'h2C8C,4);
TASK_PP(16'h2C8D,4);
TASK_PP(16'h2C8E,4);
TASK_PP(16'h2C8F,4);
TASK_PP(16'h2C90,4);
TASK_PP(16'h2C91,4);
TASK_PP(16'h2C92,4);
TASK_PP(16'h2C93,4);
TASK_PP(16'h2C94,4);
TASK_PP(16'h2C95,4);
TASK_PP(16'h2C96,4);
TASK_PP(16'h2C97,4);
TASK_PP(16'h2C98,4);
TASK_PP(16'h2C99,4);
TASK_PP(16'h2C9A,4);
TASK_PP(16'h2C9B,4);
TASK_PP(16'h2C9C,4);
TASK_PP(16'h2C9D,4);
TASK_PP(16'h2C9E,4);
TASK_PP(16'h2C9F,4);
TASK_PP(16'h2CA0,4);
TASK_PP(16'h2CA1,4);
TASK_PP(16'h2CA2,4);
TASK_PP(16'h2CA3,4);
TASK_PP(16'h2CA4,4);
TASK_PP(16'h2CA5,4);
TASK_PP(16'h2CA6,4);
TASK_PP(16'h2CA7,4);
TASK_PP(16'h2CA8,4);
TASK_PP(16'h2CA9,4);
TASK_PP(16'h2CAA,4);
TASK_PP(16'h2CAB,4);
TASK_PP(16'h2CAC,4);
TASK_PP(16'h2CAD,4);
TASK_PP(16'h2CAE,4);
TASK_PP(16'h2CAF,4);
TASK_PP(16'h2CB0,4);
TASK_PP(16'h2CB1,4);
TASK_PP(16'h2CB2,4);
TASK_PP(16'h2CB3,4);
TASK_PP(16'h2CB4,4);
TASK_PP(16'h2CB5,4);
TASK_PP(16'h2CB6,4);
TASK_PP(16'h2CB7,4);
TASK_PP(16'h2CB8,4);
TASK_PP(16'h2CB9,4);
TASK_PP(16'h2CBA,4);
TASK_PP(16'h2CBB,4);
TASK_PP(16'h2CBC,4);
TASK_PP(16'h2CBD,4);
TASK_PP(16'h2CBE,4);
TASK_PP(16'h2CBF,4);
TASK_PP(16'h2CC0,4);
TASK_PP(16'h2CC1,4);
TASK_PP(16'h2CC2,4);
TASK_PP(16'h2CC3,4);
TASK_PP(16'h2CC4,4);
TASK_PP(16'h2CC5,4);
TASK_PP(16'h2CC6,4);
TASK_PP(16'h2CC7,4);
TASK_PP(16'h2CC8,4);
TASK_PP(16'h2CC9,4);
TASK_PP(16'h2CCA,4);
TASK_PP(16'h2CCB,4);
TASK_PP(16'h2CCC,4);
TASK_PP(16'h2CCD,4);
TASK_PP(16'h2CCE,4);
TASK_PP(16'h2CCF,4);
TASK_PP(16'h2CD0,4);
TASK_PP(16'h2CD1,4);
TASK_PP(16'h2CD2,4);
TASK_PP(16'h2CD3,4);
TASK_PP(16'h2CD4,4);
TASK_PP(16'h2CD5,4);
TASK_PP(16'h2CD6,4);
TASK_PP(16'h2CD7,4);
TASK_PP(16'h2CD8,4);
TASK_PP(16'h2CD9,4);
TASK_PP(16'h2CDA,4);
TASK_PP(16'h2CDB,4);
TASK_PP(16'h2CDC,4);
TASK_PP(16'h2CDD,4);
TASK_PP(16'h2CDE,4);
TASK_PP(16'h2CDF,4);
TASK_PP(16'h2CE0,4);
TASK_PP(16'h2CE1,4);
TASK_PP(16'h2CE2,4);
TASK_PP(16'h2CE3,4);
TASK_PP(16'h2CE4,4);
TASK_PP(16'h2CE5,4);
TASK_PP(16'h2CE6,4);
TASK_PP(16'h2CE7,4);
TASK_PP(16'h2CE8,4);
TASK_PP(16'h2CE9,4);
TASK_PP(16'h2CEA,4);
TASK_PP(16'h2CEB,4);
TASK_PP(16'h2CEC,4);
TASK_PP(16'h2CED,4);
TASK_PP(16'h2CEE,4);
TASK_PP(16'h2CEF,4);
TASK_PP(16'h2CF0,4);
TASK_PP(16'h2CF1,4);
TASK_PP(16'h2CF2,4);
TASK_PP(16'h2CF3,4);
TASK_PP(16'h2CF4,4);
TASK_PP(16'h2CF5,4);
TASK_PP(16'h2CF6,4);
TASK_PP(16'h2CF7,4);
TASK_PP(16'h2CF8,4);
TASK_PP(16'h2CF9,4);
TASK_PP(16'h2CFA,4);
TASK_PP(16'h2CFB,4);
TASK_PP(16'h2CFC,4);
TASK_PP(16'h2CFD,4);
TASK_PP(16'h2CFE,4);
TASK_PP(16'h2CFF,4);
TASK_PP(16'h2D00,4);
TASK_PP(16'h2D01,4);
TASK_PP(16'h2D02,4);
TASK_PP(16'h2D03,4);
TASK_PP(16'h2D04,4);
TASK_PP(16'h2D05,4);
TASK_PP(16'h2D06,4);
TASK_PP(16'h2D07,4);
TASK_PP(16'h2D08,4);
TASK_PP(16'h2D09,4);
TASK_PP(16'h2D0A,4);
TASK_PP(16'h2D0B,4);
TASK_PP(16'h2D0C,4);
TASK_PP(16'h2D0D,4);
TASK_PP(16'h2D0E,4);
TASK_PP(16'h2D0F,4);
TASK_PP(16'h2D10,4);
TASK_PP(16'h2D11,4);
TASK_PP(16'h2D12,4);
TASK_PP(16'h2D13,4);
TASK_PP(16'h2D14,4);
TASK_PP(16'h2D15,4);
TASK_PP(16'h2D16,4);
TASK_PP(16'h2D17,4);
TASK_PP(16'h2D18,4);
TASK_PP(16'h2D19,4);
TASK_PP(16'h2D1A,4);
TASK_PP(16'h2D1B,4);
TASK_PP(16'h2D1C,4);
TASK_PP(16'h2D1D,4);
TASK_PP(16'h2D1E,4);
TASK_PP(16'h2D1F,4);
TASK_PP(16'h2D20,4);
TASK_PP(16'h2D21,4);
TASK_PP(16'h2D22,4);
TASK_PP(16'h2D23,4);
TASK_PP(16'h2D24,4);
TASK_PP(16'h2D25,4);
TASK_PP(16'h2D26,4);
TASK_PP(16'h2D27,4);
TASK_PP(16'h2D28,4);
TASK_PP(16'h2D29,4);
TASK_PP(16'h2D2A,4);
TASK_PP(16'h2D2B,4);
TASK_PP(16'h2D2C,4);
TASK_PP(16'h2D2D,4);
TASK_PP(16'h2D2E,4);
TASK_PP(16'h2D2F,4);
TASK_PP(16'h2D30,4);
TASK_PP(16'h2D31,4);
TASK_PP(16'h2D32,4);
TASK_PP(16'h2D33,4);
TASK_PP(16'h2D34,4);
TASK_PP(16'h2D35,4);
TASK_PP(16'h2D36,4);
TASK_PP(16'h2D37,4);
TASK_PP(16'h2D38,4);
TASK_PP(16'h2D39,4);
TASK_PP(16'h2D3A,4);
TASK_PP(16'h2D3B,4);
TASK_PP(16'h2D3C,4);
TASK_PP(16'h2D3D,4);
TASK_PP(16'h2D3E,4);
TASK_PP(16'h2D3F,4);
TASK_PP(16'h2D40,4);
TASK_PP(16'h2D41,4);
TASK_PP(16'h2D42,4);
TASK_PP(16'h2D43,4);
TASK_PP(16'h2D44,4);
TASK_PP(16'h2D45,4);
TASK_PP(16'h2D46,4);
TASK_PP(16'h2D47,4);
TASK_PP(16'h2D48,4);
TASK_PP(16'h2D49,4);
TASK_PP(16'h2D4A,4);
TASK_PP(16'h2D4B,4);
TASK_PP(16'h2D4C,4);
TASK_PP(16'h2D4D,4);
TASK_PP(16'h2D4E,4);
TASK_PP(16'h2D4F,4);
TASK_PP(16'h2D50,4);
TASK_PP(16'h2D51,4);
TASK_PP(16'h2D52,4);
TASK_PP(16'h2D53,4);
TASK_PP(16'h2D54,4);
TASK_PP(16'h2D55,4);
TASK_PP(16'h2D56,4);
TASK_PP(16'h2D57,4);
TASK_PP(16'h2D58,4);
TASK_PP(16'h2D59,4);
TASK_PP(16'h2D5A,4);
TASK_PP(16'h2D5B,4);
TASK_PP(16'h2D5C,4);
TASK_PP(16'h2D5D,4);
TASK_PP(16'h2D5E,4);
TASK_PP(16'h2D5F,4);
TASK_PP(16'h2D60,4);
TASK_PP(16'h2D61,4);
TASK_PP(16'h2D62,4);
TASK_PP(16'h2D63,4);
TASK_PP(16'h2D64,4);
TASK_PP(16'h2D65,4);
TASK_PP(16'h2D66,4);
TASK_PP(16'h2D67,4);
TASK_PP(16'h2D68,4);
TASK_PP(16'h2D69,4);
TASK_PP(16'h2D6A,4);
TASK_PP(16'h2D6B,4);
TASK_PP(16'h2D6C,4);
TASK_PP(16'h2D6D,4);
TASK_PP(16'h2D6E,4);
TASK_PP(16'h2D6F,4);
TASK_PP(16'h2D70,4);
TASK_PP(16'h2D71,4);
TASK_PP(16'h2D72,4);
TASK_PP(16'h2D73,4);
TASK_PP(16'h2D74,4);
TASK_PP(16'h2D75,4);
TASK_PP(16'h2D76,4);
TASK_PP(16'h2D77,4);
TASK_PP(16'h2D78,4);
TASK_PP(16'h2D79,4);
TASK_PP(16'h2D7A,4);
TASK_PP(16'h2D7B,4);
TASK_PP(16'h2D7C,4);
TASK_PP(16'h2D7D,4);
TASK_PP(16'h2D7E,4);
TASK_PP(16'h2D7F,4);
TASK_PP(16'h2D80,4);
TASK_PP(16'h2D81,4);
TASK_PP(16'h2D82,4);
TASK_PP(16'h2D83,4);
TASK_PP(16'h2D84,4);
TASK_PP(16'h2D85,4);
TASK_PP(16'h2D86,4);
TASK_PP(16'h2D87,4);
TASK_PP(16'h2D88,4);
TASK_PP(16'h2D89,4);
TASK_PP(16'h2D8A,4);
TASK_PP(16'h2D8B,4);
TASK_PP(16'h2D8C,4);
TASK_PP(16'h2D8D,4);
TASK_PP(16'h2D8E,4);
TASK_PP(16'h2D8F,4);
TASK_PP(16'h2D90,4);
TASK_PP(16'h2D91,4);
TASK_PP(16'h2D92,4);
TASK_PP(16'h2D93,4);
TASK_PP(16'h2D94,4);
TASK_PP(16'h2D95,4);
TASK_PP(16'h2D96,4);
TASK_PP(16'h2D97,4);
TASK_PP(16'h2D98,4);
TASK_PP(16'h2D99,4);
TASK_PP(16'h2D9A,4);
TASK_PP(16'h2D9B,4);
TASK_PP(16'h2D9C,4);
TASK_PP(16'h2D9D,4);
TASK_PP(16'h2D9E,4);
TASK_PP(16'h2D9F,4);
TASK_PP(16'h2DA0,4);
TASK_PP(16'h2DA1,4);
TASK_PP(16'h2DA2,4);
TASK_PP(16'h2DA3,4);
TASK_PP(16'h2DA4,4);
TASK_PP(16'h2DA5,4);
TASK_PP(16'h2DA6,4);
TASK_PP(16'h2DA7,4);
TASK_PP(16'h2DA8,4);
TASK_PP(16'h2DA9,4);
TASK_PP(16'h2DAA,4);
TASK_PP(16'h2DAB,4);
TASK_PP(16'h2DAC,4);
TASK_PP(16'h2DAD,4);
TASK_PP(16'h2DAE,4);
TASK_PP(16'h2DAF,4);
TASK_PP(16'h2DB0,4);
TASK_PP(16'h2DB1,4);
TASK_PP(16'h2DB2,4);
TASK_PP(16'h2DB3,4);
TASK_PP(16'h2DB4,4);
TASK_PP(16'h2DB5,4);
TASK_PP(16'h2DB6,4);
TASK_PP(16'h2DB7,4);
TASK_PP(16'h2DB8,4);
TASK_PP(16'h2DB9,4);
TASK_PP(16'h2DBA,4);
TASK_PP(16'h2DBB,4);
TASK_PP(16'h2DBC,4);
TASK_PP(16'h2DBD,4);
TASK_PP(16'h2DBE,4);
TASK_PP(16'h2DBF,4);
TASK_PP(16'h2DC0,4);
TASK_PP(16'h2DC1,4);
TASK_PP(16'h2DC2,4);
TASK_PP(16'h2DC3,4);
TASK_PP(16'h2DC4,4);
TASK_PP(16'h2DC5,4);
TASK_PP(16'h2DC6,4);
TASK_PP(16'h2DC7,4);
TASK_PP(16'h2DC8,4);
TASK_PP(16'h2DC9,4);
TASK_PP(16'h2DCA,4);
TASK_PP(16'h2DCB,4);
TASK_PP(16'h2DCC,4);
TASK_PP(16'h2DCD,4);
TASK_PP(16'h2DCE,4);
TASK_PP(16'h2DCF,4);
TASK_PP(16'h2DD0,4);
TASK_PP(16'h2DD1,4);
TASK_PP(16'h2DD2,4);
TASK_PP(16'h2DD3,4);
TASK_PP(16'h2DD4,4);
TASK_PP(16'h2DD5,4);
TASK_PP(16'h2DD6,4);
TASK_PP(16'h2DD7,4);
TASK_PP(16'h2DD8,4);
TASK_PP(16'h2DD9,4);
TASK_PP(16'h2DDA,4);
TASK_PP(16'h2DDB,4);
TASK_PP(16'h2DDC,4);
TASK_PP(16'h2DDD,4);
TASK_PP(16'h2DDE,4);
TASK_PP(16'h2DDF,4);
TASK_PP(16'h2DE0,4);
TASK_PP(16'h2DE1,4);
TASK_PP(16'h2DE2,4);
TASK_PP(16'h2DE3,4);
TASK_PP(16'h2DE4,4);
TASK_PP(16'h2DE5,4);
TASK_PP(16'h2DE6,4);
TASK_PP(16'h2DE7,4);
TASK_PP(16'h2DE8,4);
TASK_PP(16'h2DE9,4);
TASK_PP(16'h2DEA,4);
TASK_PP(16'h2DEB,4);
TASK_PP(16'h2DEC,4);
TASK_PP(16'h2DED,4);
TASK_PP(16'h2DEE,4);
TASK_PP(16'h2DEF,4);
TASK_PP(16'h2DF0,4);
TASK_PP(16'h2DF1,4);
TASK_PP(16'h2DF2,4);
TASK_PP(16'h2DF3,4);
TASK_PP(16'h2DF4,4);
TASK_PP(16'h2DF5,4);
TASK_PP(16'h2DF6,4);
TASK_PP(16'h2DF7,4);
TASK_PP(16'h2DF8,4);
TASK_PP(16'h2DF9,4);
TASK_PP(16'h2DFA,4);
TASK_PP(16'h2DFB,4);
TASK_PP(16'h2DFC,4);
TASK_PP(16'h2DFD,4);
TASK_PP(16'h2DFE,4);
TASK_PP(16'h2DFF,4);
TASK_PP(16'h2E00,4);
TASK_PP(16'h2E01,4);
TASK_PP(16'h2E02,4);
TASK_PP(16'h2E03,4);
TASK_PP(16'h2E04,4);
TASK_PP(16'h2E05,4);
TASK_PP(16'h2E06,4);
TASK_PP(16'h2E07,4);
TASK_PP(16'h2E08,4);
TASK_PP(16'h2E09,4);
TASK_PP(16'h2E0A,4);
TASK_PP(16'h2E0B,4);
TASK_PP(16'h2E0C,4);
TASK_PP(16'h2E0D,4);
TASK_PP(16'h2E0E,4);
TASK_PP(16'h2E0F,4);
TASK_PP(16'h2E10,4);
TASK_PP(16'h2E11,4);
TASK_PP(16'h2E12,4);
TASK_PP(16'h2E13,4);
TASK_PP(16'h2E14,4);
TASK_PP(16'h2E15,4);
TASK_PP(16'h2E16,4);
TASK_PP(16'h2E17,4);
TASK_PP(16'h2E18,4);
TASK_PP(16'h2E19,4);
TASK_PP(16'h2E1A,4);
TASK_PP(16'h2E1B,4);
TASK_PP(16'h2E1C,4);
TASK_PP(16'h2E1D,4);
TASK_PP(16'h2E1E,4);
TASK_PP(16'h2E1F,4);
TASK_PP(16'h2E20,4);
TASK_PP(16'h2E21,4);
TASK_PP(16'h2E22,4);
TASK_PP(16'h2E23,4);
TASK_PP(16'h2E24,4);
TASK_PP(16'h2E25,4);
TASK_PP(16'h2E26,4);
TASK_PP(16'h2E27,4);
TASK_PP(16'h2E28,4);
TASK_PP(16'h2E29,4);
TASK_PP(16'h2E2A,4);
TASK_PP(16'h2E2B,4);
TASK_PP(16'h2E2C,4);
TASK_PP(16'h2E2D,4);
TASK_PP(16'h2E2E,4);
TASK_PP(16'h2E2F,4);
TASK_PP(16'h2E30,4);
TASK_PP(16'h2E31,4);
TASK_PP(16'h2E32,4);
TASK_PP(16'h2E33,4);
TASK_PP(16'h2E34,4);
TASK_PP(16'h2E35,4);
TASK_PP(16'h2E36,4);
TASK_PP(16'h2E37,4);
TASK_PP(16'h2E38,4);
TASK_PP(16'h2E39,4);
TASK_PP(16'h2E3A,4);
TASK_PP(16'h2E3B,4);
TASK_PP(16'h2E3C,4);
TASK_PP(16'h2E3D,4);
TASK_PP(16'h2E3E,4);
TASK_PP(16'h2E3F,4);
TASK_PP(16'h2E40,4);
TASK_PP(16'h2E41,4);
TASK_PP(16'h2E42,4);
TASK_PP(16'h2E43,4);
TASK_PP(16'h2E44,4);
TASK_PP(16'h2E45,4);
TASK_PP(16'h2E46,4);
TASK_PP(16'h2E47,4);
TASK_PP(16'h2E48,4);
TASK_PP(16'h2E49,4);
TASK_PP(16'h2E4A,4);
TASK_PP(16'h2E4B,4);
TASK_PP(16'h2E4C,4);
TASK_PP(16'h2E4D,4);
TASK_PP(16'h2E4E,4);
TASK_PP(16'h2E4F,4);
TASK_PP(16'h2E50,4);
TASK_PP(16'h2E51,4);
TASK_PP(16'h2E52,4);
TASK_PP(16'h2E53,4);
TASK_PP(16'h2E54,4);
TASK_PP(16'h2E55,4);
TASK_PP(16'h2E56,4);
TASK_PP(16'h2E57,4);
TASK_PP(16'h2E58,4);
TASK_PP(16'h2E59,4);
TASK_PP(16'h2E5A,4);
TASK_PP(16'h2E5B,4);
TASK_PP(16'h2E5C,4);
TASK_PP(16'h2E5D,4);
TASK_PP(16'h2E5E,4);
TASK_PP(16'h2E5F,4);
TASK_PP(16'h2E60,4);
TASK_PP(16'h2E61,4);
TASK_PP(16'h2E62,4);
TASK_PP(16'h2E63,4);
TASK_PP(16'h2E64,4);
TASK_PP(16'h2E65,4);
TASK_PP(16'h2E66,4);
TASK_PP(16'h2E67,4);
TASK_PP(16'h2E68,4);
TASK_PP(16'h2E69,4);
TASK_PP(16'h2E6A,4);
TASK_PP(16'h2E6B,4);
TASK_PP(16'h2E6C,4);
TASK_PP(16'h2E6D,4);
TASK_PP(16'h2E6E,4);
TASK_PP(16'h2E6F,4);
TASK_PP(16'h2E70,4);
TASK_PP(16'h2E71,4);
TASK_PP(16'h2E72,4);
TASK_PP(16'h2E73,4);
TASK_PP(16'h2E74,4);
TASK_PP(16'h2E75,4);
TASK_PP(16'h2E76,4);
TASK_PP(16'h2E77,4);
TASK_PP(16'h2E78,4);
TASK_PP(16'h2E79,4);
TASK_PP(16'h2E7A,4);
TASK_PP(16'h2E7B,4);
TASK_PP(16'h2E7C,4);
TASK_PP(16'h2E7D,4);
TASK_PP(16'h2E7E,4);
TASK_PP(16'h2E7F,4);
TASK_PP(16'h2E80,4);
TASK_PP(16'h2E81,4);
TASK_PP(16'h2E82,4);
TASK_PP(16'h2E83,4);
TASK_PP(16'h2E84,4);
TASK_PP(16'h2E85,4);
TASK_PP(16'h2E86,4);
TASK_PP(16'h2E87,4);
TASK_PP(16'h2E88,4);
TASK_PP(16'h2E89,4);
TASK_PP(16'h2E8A,4);
TASK_PP(16'h2E8B,4);
TASK_PP(16'h2E8C,4);
TASK_PP(16'h2E8D,4);
TASK_PP(16'h2E8E,4);
TASK_PP(16'h2E8F,4);
TASK_PP(16'h2E90,4);
TASK_PP(16'h2E91,4);
TASK_PP(16'h2E92,4);
TASK_PP(16'h2E93,4);
TASK_PP(16'h2E94,4);
TASK_PP(16'h2E95,4);
TASK_PP(16'h2E96,4);
TASK_PP(16'h2E97,4);
TASK_PP(16'h2E98,4);
TASK_PP(16'h2E99,4);
TASK_PP(16'h2E9A,4);
TASK_PP(16'h2E9B,4);
TASK_PP(16'h2E9C,4);
TASK_PP(16'h2E9D,4);
TASK_PP(16'h2E9E,4);
TASK_PP(16'h2E9F,4);
TASK_PP(16'h2EA0,4);
TASK_PP(16'h2EA1,4);
TASK_PP(16'h2EA2,4);
TASK_PP(16'h2EA3,4);
TASK_PP(16'h2EA4,4);
TASK_PP(16'h2EA5,4);
TASK_PP(16'h2EA6,4);
TASK_PP(16'h2EA7,4);
TASK_PP(16'h2EA8,4);
TASK_PP(16'h2EA9,4);
TASK_PP(16'h2EAA,4);
TASK_PP(16'h2EAB,4);
TASK_PP(16'h2EAC,4);
TASK_PP(16'h2EAD,4);
TASK_PP(16'h2EAE,4);
TASK_PP(16'h2EAF,4);
TASK_PP(16'h2EB0,4);
TASK_PP(16'h2EB1,4);
TASK_PP(16'h2EB2,4);
TASK_PP(16'h2EB3,4);
TASK_PP(16'h2EB4,4);
TASK_PP(16'h2EB5,4);
TASK_PP(16'h2EB6,4);
TASK_PP(16'h2EB7,4);
TASK_PP(16'h2EB8,4);
TASK_PP(16'h2EB9,4);
TASK_PP(16'h2EBA,4);
TASK_PP(16'h2EBB,4);
TASK_PP(16'h2EBC,4);
TASK_PP(16'h2EBD,4);
TASK_PP(16'h2EBE,4);
TASK_PP(16'h2EBF,4);
TASK_PP(16'h2EC0,4);
TASK_PP(16'h2EC1,4);
TASK_PP(16'h2EC2,4);
TASK_PP(16'h2EC3,4);
TASK_PP(16'h2EC4,4);
TASK_PP(16'h2EC5,4);
TASK_PP(16'h2EC6,4);
TASK_PP(16'h2EC7,4);
TASK_PP(16'h2EC8,4);
TASK_PP(16'h2EC9,4);
TASK_PP(16'h2ECA,4);
TASK_PP(16'h2ECB,4);
TASK_PP(16'h2ECC,4);
TASK_PP(16'h2ECD,4);
TASK_PP(16'h2ECE,4);
TASK_PP(16'h2ECF,4);
TASK_PP(16'h2ED0,4);
TASK_PP(16'h2ED1,4);
TASK_PP(16'h2ED2,4);
TASK_PP(16'h2ED3,4);
TASK_PP(16'h2ED4,4);
TASK_PP(16'h2ED5,4);
TASK_PP(16'h2ED6,4);
TASK_PP(16'h2ED7,4);
TASK_PP(16'h2ED8,4);
TASK_PP(16'h2ED9,4);
TASK_PP(16'h2EDA,4);
TASK_PP(16'h2EDB,4);
TASK_PP(16'h2EDC,4);
TASK_PP(16'h2EDD,4);
TASK_PP(16'h2EDE,4);
TASK_PP(16'h2EDF,4);
TASK_PP(16'h2EE0,4);
TASK_PP(16'h2EE1,4);
TASK_PP(16'h2EE2,4);
TASK_PP(16'h2EE3,4);
TASK_PP(16'h2EE4,4);
TASK_PP(16'h2EE5,4);
TASK_PP(16'h2EE6,4);
TASK_PP(16'h2EE7,4);
TASK_PP(16'h2EE8,4);
TASK_PP(16'h2EE9,4);
TASK_PP(16'h2EEA,4);
TASK_PP(16'h2EEB,4);
TASK_PP(16'h2EEC,4);
TASK_PP(16'h2EED,4);
TASK_PP(16'h2EEE,4);
TASK_PP(16'h2EEF,4);
TASK_PP(16'h2EF0,4);
TASK_PP(16'h2EF1,4);
TASK_PP(16'h2EF2,4);
TASK_PP(16'h2EF3,4);
TASK_PP(16'h2EF4,4);
TASK_PP(16'h2EF5,4);
TASK_PP(16'h2EF6,4);
TASK_PP(16'h2EF7,4);
TASK_PP(16'h2EF8,4);
TASK_PP(16'h2EF9,4);
TASK_PP(16'h2EFA,4);
TASK_PP(16'h2EFB,4);
TASK_PP(16'h2EFC,4);
TASK_PP(16'h2EFD,4);
TASK_PP(16'h2EFE,4);
TASK_PP(16'h2EFF,4);
TASK_PP(16'h2F00,4);
TASK_PP(16'h2F01,4);
TASK_PP(16'h2F02,4);
TASK_PP(16'h2F03,4);
TASK_PP(16'h2F04,4);
TASK_PP(16'h2F05,4);
TASK_PP(16'h2F06,4);
TASK_PP(16'h2F07,4);
TASK_PP(16'h2F08,4);
TASK_PP(16'h2F09,4);
TASK_PP(16'h2F0A,4);
TASK_PP(16'h2F0B,4);
TASK_PP(16'h2F0C,4);
TASK_PP(16'h2F0D,4);
TASK_PP(16'h2F0E,4);
TASK_PP(16'h2F0F,4);
TASK_PP(16'h2F10,4);
TASK_PP(16'h2F11,4);
TASK_PP(16'h2F12,4);
TASK_PP(16'h2F13,4);
TASK_PP(16'h2F14,4);
TASK_PP(16'h2F15,4);
TASK_PP(16'h2F16,4);
TASK_PP(16'h2F17,4);
TASK_PP(16'h2F18,4);
TASK_PP(16'h2F19,4);
TASK_PP(16'h2F1A,4);
TASK_PP(16'h2F1B,4);
TASK_PP(16'h2F1C,4);
TASK_PP(16'h2F1D,4);
TASK_PP(16'h2F1E,4);
TASK_PP(16'h2F1F,4);
TASK_PP(16'h2F20,4);
TASK_PP(16'h2F21,4);
TASK_PP(16'h2F22,4);
TASK_PP(16'h2F23,4);
TASK_PP(16'h2F24,4);
TASK_PP(16'h2F25,4);
TASK_PP(16'h2F26,4);
TASK_PP(16'h2F27,4);
TASK_PP(16'h2F28,4);
TASK_PP(16'h2F29,4);
TASK_PP(16'h2F2A,4);
TASK_PP(16'h2F2B,4);
TASK_PP(16'h2F2C,4);
TASK_PP(16'h2F2D,4);
TASK_PP(16'h2F2E,4);
TASK_PP(16'h2F2F,4);
TASK_PP(16'h2F30,4);
TASK_PP(16'h2F31,4);
TASK_PP(16'h2F32,4);
TASK_PP(16'h2F33,4);
TASK_PP(16'h2F34,4);
TASK_PP(16'h2F35,4);
TASK_PP(16'h2F36,4);
TASK_PP(16'h2F37,4);
TASK_PP(16'h2F38,4);
TASK_PP(16'h2F39,4);
TASK_PP(16'h2F3A,4);
TASK_PP(16'h2F3B,4);
TASK_PP(16'h2F3C,4);
TASK_PP(16'h2F3D,4);
TASK_PP(16'h2F3E,4);
TASK_PP(16'h2F3F,4);
TASK_PP(16'h2F40,4);
TASK_PP(16'h2F41,4);
TASK_PP(16'h2F42,4);
TASK_PP(16'h2F43,4);
TASK_PP(16'h2F44,4);
TASK_PP(16'h2F45,4);
TASK_PP(16'h2F46,4);
TASK_PP(16'h2F47,4);
TASK_PP(16'h2F48,4);
TASK_PP(16'h2F49,4);
TASK_PP(16'h2F4A,4);
TASK_PP(16'h2F4B,4);
TASK_PP(16'h2F4C,4);
TASK_PP(16'h2F4D,4);
TASK_PP(16'h2F4E,4);
TASK_PP(16'h2F4F,4);
TASK_PP(16'h2F50,4);
TASK_PP(16'h2F51,4);
TASK_PP(16'h2F52,4);
TASK_PP(16'h2F53,4);
TASK_PP(16'h2F54,4);
TASK_PP(16'h2F55,4);
TASK_PP(16'h2F56,4);
TASK_PP(16'h2F57,4);
TASK_PP(16'h2F58,4);
TASK_PP(16'h2F59,4);
TASK_PP(16'h2F5A,4);
TASK_PP(16'h2F5B,4);
TASK_PP(16'h2F5C,4);
TASK_PP(16'h2F5D,4);
TASK_PP(16'h2F5E,4);
TASK_PP(16'h2F5F,4);
TASK_PP(16'h2F60,4);
TASK_PP(16'h2F61,4);
TASK_PP(16'h2F62,4);
TASK_PP(16'h2F63,4);
TASK_PP(16'h2F64,4);
TASK_PP(16'h2F65,4);
TASK_PP(16'h2F66,4);
TASK_PP(16'h2F67,4);
TASK_PP(16'h2F68,4);
TASK_PP(16'h2F69,4);
TASK_PP(16'h2F6A,4);
TASK_PP(16'h2F6B,4);
TASK_PP(16'h2F6C,4);
TASK_PP(16'h2F6D,4);
TASK_PP(16'h2F6E,4);
TASK_PP(16'h2F6F,4);
TASK_PP(16'h2F70,4);
TASK_PP(16'h2F71,4);
TASK_PP(16'h2F72,4);
TASK_PP(16'h2F73,4);
TASK_PP(16'h2F74,4);
TASK_PP(16'h2F75,4);
TASK_PP(16'h2F76,4);
TASK_PP(16'h2F77,4);
TASK_PP(16'h2F78,4);
TASK_PP(16'h2F79,4);
TASK_PP(16'h2F7A,4);
TASK_PP(16'h2F7B,4);
TASK_PP(16'h2F7C,4);
TASK_PP(16'h2F7D,4);
TASK_PP(16'h2F7E,4);
TASK_PP(16'h2F7F,4);
TASK_PP(16'h2F80,4);
TASK_PP(16'h2F81,4);
TASK_PP(16'h2F82,4);
TASK_PP(16'h2F83,4);
TASK_PP(16'h2F84,4);
TASK_PP(16'h2F85,4);
TASK_PP(16'h2F86,4);
TASK_PP(16'h2F87,4);
TASK_PP(16'h2F88,4);
TASK_PP(16'h2F89,4);
TASK_PP(16'h2F8A,4);
TASK_PP(16'h2F8B,4);
TASK_PP(16'h2F8C,4);
TASK_PP(16'h2F8D,4);
TASK_PP(16'h2F8E,4);
TASK_PP(16'h2F8F,4);
TASK_PP(16'h2F90,4);
TASK_PP(16'h2F91,4);
TASK_PP(16'h2F92,4);
TASK_PP(16'h2F93,4);
TASK_PP(16'h2F94,4);
TASK_PP(16'h2F95,4);
TASK_PP(16'h2F96,4);
TASK_PP(16'h2F97,4);
TASK_PP(16'h2F98,4);
TASK_PP(16'h2F99,4);
TASK_PP(16'h2F9A,4);
TASK_PP(16'h2F9B,4);
TASK_PP(16'h2F9C,4);
TASK_PP(16'h2F9D,4);
TASK_PP(16'h2F9E,4);
TASK_PP(16'h2F9F,4);
TASK_PP(16'h2FA0,4);
TASK_PP(16'h2FA1,4);
TASK_PP(16'h2FA2,4);
TASK_PP(16'h2FA3,4);
TASK_PP(16'h2FA4,4);
TASK_PP(16'h2FA5,4);
TASK_PP(16'h2FA6,4);
TASK_PP(16'h2FA7,4);
TASK_PP(16'h2FA8,4);
TASK_PP(16'h2FA9,4);
TASK_PP(16'h2FAA,4);
TASK_PP(16'h2FAB,4);
TASK_PP(16'h2FAC,4);
TASK_PP(16'h2FAD,4);
TASK_PP(16'h2FAE,4);
TASK_PP(16'h2FAF,4);
TASK_PP(16'h2FB0,4);
TASK_PP(16'h2FB1,4);
TASK_PP(16'h2FB2,4);
TASK_PP(16'h2FB3,4);
TASK_PP(16'h2FB4,4);
TASK_PP(16'h2FB5,4);
TASK_PP(16'h2FB6,4);
TASK_PP(16'h2FB7,4);
TASK_PP(16'h2FB8,4);
TASK_PP(16'h2FB9,4);
TASK_PP(16'h2FBA,4);
TASK_PP(16'h2FBB,4);
TASK_PP(16'h2FBC,4);
TASK_PP(16'h2FBD,4);
TASK_PP(16'h2FBE,4);
TASK_PP(16'h2FBF,4);
TASK_PP(16'h2FC0,4);
TASK_PP(16'h2FC1,4);
TASK_PP(16'h2FC2,4);
TASK_PP(16'h2FC3,4);
TASK_PP(16'h2FC4,4);
TASK_PP(16'h2FC5,4);
TASK_PP(16'h2FC6,4);
TASK_PP(16'h2FC7,4);
TASK_PP(16'h2FC8,4);
TASK_PP(16'h2FC9,4);
TASK_PP(16'h2FCA,4);
TASK_PP(16'h2FCB,4);
TASK_PP(16'h2FCC,4);
TASK_PP(16'h2FCD,4);
TASK_PP(16'h2FCE,4);
TASK_PP(16'h2FCF,4);
TASK_PP(16'h2FD0,4);
TASK_PP(16'h2FD1,4);
TASK_PP(16'h2FD2,4);
TASK_PP(16'h2FD3,4);
TASK_PP(16'h2FD4,4);
TASK_PP(16'h2FD5,4);
TASK_PP(16'h2FD6,4);
TASK_PP(16'h2FD7,4);
TASK_PP(16'h2FD8,4);
TASK_PP(16'h2FD9,4);
TASK_PP(16'h2FDA,4);
TASK_PP(16'h2FDB,4);
TASK_PP(16'h2FDC,4);
TASK_PP(16'h2FDD,4);
TASK_PP(16'h2FDE,4);
TASK_PP(16'h2FDF,4);
TASK_PP(16'h2FE0,4);
TASK_PP(16'h2FE1,4);
TASK_PP(16'h2FE2,4);
TASK_PP(16'h2FE3,4);
TASK_PP(16'h2FE4,4);
TASK_PP(16'h2FE5,4);
TASK_PP(16'h2FE6,4);
TASK_PP(16'h2FE7,4);
TASK_PP(16'h2FE8,4);
TASK_PP(16'h2FE9,4);
TASK_PP(16'h2FEA,4);
TASK_PP(16'h2FEB,4);
TASK_PP(16'h2FEC,4);
TASK_PP(16'h2FED,4);
TASK_PP(16'h2FEE,4);
TASK_PP(16'h2FEF,4);
TASK_PP(16'h2FF0,4);
TASK_PP(16'h2FF1,4);
TASK_PP(16'h2FF2,4);
TASK_PP(16'h2FF3,4);
TASK_PP(16'h2FF4,4);
TASK_PP(16'h2FF5,4);
TASK_PP(16'h2FF6,4);
TASK_PP(16'h2FF7,4);
TASK_PP(16'h2FF8,4);
TASK_PP(16'h2FF9,4);
TASK_PP(16'h2FFA,4);
TASK_PP(16'h2FFB,4);
TASK_PP(16'h2FFC,4);
TASK_PP(16'h2FFD,4);
TASK_PP(16'h2FFE,4);
TASK_PP(16'h2FFF,4);
TASK_PP(16'h3000,4);
TASK_PP(16'h3001,4);
TASK_PP(16'h3002,4);
TASK_PP(16'h3003,4);
TASK_PP(16'h3004,4);
TASK_PP(16'h3005,4);
TASK_PP(16'h3006,4);
TASK_PP(16'h3007,4);
TASK_PP(16'h3008,4);
TASK_PP(16'h3009,4);
TASK_PP(16'h300A,4);
TASK_PP(16'h300B,4);
TASK_PP(16'h300C,4);
TASK_PP(16'h300D,4);
TASK_PP(16'h300E,4);
TASK_PP(16'h300F,4);
TASK_PP(16'h3010,4);
TASK_PP(16'h3011,4);
TASK_PP(16'h3012,4);
TASK_PP(16'h3013,4);
TASK_PP(16'h3014,4);
TASK_PP(16'h3015,4);
TASK_PP(16'h3016,4);
TASK_PP(16'h3017,4);
TASK_PP(16'h3018,4);
TASK_PP(16'h3019,4);
TASK_PP(16'h301A,4);
TASK_PP(16'h301B,4);
TASK_PP(16'h301C,4);
TASK_PP(16'h301D,4);
TASK_PP(16'h301E,4);
TASK_PP(16'h301F,4);
TASK_PP(16'h3020,4);
TASK_PP(16'h3021,4);
TASK_PP(16'h3022,4);
TASK_PP(16'h3023,4);
TASK_PP(16'h3024,4);
TASK_PP(16'h3025,4);
TASK_PP(16'h3026,4);
TASK_PP(16'h3027,4);
TASK_PP(16'h3028,4);
TASK_PP(16'h3029,4);
TASK_PP(16'h302A,4);
TASK_PP(16'h302B,4);
TASK_PP(16'h302C,4);
TASK_PP(16'h302D,4);
TASK_PP(16'h302E,4);
TASK_PP(16'h302F,4);
TASK_PP(16'h3030,4);
TASK_PP(16'h3031,4);
TASK_PP(16'h3032,4);
TASK_PP(16'h3033,4);
TASK_PP(16'h3034,4);
TASK_PP(16'h3035,4);
TASK_PP(16'h3036,4);
TASK_PP(16'h3037,4);
TASK_PP(16'h3038,4);
TASK_PP(16'h3039,4);
TASK_PP(16'h303A,4);
TASK_PP(16'h303B,4);
TASK_PP(16'h303C,4);
TASK_PP(16'h303D,4);
TASK_PP(16'h303E,4);
TASK_PP(16'h303F,4);
TASK_PP(16'h3040,4);
TASK_PP(16'h3041,4);
TASK_PP(16'h3042,4);
TASK_PP(16'h3043,4);
TASK_PP(16'h3044,4);
TASK_PP(16'h3045,4);
TASK_PP(16'h3046,4);
TASK_PP(16'h3047,4);
TASK_PP(16'h3048,4);
TASK_PP(16'h3049,4);
TASK_PP(16'h304A,4);
TASK_PP(16'h304B,4);
TASK_PP(16'h304C,4);
TASK_PP(16'h304D,4);
TASK_PP(16'h304E,4);
TASK_PP(16'h304F,4);
TASK_PP(16'h3050,4);
TASK_PP(16'h3051,4);
TASK_PP(16'h3052,4);
TASK_PP(16'h3053,4);
TASK_PP(16'h3054,4);
TASK_PP(16'h3055,4);
TASK_PP(16'h3056,4);
TASK_PP(16'h3057,4);
TASK_PP(16'h3058,4);
TASK_PP(16'h3059,4);
TASK_PP(16'h305A,4);
TASK_PP(16'h305B,4);
TASK_PP(16'h305C,4);
TASK_PP(16'h305D,4);
TASK_PP(16'h305E,4);
TASK_PP(16'h305F,4);
TASK_PP(16'h3060,4);
TASK_PP(16'h3061,4);
TASK_PP(16'h3062,4);
TASK_PP(16'h3063,4);
TASK_PP(16'h3064,4);
TASK_PP(16'h3065,4);
TASK_PP(16'h3066,4);
TASK_PP(16'h3067,4);
TASK_PP(16'h3068,4);
TASK_PP(16'h3069,4);
TASK_PP(16'h306A,4);
TASK_PP(16'h306B,4);
TASK_PP(16'h306C,4);
TASK_PP(16'h306D,4);
TASK_PP(16'h306E,4);
TASK_PP(16'h306F,4);
TASK_PP(16'h3070,4);
TASK_PP(16'h3071,4);
TASK_PP(16'h3072,4);
TASK_PP(16'h3073,4);
TASK_PP(16'h3074,4);
TASK_PP(16'h3075,4);
TASK_PP(16'h3076,4);
TASK_PP(16'h3077,4);
TASK_PP(16'h3078,4);
TASK_PP(16'h3079,4);
TASK_PP(16'h307A,4);
TASK_PP(16'h307B,4);
TASK_PP(16'h307C,4);
TASK_PP(16'h307D,4);
TASK_PP(16'h307E,4);
TASK_PP(16'h307F,4);
TASK_PP(16'h3080,4);
TASK_PP(16'h3081,4);
TASK_PP(16'h3082,4);
TASK_PP(16'h3083,4);
TASK_PP(16'h3084,4);
TASK_PP(16'h3085,4);
TASK_PP(16'h3086,4);
TASK_PP(16'h3087,4);
TASK_PP(16'h3088,4);
TASK_PP(16'h3089,4);
TASK_PP(16'h308A,4);
TASK_PP(16'h308B,4);
TASK_PP(16'h308C,4);
TASK_PP(16'h308D,4);
TASK_PP(16'h308E,4);
TASK_PP(16'h308F,4);
TASK_PP(16'h3090,4);
TASK_PP(16'h3091,4);
TASK_PP(16'h3092,4);
TASK_PP(16'h3093,4);
TASK_PP(16'h3094,4);
TASK_PP(16'h3095,4);
TASK_PP(16'h3096,4);
TASK_PP(16'h3097,4);
TASK_PP(16'h3098,4);
TASK_PP(16'h3099,4);
TASK_PP(16'h309A,4);
TASK_PP(16'h309B,4);
TASK_PP(16'h309C,4);
TASK_PP(16'h309D,4);
TASK_PP(16'h309E,4);
TASK_PP(16'h309F,4);
TASK_PP(16'h30A0,4);
TASK_PP(16'h30A1,4);
TASK_PP(16'h30A2,4);
TASK_PP(16'h30A3,4);
TASK_PP(16'h30A4,4);
TASK_PP(16'h30A5,4);
TASK_PP(16'h30A6,4);
TASK_PP(16'h30A7,4);
TASK_PP(16'h30A8,4);
TASK_PP(16'h30A9,4);
TASK_PP(16'h30AA,4);
TASK_PP(16'h30AB,4);
TASK_PP(16'h30AC,4);
TASK_PP(16'h30AD,4);
TASK_PP(16'h30AE,4);
TASK_PP(16'h30AF,4);
TASK_PP(16'h30B0,4);
TASK_PP(16'h30B1,4);
TASK_PP(16'h30B2,4);
TASK_PP(16'h30B3,4);
TASK_PP(16'h30B4,4);
TASK_PP(16'h30B5,4);
TASK_PP(16'h30B6,4);
TASK_PP(16'h30B7,4);
TASK_PP(16'h30B8,4);
TASK_PP(16'h30B9,4);
TASK_PP(16'h30BA,4);
TASK_PP(16'h30BB,4);
TASK_PP(16'h30BC,4);
TASK_PP(16'h30BD,4);
TASK_PP(16'h30BE,4);
TASK_PP(16'h30BF,4);
TASK_PP(16'h30C0,4);
TASK_PP(16'h30C1,4);
TASK_PP(16'h30C2,4);
TASK_PP(16'h30C3,4);
TASK_PP(16'h30C4,4);
TASK_PP(16'h30C5,4);
TASK_PP(16'h30C6,4);
TASK_PP(16'h30C7,4);
TASK_PP(16'h30C8,4);
TASK_PP(16'h30C9,4);
TASK_PP(16'h30CA,4);
TASK_PP(16'h30CB,4);
TASK_PP(16'h30CC,4);
TASK_PP(16'h30CD,4);
TASK_PP(16'h30CE,4);
TASK_PP(16'h30CF,4);
TASK_PP(16'h30D0,4);
TASK_PP(16'h30D1,4);
TASK_PP(16'h30D2,4);
TASK_PP(16'h30D3,4);
TASK_PP(16'h30D4,4);
TASK_PP(16'h30D5,4);
TASK_PP(16'h30D6,4);
TASK_PP(16'h30D7,4);
TASK_PP(16'h30D8,4);
TASK_PP(16'h30D9,4);
TASK_PP(16'h30DA,4);
TASK_PP(16'h30DB,4);
TASK_PP(16'h30DC,4);
TASK_PP(16'h30DD,4);
TASK_PP(16'h30DE,4);
TASK_PP(16'h30DF,4);
TASK_PP(16'h30E0,4);
TASK_PP(16'h30E1,4);
TASK_PP(16'h30E2,4);
TASK_PP(16'h30E3,4);
TASK_PP(16'h30E4,4);
TASK_PP(16'h30E5,4);
TASK_PP(16'h30E6,4);
TASK_PP(16'h30E7,4);
TASK_PP(16'h30E8,4);
TASK_PP(16'h30E9,4);
TASK_PP(16'h30EA,4);
TASK_PP(16'h30EB,4);
TASK_PP(16'h30EC,4);
TASK_PP(16'h30ED,4);
TASK_PP(16'h30EE,4);
TASK_PP(16'h30EF,4);
TASK_PP(16'h30F0,4);
TASK_PP(16'h30F1,4);
TASK_PP(16'h30F2,4);
TASK_PP(16'h30F3,4);
TASK_PP(16'h30F4,4);
TASK_PP(16'h30F5,4);
TASK_PP(16'h30F6,4);
TASK_PP(16'h30F7,4);
TASK_PP(16'h30F8,4);
TASK_PP(16'h30F9,4);
TASK_PP(16'h30FA,4);
TASK_PP(16'h30FB,4);
TASK_PP(16'h30FC,4);
TASK_PP(16'h30FD,4);
TASK_PP(16'h30FE,4);
TASK_PP(16'h30FF,4);
TASK_PP(16'h3100,4);
TASK_PP(16'h3101,4);
TASK_PP(16'h3102,4);
TASK_PP(16'h3103,4);
TASK_PP(16'h3104,4);
TASK_PP(16'h3105,4);
TASK_PP(16'h3106,4);
TASK_PP(16'h3107,4);
TASK_PP(16'h3108,4);
TASK_PP(16'h3109,4);
TASK_PP(16'h310A,4);
TASK_PP(16'h310B,4);
TASK_PP(16'h310C,4);
TASK_PP(16'h310D,4);
TASK_PP(16'h310E,4);
TASK_PP(16'h310F,4);
TASK_PP(16'h3110,4);
TASK_PP(16'h3111,4);
TASK_PP(16'h3112,4);
TASK_PP(16'h3113,4);
TASK_PP(16'h3114,4);
TASK_PP(16'h3115,4);
TASK_PP(16'h3116,4);
TASK_PP(16'h3117,4);
TASK_PP(16'h3118,4);
TASK_PP(16'h3119,4);
TASK_PP(16'h311A,4);
TASK_PP(16'h311B,4);
TASK_PP(16'h311C,4);
TASK_PP(16'h311D,4);
TASK_PP(16'h311E,4);
TASK_PP(16'h311F,4);
TASK_PP(16'h3120,4);
TASK_PP(16'h3121,4);
TASK_PP(16'h3122,4);
TASK_PP(16'h3123,4);
TASK_PP(16'h3124,4);
TASK_PP(16'h3125,4);
TASK_PP(16'h3126,4);
TASK_PP(16'h3127,4);
TASK_PP(16'h3128,4);
TASK_PP(16'h3129,4);
TASK_PP(16'h312A,4);
TASK_PP(16'h312B,4);
TASK_PP(16'h312C,4);
TASK_PP(16'h312D,4);
TASK_PP(16'h312E,4);
TASK_PP(16'h312F,4);
TASK_PP(16'h3130,4);
TASK_PP(16'h3131,4);
TASK_PP(16'h3132,4);
TASK_PP(16'h3133,4);
TASK_PP(16'h3134,4);
TASK_PP(16'h3135,4);
TASK_PP(16'h3136,4);
TASK_PP(16'h3137,4);
TASK_PP(16'h3138,4);
TASK_PP(16'h3139,4);
TASK_PP(16'h313A,4);
TASK_PP(16'h313B,4);
TASK_PP(16'h313C,4);
TASK_PP(16'h313D,4);
TASK_PP(16'h313E,4);
TASK_PP(16'h313F,4);
TASK_PP(16'h3140,4);
TASK_PP(16'h3141,4);
TASK_PP(16'h3142,4);
TASK_PP(16'h3143,4);
TASK_PP(16'h3144,4);
TASK_PP(16'h3145,4);
TASK_PP(16'h3146,4);
TASK_PP(16'h3147,4);
TASK_PP(16'h3148,4);
TASK_PP(16'h3149,4);
TASK_PP(16'h314A,4);
TASK_PP(16'h314B,4);
TASK_PP(16'h314C,4);
TASK_PP(16'h314D,4);
TASK_PP(16'h314E,4);
TASK_PP(16'h314F,4);
TASK_PP(16'h3150,4);
TASK_PP(16'h3151,4);
TASK_PP(16'h3152,4);
TASK_PP(16'h3153,4);
TASK_PP(16'h3154,4);
TASK_PP(16'h3155,4);
TASK_PP(16'h3156,4);
TASK_PP(16'h3157,4);
TASK_PP(16'h3158,4);
TASK_PP(16'h3159,4);
TASK_PP(16'h315A,4);
TASK_PP(16'h315B,4);
TASK_PP(16'h315C,4);
TASK_PP(16'h315D,4);
TASK_PP(16'h315E,4);
TASK_PP(16'h315F,4);
TASK_PP(16'h3160,4);
TASK_PP(16'h3161,4);
TASK_PP(16'h3162,4);
TASK_PP(16'h3163,4);
TASK_PP(16'h3164,4);
TASK_PP(16'h3165,4);
TASK_PP(16'h3166,4);
TASK_PP(16'h3167,4);
TASK_PP(16'h3168,4);
TASK_PP(16'h3169,4);
TASK_PP(16'h316A,4);
TASK_PP(16'h316B,4);
TASK_PP(16'h316C,4);
TASK_PP(16'h316D,4);
TASK_PP(16'h316E,4);
TASK_PP(16'h316F,4);
TASK_PP(16'h3170,4);
TASK_PP(16'h3171,4);
TASK_PP(16'h3172,4);
TASK_PP(16'h3173,4);
TASK_PP(16'h3174,4);
TASK_PP(16'h3175,4);
TASK_PP(16'h3176,4);
TASK_PP(16'h3177,4);
TASK_PP(16'h3178,4);
TASK_PP(16'h3179,4);
TASK_PP(16'h317A,4);
TASK_PP(16'h317B,4);
TASK_PP(16'h317C,4);
TASK_PP(16'h317D,4);
TASK_PP(16'h317E,4);
TASK_PP(16'h317F,4);
TASK_PP(16'h3180,4);
TASK_PP(16'h3181,4);
TASK_PP(16'h3182,4);
TASK_PP(16'h3183,4);
TASK_PP(16'h3184,4);
TASK_PP(16'h3185,4);
TASK_PP(16'h3186,4);
TASK_PP(16'h3187,4);
TASK_PP(16'h3188,4);
TASK_PP(16'h3189,4);
TASK_PP(16'h318A,4);
TASK_PP(16'h318B,4);
TASK_PP(16'h318C,4);
TASK_PP(16'h318D,4);
TASK_PP(16'h318E,4);
TASK_PP(16'h318F,4);
TASK_PP(16'h3190,4);
TASK_PP(16'h3191,4);
TASK_PP(16'h3192,4);
TASK_PP(16'h3193,4);
TASK_PP(16'h3194,4);
TASK_PP(16'h3195,4);
TASK_PP(16'h3196,4);
TASK_PP(16'h3197,4);
TASK_PP(16'h3198,4);
TASK_PP(16'h3199,4);
TASK_PP(16'h319A,4);
TASK_PP(16'h319B,4);
TASK_PP(16'h319C,4);
TASK_PP(16'h319D,4);
TASK_PP(16'h319E,4);
TASK_PP(16'h319F,4);
TASK_PP(16'h31A0,4);
TASK_PP(16'h31A1,4);
TASK_PP(16'h31A2,4);
TASK_PP(16'h31A3,4);
TASK_PP(16'h31A4,4);
TASK_PP(16'h31A5,4);
TASK_PP(16'h31A6,4);
TASK_PP(16'h31A7,4);
TASK_PP(16'h31A8,4);
TASK_PP(16'h31A9,4);
TASK_PP(16'h31AA,4);
TASK_PP(16'h31AB,4);
TASK_PP(16'h31AC,4);
TASK_PP(16'h31AD,4);
TASK_PP(16'h31AE,4);
TASK_PP(16'h31AF,4);
TASK_PP(16'h31B0,4);
TASK_PP(16'h31B1,4);
TASK_PP(16'h31B2,4);
TASK_PP(16'h31B3,4);
TASK_PP(16'h31B4,4);
TASK_PP(16'h31B5,4);
TASK_PP(16'h31B6,4);
TASK_PP(16'h31B7,4);
TASK_PP(16'h31B8,4);
TASK_PP(16'h31B9,4);
TASK_PP(16'h31BA,4);
TASK_PP(16'h31BB,4);
TASK_PP(16'h31BC,4);
TASK_PP(16'h31BD,4);
TASK_PP(16'h31BE,4);
TASK_PP(16'h31BF,4);
TASK_PP(16'h31C0,4);
TASK_PP(16'h31C1,4);
TASK_PP(16'h31C2,4);
TASK_PP(16'h31C3,4);
TASK_PP(16'h31C4,4);
TASK_PP(16'h31C5,4);
TASK_PP(16'h31C6,4);
TASK_PP(16'h31C7,4);
TASK_PP(16'h31C8,4);
TASK_PP(16'h31C9,4);
TASK_PP(16'h31CA,4);
TASK_PP(16'h31CB,4);
TASK_PP(16'h31CC,4);
TASK_PP(16'h31CD,4);
TASK_PP(16'h31CE,4);
TASK_PP(16'h31CF,4);
TASK_PP(16'h31D0,4);
TASK_PP(16'h31D1,4);
TASK_PP(16'h31D2,4);
TASK_PP(16'h31D3,4);
TASK_PP(16'h31D4,4);
TASK_PP(16'h31D5,4);
TASK_PP(16'h31D6,4);
TASK_PP(16'h31D7,4);
TASK_PP(16'h31D8,4);
TASK_PP(16'h31D9,4);
TASK_PP(16'h31DA,4);
TASK_PP(16'h31DB,4);
TASK_PP(16'h31DC,4);
TASK_PP(16'h31DD,4);
TASK_PP(16'h31DE,4);
TASK_PP(16'h31DF,4);
TASK_PP(16'h31E0,4);
TASK_PP(16'h31E1,4);
TASK_PP(16'h31E2,4);
TASK_PP(16'h31E3,4);
TASK_PP(16'h31E4,4);
TASK_PP(16'h31E5,4);
TASK_PP(16'h31E6,4);
TASK_PP(16'h31E7,4);
TASK_PP(16'h31E8,4);
TASK_PP(16'h31E9,4);
TASK_PP(16'h31EA,4);
TASK_PP(16'h31EB,4);
TASK_PP(16'h31EC,4);
TASK_PP(16'h31ED,4);
TASK_PP(16'h31EE,4);
TASK_PP(16'h31EF,4);
TASK_PP(16'h31F0,4);
TASK_PP(16'h31F1,4);
TASK_PP(16'h31F2,4);
TASK_PP(16'h31F3,4);
TASK_PP(16'h31F4,4);
TASK_PP(16'h31F5,4);
TASK_PP(16'h31F6,4);
TASK_PP(16'h31F7,4);
TASK_PP(16'h31F8,4);
TASK_PP(16'h31F9,4);
TASK_PP(16'h31FA,4);
TASK_PP(16'h31FB,4);
TASK_PP(16'h31FC,4);
TASK_PP(16'h31FD,4);
TASK_PP(16'h31FE,4);
TASK_PP(16'h31FF,4);
TASK_PP(16'h3200,4);
TASK_PP(16'h3201,4);
TASK_PP(16'h3202,4);
TASK_PP(16'h3203,4);
TASK_PP(16'h3204,4);
TASK_PP(16'h3205,4);
TASK_PP(16'h3206,4);
TASK_PP(16'h3207,4);
TASK_PP(16'h3208,4);
TASK_PP(16'h3209,4);
TASK_PP(16'h320A,4);
TASK_PP(16'h320B,4);
TASK_PP(16'h320C,4);
TASK_PP(16'h320D,4);
TASK_PP(16'h320E,4);
TASK_PP(16'h320F,4);
TASK_PP(16'h3210,4);
TASK_PP(16'h3211,4);
TASK_PP(16'h3212,4);
TASK_PP(16'h3213,4);
TASK_PP(16'h3214,4);
TASK_PP(16'h3215,4);
TASK_PP(16'h3216,4);
TASK_PP(16'h3217,4);
TASK_PP(16'h3218,4);
TASK_PP(16'h3219,4);
TASK_PP(16'h321A,4);
TASK_PP(16'h321B,4);
TASK_PP(16'h321C,4);
TASK_PP(16'h321D,4);
TASK_PP(16'h321E,4);
TASK_PP(16'h321F,4);
TASK_PP(16'h3220,4);
TASK_PP(16'h3221,4);
TASK_PP(16'h3222,4);
TASK_PP(16'h3223,4);
TASK_PP(16'h3224,4);
TASK_PP(16'h3225,4);
TASK_PP(16'h3226,4);
TASK_PP(16'h3227,4);
TASK_PP(16'h3228,4);
TASK_PP(16'h3229,4);
TASK_PP(16'h322A,4);
TASK_PP(16'h322B,4);
TASK_PP(16'h322C,4);
TASK_PP(16'h322D,4);
TASK_PP(16'h322E,4);
TASK_PP(16'h322F,4);
TASK_PP(16'h3230,4);
TASK_PP(16'h3231,4);
TASK_PP(16'h3232,4);
TASK_PP(16'h3233,4);
TASK_PP(16'h3234,4);
TASK_PP(16'h3235,4);
TASK_PP(16'h3236,4);
TASK_PP(16'h3237,4);
TASK_PP(16'h3238,4);
TASK_PP(16'h3239,4);
TASK_PP(16'h323A,4);
TASK_PP(16'h323B,4);
TASK_PP(16'h323C,4);
TASK_PP(16'h323D,4);
TASK_PP(16'h323E,4);
TASK_PP(16'h323F,4);
TASK_PP(16'h3240,4);
TASK_PP(16'h3241,4);
TASK_PP(16'h3242,4);
TASK_PP(16'h3243,4);
TASK_PP(16'h3244,4);
TASK_PP(16'h3245,4);
TASK_PP(16'h3246,4);
TASK_PP(16'h3247,4);
TASK_PP(16'h3248,4);
TASK_PP(16'h3249,4);
TASK_PP(16'h324A,4);
TASK_PP(16'h324B,4);
TASK_PP(16'h324C,4);
TASK_PP(16'h324D,4);
TASK_PP(16'h324E,4);
TASK_PP(16'h324F,4);
TASK_PP(16'h3250,4);
TASK_PP(16'h3251,4);
TASK_PP(16'h3252,4);
TASK_PP(16'h3253,4);
TASK_PP(16'h3254,4);
TASK_PP(16'h3255,4);
TASK_PP(16'h3256,4);
TASK_PP(16'h3257,4);
TASK_PP(16'h3258,4);
TASK_PP(16'h3259,4);
TASK_PP(16'h325A,4);
TASK_PP(16'h325B,4);
TASK_PP(16'h325C,4);
TASK_PP(16'h325D,4);
TASK_PP(16'h325E,4);
TASK_PP(16'h325F,4);
TASK_PP(16'h3260,4);
TASK_PP(16'h3261,4);
TASK_PP(16'h3262,4);
TASK_PP(16'h3263,4);
TASK_PP(16'h3264,4);
TASK_PP(16'h3265,4);
TASK_PP(16'h3266,4);
TASK_PP(16'h3267,4);
TASK_PP(16'h3268,4);
TASK_PP(16'h3269,4);
TASK_PP(16'h326A,4);
TASK_PP(16'h326B,4);
TASK_PP(16'h326C,4);
TASK_PP(16'h326D,4);
TASK_PP(16'h326E,4);
TASK_PP(16'h326F,4);
TASK_PP(16'h3270,4);
TASK_PP(16'h3271,4);
TASK_PP(16'h3272,4);
TASK_PP(16'h3273,4);
TASK_PP(16'h3274,4);
TASK_PP(16'h3275,4);
TASK_PP(16'h3276,4);
TASK_PP(16'h3277,4);
TASK_PP(16'h3278,4);
TASK_PP(16'h3279,4);
TASK_PP(16'h327A,4);
TASK_PP(16'h327B,4);
TASK_PP(16'h327C,4);
TASK_PP(16'h327D,4);
TASK_PP(16'h327E,4);
TASK_PP(16'h327F,4);
TASK_PP(16'h3280,4);
TASK_PP(16'h3281,4);
TASK_PP(16'h3282,4);
TASK_PP(16'h3283,4);
TASK_PP(16'h3284,4);
TASK_PP(16'h3285,4);
TASK_PP(16'h3286,4);
TASK_PP(16'h3287,4);
TASK_PP(16'h3288,4);
TASK_PP(16'h3289,4);
TASK_PP(16'h328A,4);
TASK_PP(16'h328B,4);
TASK_PP(16'h328C,4);
TASK_PP(16'h328D,4);
TASK_PP(16'h328E,4);
TASK_PP(16'h328F,4);
TASK_PP(16'h3290,4);
TASK_PP(16'h3291,4);
TASK_PP(16'h3292,4);
TASK_PP(16'h3293,4);
TASK_PP(16'h3294,4);
TASK_PP(16'h3295,4);
TASK_PP(16'h3296,4);
TASK_PP(16'h3297,4);
TASK_PP(16'h3298,4);
TASK_PP(16'h3299,4);
TASK_PP(16'h329A,4);
TASK_PP(16'h329B,4);
TASK_PP(16'h329C,4);
TASK_PP(16'h329D,4);
TASK_PP(16'h329E,4);
TASK_PP(16'h329F,4);
TASK_PP(16'h32A0,4);
TASK_PP(16'h32A1,4);
TASK_PP(16'h32A2,4);
TASK_PP(16'h32A3,4);
TASK_PP(16'h32A4,4);
TASK_PP(16'h32A5,4);
TASK_PP(16'h32A6,4);
TASK_PP(16'h32A7,4);
TASK_PP(16'h32A8,4);
TASK_PP(16'h32A9,4);
TASK_PP(16'h32AA,4);
TASK_PP(16'h32AB,4);
TASK_PP(16'h32AC,4);
TASK_PP(16'h32AD,4);
TASK_PP(16'h32AE,4);
TASK_PP(16'h32AF,4);
TASK_PP(16'h32B0,4);
TASK_PP(16'h32B1,4);
TASK_PP(16'h32B2,4);
TASK_PP(16'h32B3,4);
TASK_PP(16'h32B4,4);
TASK_PP(16'h32B5,4);
TASK_PP(16'h32B6,4);
TASK_PP(16'h32B7,4);
TASK_PP(16'h32B8,4);
TASK_PP(16'h32B9,4);
TASK_PP(16'h32BA,4);
TASK_PP(16'h32BB,4);
TASK_PP(16'h32BC,4);
TASK_PP(16'h32BD,4);
TASK_PP(16'h32BE,4);
TASK_PP(16'h32BF,4);
TASK_PP(16'h32C0,4);
TASK_PP(16'h32C1,4);
TASK_PP(16'h32C2,4);
TASK_PP(16'h32C3,4);
TASK_PP(16'h32C4,4);
TASK_PP(16'h32C5,4);
TASK_PP(16'h32C6,4);
TASK_PP(16'h32C7,4);
TASK_PP(16'h32C8,4);
TASK_PP(16'h32C9,4);
TASK_PP(16'h32CA,4);
TASK_PP(16'h32CB,4);
TASK_PP(16'h32CC,4);
TASK_PP(16'h32CD,4);
TASK_PP(16'h32CE,4);
TASK_PP(16'h32CF,4);
TASK_PP(16'h32D0,4);
TASK_PP(16'h32D1,4);
TASK_PP(16'h32D2,4);
TASK_PP(16'h32D3,4);
TASK_PP(16'h32D4,4);
TASK_PP(16'h32D5,4);
TASK_PP(16'h32D6,4);
TASK_PP(16'h32D7,4);
TASK_PP(16'h32D8,4);
TASK_PP(16'h32D9,4);
TASK_PP(16'h32DA,4);
TASK_PP(16'h32DB,4);
TASK_PP(16'h32DC,4);
TASK_PP(16'h32DD,4);
TASK_PP(16'h32DE,4);
TASK_PP(16'h32DF,4);
TASK_PP(16'h32E0,4);
TASK_PP(16'h32E1,4);
TASK_PP(16'h32E2,4);
TASK_PP(16'h32E3,4);
TASK_PP(16'h32E4,4);
TASK_PP(16'h32E5,4);
TASK_PP(16'h32E6,4);
TASK_PP(16'h32E7,4);
TASK_PP(16'h32E8,4);
TASK_PP(16'h32E9,4);
TASK_PP(16'h32EA,4);
TASK_PP(16'h32EB,4);
TASK_PP(16'h32EC,4);
TASK_PP(16'h32ED,4);
TASK_PP(16'h32EE,4);
TASK_PP(16'h32EF,4);
TASK_PP(16'h32F0,4);
TASK_PP(16'h32F1,4);
TASK_PP(16'h32F2,4);
TASK_PP(16'h32F3,4);
TASK_PP(16'h32F4,4);
TASK_PP(16'h32F5,4);
TASK_PP(16'h32F6,4);
TASK_PP(16'h32F7,4);
TASK_PP(16'h32F8,4);
TASK_PP(16'h32F9,4);
TASK_PP(16'h32FA,4);
TASK_PP(16'h32FB,4);
TASK_PP(16'h32FC,4);
TASK_PP(16'h32FD,4);
TASK_PP(16'h32FE,4);
TASK_PP(16'h32FF,4);
TASK_PP(16'h3300,4);
TASK_PP(16'h3301,4);
TASK_PP(16'h3302,4);
TASK_PP(16'h3303,4);
TASK_PP(16'h3304,4);
TASK_PP(16'h3305,4);
TASK_PP(16'h3306,4);
TASK_PP(16'h3307,4);
TASK_PP(16'h3308,4);
TASK_PP(16'h3309,4);
TASK_PP(16'h330A,4);
TASK_PP(16'h330B,4);
TASK_PP(16'h330C,4);
TASK_PP(16'h330D,4);
TASK_PP(16'h330E,4);
TASK_PP(16'h330F,4);
TASK_PP(16'h3310,4);
TASK_PP(16'h3311,4);
TASK_PP(16'h3312,4);
TASK_PP(16'h3313,4);
TASK_PP(16'h3314,4);
TASK_PP(16'h3315,4);
TASK_PP(16'h3316,4);
TASK_PP(16'h3317,4);
TASK_PP(16'h3318,4);
TASK_PP(16'h3319,4);
TASK_PP(16'h331A,4);
TASK_PP(16'h331B,4);
TASK_PP(16'h331C,4);
TASK_PP(16'h331D,4);
TASK_PP(16'h331E,4);
TASK_PP(16'h331F,4);
TASK_PP(16'h3320,4);
TASK_PP(16'h3321,4);
TASK_PP(16'h3322,4);
TASK_PP(16'h3323,4);
TASK_PP(16'h3324,4);
TASK_PP(16'h3325,4);
TASK_PP(16'h3326,4);
TASK_PP(16'h3327,4);
TASK_PP(16'h3328,4);
TASK_PP(16'h3329,4);
TASK_PP(16'h332A,4);
TASK_PP(16'h332B,4);
TASK_PP(16'h332C,4);
TASK_PP(16'h332D,4);
TASK_PP(16'h332E,4);
TASK_PP(16'h332F,4);
TASK_PP(16'h3330,4);
TASK_PP(16'h3331,4);
TASK_PP(16'h3332,4);
TASK_PP(16'h3333,4);
TASK_PP(16'h3334,4);
TASK_PP(16'h3335,4);
TASK_PP(16'h3336,4);
TASK_PP(16'h3337,4);
TASK_PP(16'h3338,4);
TASK_PP(16'h3339,4);
TASK_PP(16'h333A,4);
TASK_PP(16'h333B,4);
TASK_PP(16'h333C,4);
TASK_PP(16'h333D,4);
TASK_PP(16'h333E,4);
TASK_PP(16'h333F,4);
TASK_PP(16'h3340,4);
TASK_PP(16'h3341,4);
TASK_PP(16'h3342,4);
TASK_PP(16'h3343,4);
TASK_PP(16'h3344,4);
TASK_PP(16'h3345,4);
TASK_PP(16'h3346,4);
TASK_PP(16'h3347,4);
TASK_PP(16'h3348,4);
TASK_PP(16'h3349,4);
TASK_PP(16'h334A,4);
TASK_PP(16'h334B,4);
TASK_PP(16'h334C,4);
TASK_PP(16'h334D,4);
TASK_PP(16'h334E,4);
TASK_PP(16'h334F,4);
TASK_PP(16'h3350,4);
TASK_PP(16'h3351,4);
TASK_PP(16'h3352,4);
TASK_PP(16'h3353,4);
TASK_PP(16'h3354,4);
TASK_PP(16'h3355,4);
TASK_PP(16'h3356,4);
TASK_PP(16'h3357,4);
TASK_PP(16'h3358,4);
TASK_PP(16'h3359,4);
TASK_PP(16'h335A,4);
TASK_PP(16'h335B,4);
TASK_PP(16'h335C,4);
TASK_PP(16'h335D,4);
TASK_PP(16'h335E,4);
TASK_PP(16'h335F,4);
TASK_PP(16'h3360,4);
TASK_PP(16'h3361,4);
TASK_PP(16'h3362,4);
TASK_PP(16'h3363,4);
TASK_PP(16'h3364,4);
TASK_PP(16'h3365,4);
TASK_PP(16'h3366,4);
TASK_PP(16'h3367,4);
TASK_PP(16'h3368,4);
TASK_PP(16'h3369,4);
TASK_PP(16'h336A,4);
TASK_PP(16'h336B,4);
TASK_PP(16'h336C,4);
TASK_PP(16'h336D,4);
TASK_PP(16'h336E,4);
TASK_PP(16'h336F,4);
TASK_PP(16'h3370,4);
TASK_PP(16'h3371,4);
TASK_PP(16'h3372,4);
TASK_PP(16'h3373,4);
TASK_PP(16'h3374,4);
TASK_PP(16'h3375,4);
TASK_PP(16'h3376,4);
TASK_PP(16'h3377,4);
TASK_PP(16'h3378,4);
TASK_PP(16'h3379,4);
TASK_PP(16'h337A,4);
TASK_PP(16'h337B,4);
TASK_PP(16'h337C,4);
TASK_PP(16'h337D,4);
TASK_PP(16'h337E,4);
TASK_PP(16'h337F,4);
TASK_PP(16'h3380,4);
TASK_PP(16'h3381,4);
TASK_PP(16'h3382,4);
TASK_PP(16'h3383,4);
TASK_PP(16'h3384,4);
TASK_PP(16'h3385,4);
TASK_PP(16'h3386,4);
TASK_PP(16'h3387,4);
TASK_PP(16'h3388,4);
TASK_PP(16'h3389,4);
TASK_PP(16'h338A,4);
TASK_PP(16'h338B,4);
TASK_PP(16'h338C,4);
TASK_PP(16'h338D,4);
TASK_PP(16'h338E,4);
TASK_PP(16'h338F,4);
TASK_PP(16'h3390,4);
TASK_PP(16'h3391,4);
TASK_PP(16'h3392,4);
TASK_PP(16'h3393,4);
TASK_PP(16'h3394,4);
TASK_PP(16'h3395,4);
TASK_PP(16'h3396,4);
TASK_PP(16'h3397,4);
TASK_PP(16'h3398,4);
TASK_PP(16'h3399,4);
TASK_PP(16'h339A,4);
TASK_PP(16'h339B,4);
TASK_PP(16'h339C,4);
TASK_PP(16'h339D,4);
TASK_PP(16'h339E,4);
TASK_PP(16'h339F,4);
TASK_PP(16'h33A0,4);
TASK_PP(16'h33A1,4);
TASK_PP(16'h33A2,4);
TASK_PP(16'h33A3,4);
TASK_PP(16'h33A4,4);
TASK_PP(16'h33A5,4);
TASK_PP(16'h33A6,4);
TASK_PP(16'h33A7,4);
TASK_PP(16'h33A8,4);
TASK_PP(16'h33A9,4);
TASK_PP(16'h33AA,4);
TASK_PP(16'h33AB,4);
TASK_PP(16'h33AC,4);
TASK_PP(16'h33AD,4);
TASK_PP(16'h33AE,4);
TASK_PP(16'h33AF,4);
TASK_PP(16'h33B0,4);
TASK_PP(16'h33B1,4);
TASK_PP(16'h33B2,4);
TASK_PP(16'h33B3,4);
TASK_PP(16'h33B4,4);
TASK_PP(16'h33B5,4);
TASK_PP(16'h33B6,4);
TASK_PP(16'h33B7,4);
TASK_PP(16'h33B8,4);
TASK_PP(16'h33B9,4);
TASK_PP(16'h33BA,4);
TASK_PP(16'h33BB,4);
TASK_PP(16'h33BC,4);
TASK_PP(16'h33BD,4);
TASK_PP(16'h33BE,4);
TASK_PP(16'h33BF,4);
TASK_PP(16'h33C0,4);
TASK_PP(16'h33C1,4);
TASK_PP(16'h33C2,4);
TASK_PP(16'h33C3,4);
TASK_PP(16'h33C4,4);
TASK_PP(16'h33C5,4);
TASK_PP(16'h33C6,4);
TASK_PP(16'h33C7,4);
TASK_PP(16'h33C8,4);
TASK_PP(16'h33C9,4);
TASK_PP(16'h33CA,4);
TASK_PP(16'h33CB,4);
TASK_PP(16'h33CC,4);
TASK_PP(16'h33CD,4);
TASK_PP(16'h33CE,4);
TASK_PP(16'h33CF,4);
TASK_PP(16'h33D0,4);
TASK_PP(16'h33D1,4);
TASK_PP(16'h33D2,4);
TASK_PP(16'h33D3,4);
TASK_PP(16'h33D4,4);
TASK_PP(16'h33D5,4);
TASK_PP(16'h33D6,4);
TASK_PP(16'h33D7,4);
TASK_PP(16'h33D8,4);
TASK_PP(16'h33D9,4);
TASK_PP(16'h33DA,4);
TASK_PP(16'h33DB,4);
TASK_PP(16'h33DC,4);
TASK_PP(16'h33DD,4);
TASK_PP(16'h33DE,4);
TASK_PP(16'h33DF,4);
TASK_PP(16'h33E0,4);
TASK_PP(16'h33E1,4);
TASK_PP(16'h33E2,4);
TASK_PP(16'h33E3,4);
TASK_PP(16'h33E4,4);
TASK_PP(16'h33E5,4);
TASK_PP(16'h33E6,4);
TASK_PP(16'h33E7,4);
TASK_PP(16'h33E8,4);
TASK_PP(16'h33E9,4);
TASK_PP(16'h33EA,4);
TASK_PP(16'h33EB,4);
TASK_PP(16'h33EC,4);
TASK_PP(16'h33ED,4);
TASK_PP(16'h33EE,4);
TASK_PP(16'h33EF,4);
TASK_PP(16'h33F0,4);
TASK_PP(16'h33F1,4);
TASK_PP(16'h33F2,4);
TASK_PP(16'h33F3,4);
TASK_PP(16'h33F4,4);
TASK_PP(16'h33F5,4);
TASK_PP(16'h33F6,4);
TASK_PP(16'h33F7,4);
TASK_PP(16'h33F8,4);
TASK_PP(16'h33F9,4);
TASK_PP(16'h33FA,4);
TASK_PP(16'h33FB,4);
TASK_PP(16'h33FC,4);
TASK_PP(16'h33FD,4);
TASK_PP(16'h33FE,4);
TASK_PP(16'h33FF,4);
TASK_PP(16'h3400,4);
TASK_PP(16'h3401,4);
TASK_PP(16'h3402,4);
TASK_PP(16'h3403,4);
TASK_PP(16'h3404,4);
TASK_PP(16'h3405,4);
TASK_PP(16'h3406,4);
TASK_PP(16'h3407,4);
TASK_PP(16'h3408,4);
TASK_PP(16'h3409,4);
TASK_PP(16'h340A,4);
TASK_PP(16'h340B,4);
TASK_PP(16'h340C,4);
TASK_PP(16'h340D,4);
TASK_PP(16'h340E,4);
TASK_PP(16'h340F,4);
TASK_PP(16'h3410,4);
TASK_PP(16'h3411,4);
TASK_PP(16'h3412,4);
TASK_PP(16'h3413,4);
TASK_PP(16'h3414,4);
TASK_PP(16'h3415,4);
TASK_PP(16'h3416,4);
TASK_PP(16'h3417,4);
TASK_PP(16'h3418,4);
TASK_PP(16'h3419,4);
TASK_PP(16'h341A,4);
TASK_PP(16'h341B,4);
TASK_PP(16'h341C,4);
TASK_PP(16'h341D,4);
TASK_PP(16'h341E,4);
TASK_PP(16'h341F,4);
TASK_PP(16'h3420,4);
TASK_PP(16'h3421,4);
TASK_PP(16'h3422,4);
TASK_PP(16'h3423,4);
TASK_PP(16'h3424,4);
TASK_PP(16'h3425,4);
TASK_PP(16'h3426,4);
TASK_PP(16'h3427,4);
TASK_PP(16'h3428,4);
TASK_PP(16'h3429,4);
TASK_PP(16'h342A,4);
TASK_PP(16'h342B,4);
TASK_PP(16'h342C,4);
TASK_PP(16'h342D,4);
TASK_PP(16'h342E,4);
TASK_PP(16'h342F,4);
TASK_PP(16'h3430,4);
TASK_PP(16'h3431,4);
TASK_PP(16'h3432,4);
TASK_PP(16'h3433,4);
TASK_PP(16'h3434,4);
TASK_PP(16'h3435,4);
TASK_PP(16'h3436,4);
TASK_PP(16'h3437,4);
TASK_PP(16'h3438,4);
TASK_PP(16'h3439,4);
TASK_PP(16'h343A,4);
TASK_PP(16'h343B,4);
TASK_PP(16'h343C,4);
TASK_PP(16'h343D,4);
TASK_PP(16'h343E,4);
TASK_PP(16'h343F,4);
TASK_PP(16'h3440,4);
TASK_PP(16'h3441,4);
TASK_PP(16'h3442,4);
TASK_PP(16'h3443,4);
TASK_PP(16'h3444,4);
TASK_PP(16'h3445,4);
TASK_PP(16'h3446,4);
TASK_PP(16'h3447,4);
TASK_PP(16'h3448,4);
TASK_PP(16'h3449,4);
TASK_PP(16'h344A,4);
TASK_PP(16'h344B,4);
TASK_PP(16'h344C,4);
TASK_PP(16'h344D,4);
TASK_PP(16'h344E,4);
TASK_PP(16'h344F,4);
TASK_PP(16'h3450,4);
TASK_PP(16'h3451,4);
TASK_PP(16'h3452,4);
TASK_PP(16'h3453,4);
TASK_PP(16'h3454,4);
TASK_PP(16'h3455,4);
TASK_PP(16'h3456,4);
TASK_PP(16'h3457,4);
TASK_PP(16'h3458,4);
TASK_PP(16'h3459,4);
TASK_PP(16'h345A,4);
TASK_PP(16'h345B,4);
TASK_PP(16'h345C,4);
TASK_PP(16'h345D,4);
TASK_PP(16'h345E,4);
TASK_PP(16'h345F,4);
TASK_PP(16'h3460,4);
TASK_PP(16'h3461,4);
TASK_PP(16'h3462,4);
TASK_PP(16'h3463,4);
TASK_PP(16'h3464,4);
TASK_PP(16'h3465,4);
TASK_PP(16'h3466,4);
TASK_PP(16'h3467,4);
TASK_PP(16'h3468,4);
TASK_PP(16'h3469,4);
TASK_PP(16'h346A,4);
TASK_PP(16'h346B,4);
TASK_PP(16'h346C,4);
TASK_PP(16'h346D,4);
TASK_PP(16'h346E,4);
TASK_PP(16'h346F,4);
TASK_PP(16'h3470,4);
TASK_PP(16'h3471,4);
TASK_PP(16'h3472,4);
TASK_PP(16'h3473,4);
TASK_PP(16'h3474,4);
TASK_PP(16'h3475,4);
TASK_PP(16'h3476,4);
TASK_PP(16'h3477,4);
TASK_PP(16'h3478,4);
TASK_PP(16'h3479,4);
TASK_PP(16'h347A,4);
TASK_PP(16'h347B,4);
TASK_PP(16'h347C,4);
TASK_PP(16'h347D,4);
TASK_PP(16'h347E,4);
TASK_PP(16'h347F,4);
TASK_PP(16'h3480,4);
TASK_PP(16'h3481,4);
TASK_PP(16'h3482,4);
TASK_PP(16'h3483,4);
TASK_PP(16'h3484,4);
TASK_PP(16'h3485,4);
TASK_PP(16'h3486,4);
TASK_PP(16'h3487,4);
TASK_PP(16'h3488,4);
TASK_PP(16'h3489,4);
TASK_PP(16'h348A,4);
TASK_PP(16'h348B,4);
TASK_PP(16'h348C,4);
TASK_PP(16'h348D,4);
TASK_PP(16'h348E,4);
TASK_PP(16'h348F,4);
TASK_PP(16'h3490,4);
TASK_PP(16'h3491,4);
TASK_PP(16'h3492,4);
TASK_PP(16'h3493,4);
TASK_PP(16'h3494,4);
TASK_PP(16'h3495,4);
TASK_PP(16'h3496,4);
TASK_PP(16'h3497,4);
TASK_PP(16'h3498,4);
TASK_PP(16'h3499,4);
TASK_PP(16'h349A,4);
TASK_PP(16'h349B,4);
TASK_PP(16'h349C,4);
TASK_PP(16'h349D,4);
TASK_PP(16'h349E,4);
TASK_PP(16'h349F,4);
TASK_PP(16'h34A0,4);
TASK_PP(16'h34A1,4);
TASK_PP(16'h34A2,4);
TASK_PP(16'h34A3,4);
TASK_PP(16'h34A4,4);
TASK_PP(16'h34A5,4);
TASK_PP(16'h34A6,4);
TASK_PP(16'h34A7,4);
TASK_PP(16'h34A8,4);
TASK_PP(16'h34A9,4);
TASK_PP(16'h34AA,4);
TASK_PP(16'h34AB,4);
TASK_PP(16'h34AC,4);
TASK_PP(16'h34AD,4);
TASK_PP(16'h34AE,4);
TASK_PP(16'h34AF,4);
TASK_PP(16'h34B0,4);
TASK_PP(16'h34B1,4);
TASK_PP(16'h34B2,4);
TASK_PP(16'h34B3,4);
TASK_PP(16'h34B4,4);
TASK_PP(16'h34B5,4);
TASK_PP(16'h34B6,4);
TASK_PP(16'h34B7,4);
TASK_PP(16'h34B8,4);
TASK_PP(16'h34B9,4);
TASK_PP(16'h34BA,4);
TASK_PP(16'h34BB,4);
TASK_PP(16'h34BC,4);
TASK_PP(16'h34BD,4);
TASK_PP(16'h34BE,4);
TASK_PP(16'h34BF,4);
TASK_PP(16'h34C0,4);
TASK_PP(16'h34C1,4);
TASK_PP(16'h34C2,4);
TASK_PP(16'h34C3,4);
TASK_PP(16'h34C4,4);
TASK_PP(16'h34C5,4);
TASK_PP(16'h34C6,4);
TASK_PP(16'h34C7,4);
TASK_PP(16'h34C8,4);
TASK_PP(16'h34C9,4);
TASK_PP(16'h34CA,4);
TASK_PP(16'h34CB,4);
TASK_PP(16'h34CC,4);
TASK_PP(16'h34CD,4);
TASK_PP(16'h34CE,4);
TASK_PP(16'h34CF,4);
TASK_PP(16'h34D0,4);
TASK_PP(16'h34D1,4);
TASK_PP(16'h34D2,4);
TASK_PP(16'h34D3,4);
TASK_PP(16'h34D4,4);
TASK_PP(16'h34D5,4);
TASK_PP(16'h34D6,4);
TASK_PP(16'h34D7,4);
TASK_PP(16'h34D8,4);
TASK_PP(16'h34D9,4);
TASK_PP(16'h34DA,4);
TASK_PP(16'h34DB,4);
TASK_PP(16'h34DC,4);
TASK_PP(16'h34DD,4);
TASK_PP(16'h34DE,4);
TASK_PP(16'h34DF,4);
TASK_PP(16'h34E0,4);
TASK_PP(16'h34E1,4);
TASK_PP(16'h34E2,4);
TASK_PP(16'h34E3,4);
TASK_PP(16'h34E4,4);
TASK_PP(16'h34E5,4);
TASK_PP(16'h34E6,4);
TASK_PP(16'h34E7,4);
TASK_PP(16'h34E8,4);
TASK_PP(16'h34E9,4);
TASK_PP(16'h34EA,4);
TASK_PP(16'h34EB,4);
TASK_PP(16'h34EC,4);
TASK_PP(16'h34ED,4);
TASK_PP(16'h34EE,4);
TASK_PP(16'h34EF,4);
TASK_PP(16'h34F0,4);
TASK_PP(16'h34F1,4);
TASK_PP(16'h34F2,4);
TASK_PP(16'h34F3,4);
TASK_PP(16'h34F4,4);
TASK_PP(16'h34F5,4);
TASK_PP(16'h34F6,4);
TASK_PP(16'h34F7,4);
TASK_PP(16'h34F8,4);
TASK_PP(16'h34F9,4);
TASK_PP(16'h34FA,4);
TASK_PP(16'h34FB,4);
TASK_PP(16'h34FC,4);
TASK_PP(16'h34FD,4);
TASK_PP(16'h34FE,4);
TASK_PP(16'h34FF,4);
TASK_PP(16'h3500,4);
TASK_PP(16'h3501,4);
TASK_PP(16'h3502,4);
TASK_PP(16'h3503,4);
TASK_PP(16'h3504,4);
TASK_PP(16'h3505,4);
TASK_PP(16'h3506,4);
TASK_PP(16'h3507,4);
TASK_PP(16'h3508,4);
TASK_PP(16'h3509,4);
TASK_PP(16'h350A,4);
TASK_PP(16'h350B,4);
TASK_PP(16'h350C,4);
TASK_PP(16'h350D,4);
TASK_PP(16'h350E,4);
TASK_PP(16'h350F,4);
TASK_PP(16'h3510,4);
TASK_PP(16'h3511,4);
TASK_PP(16'h3512,4);
TASK_PP(16'h3513,4);
TASK_PP(16'h3514,4);
TASK_PP(16'h3515,4);
TASK_PP(16'h3516,4);
TASK_PP(16'h3517,4);
TASK_PP(16'h3518,4);
TASK_PP(16'h3519,4);
TASK_PP(16'h351A,4);
TASK_PP(16'h351B,4);
TASK_PP(16'h351C,4);
TASK_PP(16'h351D,4);
TASK_PP(16'h351E,4);
TASK_PP(16'h351F,4);
TASK_PP(16'h3520,4);
TASK_PP(16'h3521,4);
TASK_PP(16'h3522,4);
TASK_PP(16'h3523,4);
TASK_PP(16'h3524,4);
TASK_PP(16'h3525,4);
TASK_PP(16'h3526,4);
TASK_PP(16'h3527,4);
TASK_PP(16'h3528,4);
TASK_PP(16'h3529,4);
TASK_PP(16'h352A,4);
TASK_PP(16'h352B,4);
TASK_PP(16'h352C,4);
TASK_PP(16'h352D,4);
TASK_PP(16'h352E,4);
TASK_PP(16'h352F,4);
TASK_PP(16'h3530,4);
TASK_PP(16'h3531,4);
TASK_PP(16'h3532,4);
TASK_PP(16'h3533,4);
TASK_PP(16'h3534,4);
TASK_PP(16'h3535,4);
TASK_PP(16'h3536,4);
TASK_PP(16'h3537,4);
TASK_PP(16'h3538,4);
TASK_PP(16'h3539,4);
TASK_PP(16'h353A,4);
TASK_PP(16'h353B,4);
TASK_PP(16'h353C,4);
TASK_PP(16'h353D,4);
TASK_PP(16'h353E,4);
TASK_PP(16'h353F,4);
TASK_PP(16'h3540,4);
TASK_PP(16'h3541,4);
TASK_PP(16'h3542,4);
TASK_PP(16'h3543,4);
TASK_PP(16'h3544,4);
TASK_PP(16'h3545,4);
TASK_PP(16'h3546,4);
TASK_PP(16'h3547,4);
TASK_PP(16'h3548,4);
TASK_PP(16'h3549,4);
TASK_PP(16'h354A,4);
TASK_PP(16'h354B,4);
TASK_PP(16'h354C,4);
TASK_PP(16'h354D,4);
TASK_PP(16'h354E,4);
TASK_PP(16'h354F,4);
TASK_PP(16'h3550,4);
TASK_PP(16'h3551,4);
TASK_PP(16'h3552,4);
TASK_PP(16'h3553,4);
TASK_PP(16'h3554,4);
TASK_PP(16'h3555,4);
TASK_PP(16'h3556,4);
TASK_PP(16'h3557,4);
TASK_PP(16'h3558,4);
TASK_PP(16'h3559,4);
TASK_PP(16'h355A,4);
TASK_PP(16'h355B,4);
TASK_PP(16'h355C,4);
TASK_PP(16'h355D,4);
TASK_PP(16'h355E,4);
TASK_PP(16'h355F,4);
TASK_PP(16'h3560,4);
TASK_PP(16'h3561,4);
TASK_PP(16'h3562,4);
TASK_PP(16'h3563,4);
TASK_PP(16'h3564,4);
TASK_PP(16'h3565,4);
TASK_PP(16'h3566,4);
TASK_PP(16'h3567,4);
TASK_PP(16'h3568,4);
TASK_PP(16'h3569,4);
TASK_PP(16'h356A,4);
TASK_PP(16'h356B,4);
TASK_PP(16'h356C,4);
TASK_PP(16'h356D,4);
TASK_PP(16'h356E,4);
TASK_PP(16'h356F,4);
TASK_PP(16'h3570,4);
TASK_PP(16'h3571,4);
TASK_PP(16'h3572,4);
TASK_PP(16'h3573,4);
TASK_PP(16'h3574,4);
TASK_PP(16'h3575,4);
TASK_PP(16'h3576,4);
TASK_PP(16'h3577,4);
TASK_PP(16'h3578,4);
TASK_PP(16'h3579,4);
TASK_PP(16'h357A,4);
TASK_PP(16'h357B,4);
TASK_PP(16'h357C,4);
TASK_PP(16'h357D,4);
TASK_PP(16'h357E,4);
TASK_PP(16'h357F,4);
TASK_PP(16'h3580,4);
TASK_PP(16'h3581,4);
TASK_PP(16'h3582,4);
TASK_PP(16'h3583,4);
TASK_PP(16'h3584,4);
TASK_PP(16'h3585,4);
TASK_PP(16'h3586,4);
TASK_PP(16'h3587,4);
TASK_PP(16'h3588,4);
TASK_PP(16'h3589,4);
TASK_PP(16'h358A,4);
TASK_PP(16'h358B,4);
TASK_PP(16'h358C,4);
TASK_PP(16'h358D,4);
TASK_PP(16'h358E,4);
TASK_PP(16'h358F,4);
TASK_PP(16'h3590,4);
TASK_PP(16'h3591,4);
TASK_PP(16'h3592,4);
TASK_PP(16'h3593,4);
TASK_PP(16'h3594,4);
TASK_PP(16'h3595,4);
TASK_PP(16'h3596,4);
TASK_PP(16'h3597,4);
TASK_PP(16'h3598,4);
TASK_PP(16'h3599,4);
TASK_PP(16'h359A,4);
TASK_PP(16'h359B,4);
TASK_PP(16'h359C,4);
TASK_PP(16'h359D,4);
TASK_PP(16'h359E,4);
TASK_PP(16'h359F,4);
TASK_PP(16'h35A0,4);
TASK_PP(16'h35A1,4);
TASK_PP(16'h35A2,4);
TASK_PP(16'h35A3,4);
TASK_PP(16'h35A4,4);
TASK_PP(16'h35A5,4);
TASK_PP(16'h35A6,4);
TASK_PP(16'h35A7,4);
TASK_PP(16'h35A8,4);
TASK_PP(16'h35A9,4);
TASK_PP(16'h35AA,4);
TASK_PP(16'h35AB,4);
TASK_PP(16'h35AC,4);
TASK_PP(16'h35AD,4);
TASK_PP(16'h35AE,4);
TASK_PP(16'h35AF,4);
TASK_PP(16'h35B0,4);
TASK_PP(16'h35B1,4);
TASK_PP(16'h35B2,4);
TASK_PP(16'h35B3,4);
TASK_PP(16'h35B4,4);
TASK_PP(16'h35B5,4);
TASK_PP(16'h35B6,4);
TASK_PP(16'h35B7,4);
TASK_PP(16'h35B8,4);
TASK_PP(16'h35B9,4);
TASK_PP(16'h35BA,4);
TASK_PP(16'h35BB,4);
TASK_PP(16'h35BC,4);
TASK_PP(16'h35BD,4);
TASK_PP(16'h35BE,4);
TASK_PP(16'h35BF,4);
TASK_PP(16'h35C0,4);
TASK_PP(16'h35C1,4);
TASK_PP(16'h35C2,4);
TASK_PP(16'h35C3,4);
TASK_PP(16'h35C4,4);
TASK_PP(16'h35C5,4);
TASK_PP(16'h35C6,4);
TASK_PP(16'h35C7,4);
TASK_PP(16'h35C8,4);
TASK_PP(16'h35C9,4);
TASK_PP(16'h35CA,4);
TASK_PP(16'h35CB,4);
TASK_PP(16'h35CC,4);
TASK_PP(16'h35CD,4);
TASK_PP(16'h35CE,4);
TASK_PP(16'h35CF,4);
TASK_PP(16'h35D0,4);
TASK_PP(16'h35D1,4);
TASK_PP(16'h35D2,4);
TASK_PP(16'h35D3,4);
TASK_PP(16'h35D4,4);
TASK_PP(16'h35D5,4);
TASK_PP(16'h35D6,4);
TASK_PP(16'h35D7,4);
TASK_PP(16'h35D8,4);
TASK_PP(16'h35D9,4);
TASK_PP(16'h35DA,4);
TASK_PP(16'h35DB,4);
TASK_PP(16'h35DC,4);
TASK_PP(16'h35DD,4);
TASK_PP(16'h35DE,4);
TASK_PP(16'h35DF,4);
TASK_PP(16'h35E0,4);
TASK_PP(16'h35E1,4);
TASK_PP(16'h35E2,4);
TASK_PP(16'h35E3,4);
TASK_PP(16'h35E4,4);
TASK_PP(16'h35E5,4);
TASK_PP(16'h35E6,4);
TASK_PP(16'h35E7,4);
TASK_PP(16'h35E8,4);
TASK_PP(16'h35E9,4);
TASK_PP(16'h35EA,4);
TASK_PP(16'h35EB,4);
TASK_PP(16'h35EC,4);
TASK_PP(16'h35ED,4);
TASK_PP(16'h35EE,4);
TASK_PP(16'h35EF,4);
TASK_PP(16'h35F0,4);
TASK_PP(16'h35F1,4);
TASK_PP(16'h35F2,4);
TASK_PP(16'h35F3,4);
TASK_PP(16'h35F4,4);
TASK_PP(16'h35F5,4);
TASK_PP(16'h35F6,4);
TASK_PP(16'h35F7,4);
TASK_PP(16'h35F8,4);
TASK_PP(16'h35F9,4);
TASK_PP(16'h35FA,4);
TASK_PP(16'h35FB,4);
TASK_PP(16'h35FC,4);
TASK_PP(16'h35FD,4);
TASK_PP(16'h35FE,4);
TASK_PP(16'h35FF,4);
TASK_PP(16'h3600,4);
TASK_PP(16'h3601,4);
TASK_PP(16'h3602,4);
TASK_PP(16'h3603,4);
TASK_PP(16'h3604,4);
TASK_PP(16'h3605,4);
TASK_PP(16'h3606,4);
TASK_PP(16'h3607,4);
TASK_PP(16'h3608,4);
TASK_PP(16'h3609,4);
TASK_PP(16'h360A,4);
TASK_PP(16'h360B,4);
TASK_PP(16'h360C,4);
TASK_PP(16'h360D,4);
TASK_PP(16'h360E,4);
TASK_PP(16'h360F,4);
TASK_PP(16'h3610,4);
TASK_PP(16'h3611,4);
TASK_PP(16'h3612,4);
TASK_PP(16'h3613,4);
TASK_PP(16'h3614,4);
TASK_PP(16'h3615,4);
TASK_PP(16'h3616,4);
TASK_PP(16'h3617,4);
TASK_PP(16'h3618,4);
TASK_PP(16'h3619,4);
TASK_PP(16'h361A,4);
TASK_PP(16'h361B,4);
TASK_PP(16'h361C,4);
TASK_PP(16'h361D,4);
TASK_PP(16'h361E,4);
TASK_PP(16'h361F,4);
TASK_PP(16'h3620,4);
TASK_PP(16'h3621,4);
TASK_PP(16'h3622,4);
TASK_PP(16'h3623,4);
TASK_PP(16'h3624,4);
TASK_PP(16'h3625,4);
TASK_PP(16'h3626,4);
TASK_PP(16'h3627,4);
TASK_PP(16'h3628,4);
TASK_PP(16'h3629,4);
TASK_PP(16'h362A,4);
TASK_PP(16'h362B,4);
TASK_PP(16'h362C,4);
TASK_PP(16'h362D,4);
TASK_PP(16'h362E,4);
TASK_PP(16'h362F,4);
TASK_PP(16'h3630,4);
TASK_PP(16'h3631,4);
TASK_PP(16'h3632,4);
TASK_PP(16'h3633,4);
TASK_PP(16'h3634,4);
TASK_PP(16'h3635,4);
TASK_PP(16'h3636,4);
TASK_PP(16'h3637,4);
TASK_PP(16'h3638,4);
TASK_PP(16'h3639,4);
TASK_PP(16'h363A,4);
TASK_PP(16'h363B,4);
TASK_PP(16'h363C,4);
TASK_PP(16'h363D,4);
TASK_PP(16'h363E,4);
TASK_PP(16'h363F,4);
TASK_PP(16'h3640,4);
TASK_PP(16'h3641,4);
TASK_PP(16'h3642,4);
TASK_PP(16'h3643,4);
TASK_PP(16'h3644,4);
TASK_PP(16'h3645,4);
TASK_PP(16'h3646,4);
TASK_PP(16'h3647,4);
TASK_PP(16'h3648,4);
TASK_PP(16'h3649,4);
TASK_PP(16'h364A,4);
TASK_PP(16'h364B,4);
TASK_PP(16'h364C,4);
TASK_PP(16'h364D,4);
TASK_PP(16'h364E,4);
TASK_PP(16'h364F,4);
TASK_PP(16'h3650,4);
TASK_PP(16'h3651,4);
TASK_PP(16'h3652,4);
TASK_PP(16'h3653,4);
TASK_PP(16'h3654,4);
TASK_PP(16'h3655,4);
TASK_PP(16'h3656,4);
TASK_PP(16'h3657,4);
TASK_PP(16'h3658,4);
TASK_PP(16'h3659,4);
TASK_PP(16'h365A,4);
TASK_PP(16'h365B,4);
TASK_PP(16'h365C,4);
TASK_PP(16'h365D,4);
TASK_PP(16'h365E,4);
TASK_PP(16'h365F,4);
TASK_PP(16'h3660,4);
TASK_PP(16'h3661,4);
TASK_PP(16'h3662,4);
TASK_PP(16'h3663,4);
TASK_PP(16'h3664,4);
TASK_PP(16'h3665,4);
TASK_PP(16'h3666,4);
TASK_PP(16'h3667,4);
TASK_PP(16'h3668,4);
TASK_PP(16'h3669,4);
TASK_PP(16'h366A,4);
TASK_PP(16'h366B,4);
TASK_PP(16'h366C,4);
TASK_PP(16'h366D,4);
TASK_PP(16'h366E,4);
TASK_PP(16'h366F,4);
TASK_PP(16'h3670,4);
TASK_PP(16'h3671,4);
TASK_PP(16'h3672,4);
TASK_PP(16'h3673,4);
TASK_PP(16'h3674,4);
TASK_PP(16'h3675,4);
TASK_PP(16'h3676,4);
TASK_PP(16'h3677,4);
TASK_PP(16'h3678,4);
TASK_PP(16'h3679,4);
TASK_PP(16'h367A,4);
TASK_PP(16'h367B,4);
TASK_PP(16'h367C,4);
TASK_PP(16'h367D,4);
TASK_PP(16'h367E,4);
TASK_PP(16'h367F,4);
TASK_PP(16'h3680,4);
TASK_PP(16'h3681,4);
TASK_PP(16'h3682,4);
TASK_PP(16'h3683,4);
TASK_PP(16'h3684,4);
TASK_PP(16'h3685,4);
TASK_PP(16'h3686,4);
TASK_PP(16'h3687,4);
TASK_PP(16'h3688,4);
TASK_PP(16'h3689,4);
TASK_PP(16'h368A,4);
TASK_PP(16'h368B,4);
TASK_PP(16'h368C,4);
TASK_PP(16'h368D,4);
TASK_PP(16'h368E,4);
TASK_PP(16'h368F,4);
TASK_PP(16'h3690,4);
TASK_PP(16'h3691,4);
TASK_PP(16'h3692,4);
TASK_PP(16'h3693,4);
TASK_PP(16'h3694,4);
TASK_PP(16'h3695,4);
TASK_PP(16'h3696,4);
TASK_PP(16'h3697,4);
TASK_PP(16'h3698,4);
TASK_PP(16'h3699,4);
TASK_PP(16'h369A,4);
TASK_PP(16'h369B,4);
TASK_PP(16'h369C,4);
TASK_PP(16'h369D,4);
TASK_PP(16'h369E,4);
TASK_PP(16'h369F,4);
TASK_PP(16'h36A0,4);
TASK_PP(16'h36A1,4);
TASK_PP(16'h36A2,4);
TASK_PP(16'h36A3,4);
TASK_PP(16'h36A4,4);
TASK_PP(16'h36A5,4);
TASK_PP(16'h36A6,4);
TASK_PP(16'h36A7,4);
TASK_PP(16'h36A8,4);
TASK_PP(16'h36A9,4);
TASK_PP(16'h36AA,4);
TASK_PP(16'h36AB,4);
TASK_PP(16'h36AC,4);
TASK_PP(16'h36AD,4);
TASK_PP(16'h36AE,4);
TASK_PP(16'h36AF,4);
TASK_PP(16'h36B0,4);
TASK_PP(16'h36B1,4);
TASK_PP(16'h36B2,4);
TASK_PP(16'h36B3,4);
TASK_PP(16'h36B4,4);
TASK_PP(16'h36B5,4);
TASK_PP(16'h36B6,4);
TASK_PP(16'h36B7,4);
TASK_PP(16'h36B8,4);
TASK_PP(16'h36B9,4);
TASK_PP(16'h36BA,4);
TASK_PP(16'h36BB,4);
TASK_PP(16'h36BC,4);
TASK_PP(16'h36BD,4);
TASK_PP(16'h36BE,4);
TASK_PP(16'h36BF,4);
TASK_PP(16'h36C0,4);
TASK_PP(16'h36C1,4);
TASK_PP(16'h36C2,4);
TASK_PP(16'h36C3,4);
TASK_PP(16'h36C4,4);
TASK_PP(16'h36C5,4);
TASK_PP(16'h36C6,4);
TASK_PP(16'h36C7,4);
TASK_PP(16'h36C8,4);
TASK_PP(16'h36C9,4);
TASK_PP(16'h36CA,4);
TASK_PP(16'h36CB,4);
TASK_PP(16'h36CC,4);
TASK_PP(16'h36CD,4);
TASK_PP(16'h36CE,4);
TASK_PP(16'h36CF,4);
TASK_PP(16'h36D0,4);
TASK_PP(16'h36D1,4);
TASK_PP(16'h36D2,4);
TASK_PP(16'h36D3,4);
TASK_PP(16'h36D4,4);
TASK_PP(16'h36D5,4);
TASK_PP(16'h36D6,4);
TASK_PP(16'h36D7,4);
TASK_PP(16'h36D8,4);
TASK_PP(16'h36D9,4);
TASK_PP(16'h36DA,4);
TASK_PP(16'h36DB,4);
TASK_PP(16'h36DC,4);
TASK_PP(16'h36DD,4);
TASK_PP(16'h36DE,4);
TASK_PP(16'h36DF,4);
TASK_PP(16'h36E0,4);
TASK_PP(16'h36E1,4);
TASK_PP(16'h36E2,4);
TASK_PP(16'h36E3,4);
TASK_PP(16'h36E4,4);
TASK_PP(16'h36E5,4);
TASK_PP(16'h36E6,4);
TASK_PP(16'h36E7,4);
TASK_PP(16'h36E8,4);
TASK_PP(16'h36E9,4);
TASK_PP(16'h36EA,4);
TASK_PP(16'h36EB,4);
TASK_PP(16'h36EC,4);
TASK_PP(16'h36ED,4);
TASK_PP(16'h36EE,4);
TASK_PP(16'h36EF,4);
TASK_PP(16'h36F0,4);
TASK_PP(16'h36F1,4);
TASK_PP(16'h36F2,4);
TASK_PP(16'h36F3,4);
TASK_PP(16'h36F4,4);
TASK_PP(16'h36F5,4);
TASK_PP(16'h36F6,4);
TASK_PP(16'h36F7,4);
TASK_PP(16'h36F8,4);
TASK_PP(16'h36F9,4);
TASK_PP(16'h36FA,4);
TASK_PP(16'h36FB,4);
TASK_PP(16'h36FC,4);
TASK_PP(16'h36FD,4);
TASK_PP(16'h36FE,4);
TASK_PP(16'h36FF,4);
TASK_PP(16'h3700,4);
TASK_PP(16'h3701,4);
TASK_PP(16'h3702,4);
TASK_PP(16'h3703,4);
TASK_PP(16'h3704,4);
TASK_PP(16'h3705,4);
TASK_PP(16'h3706,4);
TASK_PP(16'h3707,4);
TASK_PP(16'h3708,4);
TASK_PP(16'h3709,4);
TASK_PP(16'h370A,4);
TASK_PP(16'h370B,4);
TASK_PP(16'h370C,4);
TASK_PP(16'h370D,4);
TASK_PP(16'h370E,4);
TASK_PP(16'h370F,4);
TASK_PP(16'h3710,4);
TASK_PP(16'h3711,4);
TASK_PP(16'h3712,4);
TASK_PP(16'h3713,4);
TASK_PP(16'h3714,4);
TASK_PP(16'h3715,4);
TASK_PP(16'h3716,4);
TASK_PP(16'h3717,4);
TASK_PP(16'h3718,4);
TASK_PP(16'h3719,4);
TASK_PP(16'h371A,4);
TASK_PP(16'h371B,4);
TASK_PP(16'h371C,4);
TASK_PP(16'h371D,4);
TASK_PP(16'h371E,4);
TASK_PP(16'h371F,4);
TASK_PP(16'h3720,4);
TASK_PP(16'h3721,4);
TASK_PP(16'h3722,4);
TASK_PP(16'h3723,4);
TASK_PP(16'h3724,4);
TASK_PP(16'h3725,4);
TASK_PP(16'h3726,4);
TASK_PP(16'h3727,4);
TASK_PP(16'h3728,4);
TASK_PP(16'h3729,4);
TASK_PP(16'h372A,4);
TASK_PP(16'h372B,4);
TASK_PP(16'h372C,4);
TASK_PP(16'h372D,4);
TASK_PP(16'h372E,4);
TASK_PP(16'h372F,4);
TASK_PP(16'h3730,4);
TASK_PP(16'h3731,4);
TASK_PP(16'h3732,4);
TASK_PP(16'h3733,4);
TASK_PP(16'h3734,4);
TASK_PP(16'h3735,4);
TASK_PP(16'h3736,4);
TASK_PP(16'h3737,4);
TASK_PP(16'h3738,4);
TASK_PP(16'h3739,4);
TASK_PP(16'h373A,4);
TASK_PP(16'h373B,4);
TASK_PP(16'h373C,4);
TASK_PP(16'h373D,4);
TASK_PP(16'h373E,4);
TASK_PP(16'h373F,4);
TASK_PP(16'h3740,4);
TASK_PP(16'h3741,4);
TASK_PP(16'h3742,4);
TASK_PP(16'h3743,4);
TASK_PP(16'h3744,4);
TASK_PP(16'h3745,4);
TASK_PP(16'h3746,4);
TASK_PP(16'h3747,4);
TASK_PP(16'h3748,4);
TASK_PP(16'h3749,4);
TASK_PP(16'h374A,4);
TASK_PP(16'h374B,4);
TASK_PP(16'h374C,4);
TASK_PP(16'h374D,4);
TASK_PP(16'h374E,4);
TASK_PP(16'h374F,4);
TASK_PP(16'h3750,4);
TASK_PP(16'h3751,4);
TASK_PP(16'h3752,4);
TASK_PP(16'h3753,4);
TASK_PP(16'h3754,4);
TASK_PP(16'h3755,4);
TASK_PP(16'h3756,4);
TASK_PP(16'h3757,4);
TASK_PP(16'h3758,4);
TASK_PP(16'h3759,4);
TASK_PP(16'h375A,4);
TASK_PP(16'h375B,4);
TASK_PP(16'h375C,4);
TASK_PP(16'h375D,4);
TASK_PP(16'h375E,4);
TASK_PP(16'h375F,4);
TASK_PP(16'h3760,4);
TASK_PP(16'h3761,4);
TASK_PP(16'h3762,4);
TASK_PP(16'h3763,4);
TASK_PP(16'h3764,4);
TASK_PP(16'h3765,4);
TASK_PP(16'h3766,4);
TASK_PP(16'h3767,4);
TASK_PP(16'h3768,4);
TASK_PP(16'h3769,4);
TASK_PP(16'h376A,4);
TASK_PP(16'h376B,4);
TASK_PP(16'h376C,4);
TASK_PP(16'h376D,4);
TASK_PP(16'h376E,4);
TASK_PP(16'h376F,4);
TASK_PP(16'h3770,4);
TASK_PP(16'h3771,4);
TASK_PP(16'h3772,4);
TASK_PP(16'h3773,4);
TASK_PP(16'h3774,4);
TASK_PP(16'h3775,4);
TASK_PP(16'h3776,4);
TASK_PP(16'h3777,4);
TASK_PP(16'h3778,4);
TASK_PP(16'h3779,4);
TASK_PP(16'h377A,4);
TASK_PP(16'h377B,4);
TASK_PP(16'h377C,4);
TASK_PP(16'h377D,4);
TASK_PP(16'h377E,4);
TASK_PP(16'h377F,4);
TASK_PP(16'h3780,4);
TASK_PP(16'h3781,4);
TASK_PP(16'h3782,4);
TASK_PP(16'h3783,4);
TASK_PP(16'h3784,4);
TASK_PP(16'h3785,4);
TASK_PP(16'h3786,4);
TASK_PP(16'h3787,4);
TASK_PP(16'h3788,4);
TASK_PP(16'h3789,4);
TASK_PP(16'h378A,4);
TASK_PP(16'h378B,4);
TASK_PP(16'h378C,4);
TASK_PP(16'h378D,4);
TASK_PP(16'h378E,4);
TASK_PP(16'h378F,4);
TASK_PP(16'h3790,4);
TASK_PP(16'h3791,4);
TASK_PP(16'h3792,4);
TASK_PP(16'h3793,4);
TASK_PP(16'h3794,4);
TASK_PP(16'h3795,4);
TASK_PP(16'h3796,4);
TASK_PP(16'h3797,4);
TASK_PP(16'h3798,4);
TASK_PP(16'h3799,4);
TASK_PP(16'h379A,4);
TASK_PP(16'h379B,4);
TASK_PP(16'h379C,4);
TASK_PP(16'h379D,4);
TASK_PP(16'h379E,4);
TASK_PP(16'h379F,4);
TASK_PP(16'h37A0,4);
TASK_PP(16'h37A1,4);
TASK_PP(16'h37A2,4);
TASK_PP(16'h37A3,4);
TASK_PP(16'h37A4,4);
TASK_PP(16'h37A5,4);
TASK_PP(16'h37A6,4);
TASK_PP(16'h37A7,4);
TASK_PP(16'h37A8,4);
TASK_PP(16'h37A9,4);
TASK_PP(16'h37AA,4);
TASK_PP(16'h37AB,4);
TASK_PP(16'h37AC,4);
TASK_PP(16'h37AD,4);
TASK_PP(16'h37AE,4);
TASK_PP(16'h37AF,4);
TASK_PP(16'h37B0,4);
TASK_PP(16'h37B1,4);
TASK_PP(16'h37B2,4);
TASK_PP(16'h37B3,4);
TASK_PP(16'h37B4,4);
TASK_PP(16'h37B5,4);
TASK_PP(16'h37B6,4);
TASK_PP(16'h37B7,4);
TASK_PP(16'h37B8,4);
TASK_PP(16'h37B9,4);
TASK_PP(16'h37BA,4);
TASK_PP(16'h37BB,4);
TASK_PP(16'h37BC,4);
TASK_PP(16'h37BD,4);
TASK_PP(16'h37BE,4);
TASK_PP(16'h37BF,4);
TASK_PP(16'h37C0,4);
TASK_PP(16'h37C1,4);
TASK_PP(16'h37C2,4);
TASK_PP(16'h37C3,4);
TASK_PP(16'h37C4,4);
TASK_PP(16'h37C5,4);
TASK_PP(16'h37C6,4);
TASK_PP(16'h37C7,4);
TASK_PP(16'h37C8,4);
TASK_PP(16'h37C9,4);
TASK_PP(16'h37CA,4);
TASK_PP(16'h37CB,4);
TASK_PP(16'h37CC,4);
TASK_PP(16'h37CD,4);
TASK_PP(16'h37CE,4);
TASK_PP(16'h37CF,4);
TASK_PP(16'h37D0,4);
TASK_PP(16'h37D1,4);
TASK_PP(16'h37D2,4);
TASK_PP(16'h37D3,4);
TASK_PP(16'h37D4,4);
TASK_PP(16'h37D5,4);
TASK_PP(16'h37D6,4);
TASK_PP(16'h37D7,4);
TASK_PP(16'h37D8,4);
TASK_PP(16'h37D9,4);
TASK_PP(16'h37DA,4);
TASK_PP(16'h37DB,4);
TASK_PP(16'h37DC,4);
TASK_PP(16'h37DD,4);
TASK_PP(16'h37DE,4);
TASK_PP(16'h37DF,4);
TASK_PP(16'h37E0,4);
TASK_PP(16'h37E1,4);
TASK_PP(16'h37E2,4);
TASK_PP(16'h37E3,4);
TASK_PP(16'h37E4,4);
TASK_PP(16'h37E5,4);
TASK_PP(16'h37E6,4);
TASK_PP(16'h37E7,4);
TASK_PP(16'h37E8,4);
TASK_PP(16'h37E9,4);
TASK_PP(16'h37EA,4);
TASK_PP(16'h37EB,4);
TASK_PP(16'h37EC,4);
TASK_PP(16'h37ED,4);
TASK_PP(16'h37EE,4);
TASK_PP(16'h37EF,4);
TASK_PP(16'h37F0,4);
TASK_PP(16'h37F1,4);
TASK_PP(16'h37F2,4);
TASK_PP(16'h37F3,4);
TASK_PP(16'h37F4,4);
TASK_PP(16'h37F5,4);
TASK_PP(16'h37F6,4);
TASK_PP(16'h37F7,4);
TASK_PP(16'h37F8,4);
TASK_PP(16'h37F9,4);
TASK_PP(16'h37FA,4);
TASK_PP(16'h37FB,4);
TASK_PP(16'h37FC,4);
TASK_PP(16'h37FD,4);
TASK_PP(16'h37FE,4);
TASK_PP(16'h37FF,4);
TASK_PP(16'h3800,4);
TASK_PP(16'h3801,4);
TASK_PP(16'h3802,4);
TASK_PP(16'h3803,4);
TASK_PP(16'h3804,4);
TASK_PP(16'h3805,4);
TASK_PP(16'h3806,4);
TASK_PP(16'h3807,4);
TASK_PP(16'h3808,4);
TASK_PP(16'h3809,4);
TASK_PP(16'h380A,4);
TASK_PP(16'h380B,4);
TASK_PP(16'h380C,4);
TASK_PP(16'h380D,4);
TASK_PP(16'h380E,4);
TASK_PP(16'h380F,4);
TASK_PP(16'h3810,4);
TASK_PP(16'h3811,4);
TASK_PP(16'h3812,4);
TASK_PP(16'h3813,4);
TASK_PP(16'h3814,4);
TASK_PP(16'h3815,4);
TASK_PP(16'h3816,4);
TASK_PP(16'h3817,4);
TASK_PP(16'h3818,4);
TASK_PP(16'h3819,4);
TASK_PP(16'h381A,4);
TASK_PP(16'h381B,4);
TASK_PP(16'h381C,4);
TASK_PP(16'h381D,4);
TASK_PP(16'h381E,4);
TASK_PP(16'h381F,4);
TASK_PP(16'h3820,4);
TASK_PP(16'h3821,4);
TASK_PP(16'h3822,4);
TASK_PP(16'h3823,4);
TASK_PP(16'h3824,4);
TASK_PP(16'h3825,4);
TASK_PP(16'h3826,4);
TASK_PP(16'h3827,4);
TASK_PP(16'h3828,4);
TASK_PP(16'h3829,4);
TASK_PP(16'h382A,4);
TASK_PP(16'h382B,4);
TASK_PP(16'h382C,4);
TASK_PP(16'h382D,4);
TASK_PP(16'h382E,4);
TASK_PP(16'h382F,4);
TASK_PP(16'h3830,4);
TASK_PP(16'h3831,4);
TASK_PP(16'h3832,4);
TASK_PP(16'h3833,4);
TASK_PP(16'h3834,4);
TASK_PP(16'h3835,4);
TASK_PP(16'h3836,4);
TASK_PP(16'h3837,4);
TASK_PP(16'h3838,4);
TASK_PP(16'h3839,4);
TASK_PP(16'h383A,4);
TASK_PP(16'h383B,4);
TASK_PP(16'h383C,4);
TASK_PP(16'h383D,4);
TASK_PP(16'h383E,4);
TASK_PP(16'h383F,4);
TASK_PP(16'h3840,4);
TASK_PP(16'h3841,4);
TASK_PP(16'h3842,4);
TASK_PP(16'h3843,4);
TASK_PP(16'h3844,4);
TASK_PP(16'h3845,4);
TASK_PP(16'h3846,4);
TASK_PP(16'h3847,4);
TASK_PP(16'h3848,4);
TASK_PP(16'h3849,4);
TASK_PP(16'h384A,4);
TASK_PP(16'h384B,4);
TASK_PP(16'h384C,4);
TASK_PP(16'h384D,4);
TASK_PP(16'h384E,4);
TASK_PP(16'h384F,4);
TASK_PP(16'h3850,4);
TASK_PP(16'h3851,4);
TASK_PP(16'h3852,4);
TASK_PP(16'h3853,4);
TASK_PP(16'h3854,4);
TASK_PP(16'h3855,4);
TASK_PP(16'h3856,4);
TASK_PP(16'h3857,4);
TASK_PP(16'h3858,4);
TASK_PP(16'h3859,4);
TASK_PP(16'h385A,4);
TASK_PP(16'h385B,4);
TASK_PP(16'h385C,4);
TASK_PP(16'h385D,4);
TASK_PP(16'h385E,4);
TASK_PP(16'h385F,4);
TASK_PP(16'h3860,4);
TASK_PP(16'h3861,4);
TASK_PP(16'h3862,4);
TASK_PP(16'h3863,4);
TASK_PP(16'h3864,4);
TASK_PP(16'h3865,4);
TASK_PP(16'h3866,4);
TASK_PP(16'h3867,4);
TASK_PP(16'h3868,4);
TASK_PP(16'h3869,4);
TASK_PP(16'h386A,4);
TASK_PP(16'h386B,4);
TASK_PP(16'h386C,4);
TASK_PP(16'h386D,4);
TASK_PP(16'h386E,4);
TASK_PP(16'h386F,4);
TASK_PP(16'h3870,4);
TASK_PP(16'h3871,4);
TASK_PP(16'h3872,4);
TASK_PP(16'h3873,4);
TASK_PP(16'h3874,4);
TASK_PP(16'h3875,4);
TASK_PP(16'h3876,4);
TASK_PP(16'h3877,4);
TASK_PP(16'h3878,4);
TASK_PP(16'h3879,4);
TASK_PP(16'h387A,4);
TASK_PP(16'h387B,4);
TASK_PP(16'h387C,4);
TASK_PP(16'h387D,4);
TASK_PP(16'h387E,4);
TASK_PP(16'h387F,4);
TASK_PP(16'h3880,4);
TASK_PP(16'h3881,4);
TASK_PP(16'h3882,4);
TASK_PP(16'h3883,4);
TASK_PP(16'h3884,4);
TASK_PP(16'h3885,4);
TASK_PP(16'h3886,4);
TASK_PP(16'h3887,4);
TASK_PP(16'h3888,4);
TASK_PP(16'h3889,4);
TASK_PP(16'h388A,4);
TASK_PP(16'h388B,4);
TASK_PP(16'h388C,4);
TASK_PP(16'h388D,4);
TASK_PP(16'h388E,4);
TASK_PP(16'h388F,4);
TASK_PP(16'h3890,4);
TASK_PP(16'h3891,4);
TASK_PP(16'h3892,4);
TASK_PP(16'h3893,4);
TASK_PP(16'h3894,4);
TASK_PP(16'h3895,4);
TASK_PP(16'h3896,4);
TASK_PP(16'h3897,4);
TASK_PP(16'h3898,4);
TASK_PP(16'h3899,4);
TASK_PP(16'h389A,4);
TASK_PP(16'h389B,4);
TASK_PP(16'h389C,4);
TASK_PP(16'h389D,4);
TASK_PP(16'h389E,4);
TASK_PP(16'h389F,4);
TASK_PP(16'h38A0,4);
TASK_PP(16'h38A1,4);
TASK_PP(16'h38A2,4);
TASK_PP(16'h38A3,4);
TASK_PP(16'h38A4,4);
TASK_PP(16'h38A5,4);
TASK_PP(16'h38A6,4);
TASK_PP(16'h38A7,4);
TASK_PP(16'h38A8,4);
TASK_PP(16'h38A9,4);
TASK_PP(16'h38AA,4);
TASK_PP(16'h38AB,4);
TASK_PP(16'h38AC,4);
TASK_PP(16'h38AD,4);
TASK_PP(16'h38AE,4);
TASK_PP(16'h38AF,4);
TASK_PP(16'h38B0,4);
TASK_PP(16'h38B1,4);
TASK_PP(16'h38B2,4);
TASK_PP(16'h38B3,4);
TASK_PP(16'h38B4,4);
TASK_PP(16'h38B5,4);
TASK_PP(16'h38B6,4);
TASK_PP(16'h38B7,4);
TASK_PP(16'h38B8,4);
TASK_PP(16'h38B9,4);
TASK_PP(16'h38BA,4);
TASK_PP(16'h38BB,4);
TASK_PP(16'h38BC,4);
TASK_PP(16'h38BD,4);
TASK_PP(16'h38BE,4);
TASK_PP(16'h38BF,4);
TASK_PP(16'h38C0,4);
TASK_PP(16'h38C1,4);
TASK_PP(16'h38C2,4);
TASK_PP(16'h38C3,4);
TASK_PP(16'h38C4,4);
TASK_PP(16'h38C5,4);
TASK_PP(16'h38C6,4);
TASK_PP(16'h38C7,4);
TASK_PP(16'h38C8,4);
TASK_PP(16'h38C9,4);
TASK_PP(16'h38CA,4);
TASK_PP(16'h38CB,4);
TASK_PP(16'h38CC,4);
TASK_PP(16'h38CD,4);
TASK_PP(16'h38CE,4);
TASK_PP(16'h38CF,4);
TASK_PP(16'h38D0,4);
TASK_PP(16'h38D1,4);
TASK_PP(16'h38D2,4);
TASK_PP(16'h38D3,4);
TASK_PP(16'h38D4,4);
TASK_PP(16'h38D5,4);
TASK_PP(16'h38D6,4);
TASK_PP(16'h38D7,4);
TASK_PP(16'h38D8,4);
TASK_PP(16'h38D9,4);
TASK_PP(16'h38DA,4);
TASK_PP(16'h38DB,4);
TASK_PP(16'h38DC,4);
TASK_PP(16'h38DD,4);
TASK_PP(16'h38DE,4);
TASK_PP(16'h38DF,4);
TASK_PP(16'h38E0,4);
TASK_PP(16'h38E1,4);
TASK_PP(16'h38E2,4);
TASK_PP(16'h38E3,4);
TASK_PP(16'h38E4,4);
TASK_PP(16'h38E5,4);
TASK_PP(16'h38E6,4);
TASK_PP(16'h38E7,4);
TASK_PP(16'h38E8,4);
TASK_PP(16'h38E9,4);
TASK_PP(16'h38EA,4);
TASK_PP(16'h38EB,4);
TASK_PP(16'h38EC,4);
TASK_PP(16'h38ED,4);
TASK_PP(16'h38EE,4);
TASK_PP(16'h38EF,4);
TASK_PP(16'h38F0,4);
TASK_PP(16'h38F1,4);
TASK_PP(16'h38F2,4);
TASK_PP(16'h38F3,4);
TASK_PP(16'h38F4,4);
TASK_PP(16'h38F5,4);
TASK_PP(16'h38F6,4);
TASK_PP(16'h38F7,4);
TASK_PP(16'h38F8,4);
TASK_PP(16'h38F9,4);
TASK_PP(16'h38FA,4);
TASK_PP(16'h38FB,4);
TASK_PP(16'h38FC,4);
TASK_PP(16'h38FD,4);
TASK_PP(16'h38FE,4);
TASK_PP(16'h38FF,4);
TASK_PP(16'h3900,4);
TASK_PP(16'h3901,4);
TASK_PP(16'h3902,4);
TASK_PP(16'h3903,4);
TASK_PP(16'h3904,4);
TASK_PP(16'h3905,4);
TASK_PP(16'h3906,4);
TASK_PP(16'h3907,4);
TASK_PP(16'h3908,4);
TASK_PP(16'h3909,4);
TASK_PP(16'h390A,4);
TASK_PP(16'h390B,4);
TASK_PP(16'h390C,4);
TASK_PP(16'h390D,4);
TASK_PP(16'h390E,4);
TASK_PP(16'h390F,4);
TASK_PP(16'h3910,4);
TASK_PP(16'h3911,4);
TASK_PP(16'h3912,4);
TASK_PP(16'h3913,4);
TASK_PP(16'h3914,4);
TASK_PP(16'h3915,4);
TASK_PP(16'h3916,4);
TASK_PP(16'h3917,4);
TASK_PP(16'h3918,4);
TASK_PP(16'h3919,4);
TASK_PP(16'h391A,4);
TASK_PP(16'h391B,4);
TASK_PP(16'h391C,4);
TASK_PP(16'h391D,4);
TASK_PP(16'h391E,4);
TASK_PP(16'h391F,4);
TASK_PP(16'h3920,4);
TASK_PP(16'h3921,4);
TASK_PP(16'h3922,4);
TASK_PP(16'h3923,4);
TASK_PP(16'h3924,4);
TASK_PP(16'h3925,4);
TASK_PP(16'h3926,4);
TASK_PP(16'h3927,4);
TASK_PP(16'h3928,4);
TASK_PP(16'h3929,4);
TASK_PP(16'h392A,4);
TASK_PP(16'h392B,4);
TASK_PP(16'h392C,4);
TASK_PP(16'h392D,4);
TASK_PP(16'h392E,4);
TASK_PP(16'h392F,4);
TASK_PP(16'h3930,4);
TASK_PP(16'h3931,4);
TASK_PP(16'h3932,4);
TASK_PP(16'h3933,4);
TASK_PP(16'h3934,4);
TASK_PP(16'h3935,4);
TASK_PP(16'h3936,4);
TASK_PP(16'h3937,4);
TASK_PP(16'h3938,4);
TASK_PP(16'h3939,4);
TASK_PP(16'h393A,4);
TASK_PP(16'h393B,4);
TASK_PP(16'h393C,4);
TASK_PP(16'h393D,4);
TASK_PP(16'h393E,4);
TASK_PP(16'h393F,4);
TASK_PP(16'h3940,4);
TASK_PP(16'h3941,4);
TASK_PP(16'h3942,4);
TASK_PP(16'h3943,4);
TASK_PP(16'h3944,4);
TASK_PP(16'h3945,4);
TASK_PP(16'h3946,4);
TASK_PP(16'h3947,4);
TASK_PP(16'h3948,4);
TASK_PP(16'h3949,4);
TASK_PP(16'h394A,4);
TASK_PP(16'h394B,4);
TASK_PP(16'h394C,4);
TASK_PP(16'h394D,4);
TASK_PP(16'h394E,4);
TASK_PP(16'h394F,4);
TASK_PP(16'h3950,4);
TASK_PP(16'h3951,4);
TASK_PP(16'h3952,4);
TASK_PP(16'h3953,4);
TASK_PP(16'h3954,4);
TASK_PP(16'h3955,4);
TASK_PP(16'h3956,4);
TASK_PP(16'h3957,4);
TASK_PP(16'h3958,4);
TASK_PP(16'h3959,4);
TASK_PP(16'h395A,4);
TASK_PP(16'h395B,4);
TASK_PP(16'h395C,4);
TASK_PP(16'h395D,4);
TASK_PP(16'h395E,4);
TASK_PP(16'h395F,4);
TASK_PP(16'h3960,4);
TASK_PP(16'h3961,4);
TASK_PP(16'h3962,4);
TASK_PP(16'h3963,4);
TASK_PP(16'h3964,4);
TASK_PP(16'h3965,4);
TASK_PP(16'h3966,4);
TASK_PP(16'h3967,4);
TASK_PP(16'h3968,4);
TASK_PP(16'h3969,4);
TASK_PP(16'h396A,4);
TASK_PP(16'h396B,4);
TASK_PP(16'h396C,4);
TASK_PP(16'h396D,4);
TASK_PP(16'h396E,4);
TASK_PP(16'h396F,4);
TASK_PP(16'h3970,4);
TASK_PP(16'h3971,4);
TASK_PP(16'h3972,4);
TASK_PP(16'h3973,4);
TASK_PP(16'h3974,4);
TASK_PP(16'h3975,4);
TASK_PP(16'h3976,4);
TASK_PP(16'h3977,4);
TASK_PP(16'h3978,4);
TASK_PP(16'h3979,4);
TASK_PP(16'h397A,4);
TASK_PP(16'h397B,4);
TASK_PP(16'h397C,4);
TASK_PP(16'h397D,4);
TASK_PP(16'h397E,4);
TASK_PP(16'h397F,4);
TASK_PP(16'h3980,4);
TASK_PP(16'h3981,4);
TASK_PP(16'h3982,4);
TASK_PP(16'h3983,4);
TASK_PP(16'h3984,4);
TASK_PP(16'h3985,4);
TASK_PP(16'h3986,4);
TASK_PP(16'h3987,4);
TASK_PP(16'h3988,4);
TASK_PP(16'h3989,4);
TASK_PP(16'h398A,4);
TASK_PP(16'h398B,4);
TASK_PP(16'h398C,4);
TASK_PP(16'h398D,4);
TASK_PP(16'h398E,4);
TASK_PP(16'h398F,4);
TASK_PP(16'h3990,4);
TASK_PP(16'h3991,4);
TASK_PP(16'h3992,4);
TASK_PP(16'h3993,4);
TASK_PP(16'h3994,4);
TASK_PP(16'h3995,4);
TASK_PP(16'h3996,4);
TASK_PP(16'h3997,4);
TASK_PP(16'h3998,4);
TASK_PP(16'h3999,4);
TASK_PP(16'h399A,4);
TASK_PP(16'h399B,4);
TASK_PP(16'h399C,4);
TASK_PP(16'h399D,4);
TASK_PP(16'h399E,4);
TASK_PP(16'h399F,4);
TASK_PP(16'h39A0,4);
TASK_PP(16'h39A1,4);
TASK_PP(16'h39A2,4);
TASK_PP(16'h39A3,4);
TASK_PP(16'h39A4,4);
TASK_PP(16'h39A5,4);
TASK_PP(16'h39A6,4);
TASK_PP(16'h39A7,4);
TASK_PP(16'h39A8,4);
TASK_PP(16'h39A9,4);
TASK_PP(16'h39AA,4);
TASK_PP(16'h39AB,4);
TASK_PP(16'h39AC,4);
TASK_PP(16'h39AD,4);
TASK_PP(16'h39AE,4);
TASK_PP(16'h39AF,4);
TASK_PP(16'h39B0,4);
TASK_PP(16'h39B1,4);
TASK_PP(16'h39B2,4);
TASK_PP(16'h39B3,4);
TASK_PP(16'h39B4,4);
TASK_PP(16'h39B5,4);
TASK_PP(16'h39B6,4);
TASK_PP(16'h39B7,4);
TASK_PP(16'h39B8,4);
TASK_PP(16'h39B9,4);
TASK_PP(16'h39BA,4);
TASK_PP(16'h39BB,4);
TASK_PP(16'h39BC,4);
TASK_PP(16'h39BD,4);
TASK_PP(16'h39BE,4);
TASK_PP(16'h39BF,4);
TASK_PP(16'h39C0,4);
TASK_PP(16'h39C1,4);
TASK_PP(16'h39C2,4);
TASK_PP(16'h39C3,4);
TASK_PP(16'h39C4,4);
TASK_PP(16'h39C5,4);
TASK_PP(16'h39C6,4);
TASK_PP(16'h39C7,4);
TASK_PP(16'h39C8,4);
TASK_PP(16'h39C9,4);
TASK_PP(16'h39CA,4);
TASK_PP(16'h39CB,4);
TASK_PP(16'h39CC,4);
TASK_PP(16'h39CD,4);
TASK_PP(16'h39CE,4);
TASK_PP(16'h39CF,4);
TASK_PP(16'h39D0,4);
TASK_PP(16'h39D1,4);
TASK_PP(16'h39D2,4);
TASK_PP(16'h39D3,4);
TASK_PP(16'h39D4,4);
TASK_PP(16'h39D5,4);
TASK_PP(16'h39D6,4);
TASK_PP(16'h39D7,4);
TASK_PP(16'h39D8,4);
TASK_PP(16'h39D9,4);
TASK_PP(16'h39DA,4);
TASK_PP(16'h39DB,4);
TASK_PP(16'h39DC,4);
TASK_PP(16'h39DD,4);
TASK_PP(16'h39DE,4);
TASK_PP(16'h39DF,4);
TASK_PP(16'h39E0,4);
TASK_PP(16'h39E1,4);
TASK_PP(16'h39E2,4);
TASK_PP(16'h39E3,4);
TASK_PP(16'h39E4,4);
TASK_PP(16'h39E5,4);
TASK_PP(16'h39E6,4);
TASK_PP(16'h39E7,4);
TASK_PP(16'h39E8,4);
TASK_PP(16'h39E9,4);
TASK_PP(16'h39EA,4);
TASK_PP(16'h39EB,4);
TASK_PP(16'h39EC,4);
TASK_PP(16'h39ED,4);
TASK_PP(16'h39EE,4);
TASK_PP(16'h39EF,4);
TASK_PP(16'h39F0,4);
TASK_PP(16'h39F1,4);
TASK_PP(16'h39F2,4);
TASK_PP(16'h39F3,4);
TASK_PP(16'h39F4,4);
TASK_PP(16'h39F5,4);
TASK_PP(16'h39F6,4);
TASK_PP(16'h39F7,4);
TASK_PP(16'h39F8,4);
TASK_PP(16'h39F9,4);
TASK_PP(16'h39FA,4);
TASK_PP(16'h39FB,4);
TASK_PP(16'h39FC,4);
TASK_PP(16'h39FD,4);
TASK_PP(16'h39FE,4);
TASK_PP(16'h39FF,4);
TASK_PP(16'h3A00,4);
TASK_PP(16'h3A01,4);
TASK_PP(16'h3A02,4);
TASK_PP(16'h3A03,4);
TASK_PP(16'h3A04,4);
TASK_PP(16'h3A05,4);
TASK_PP(16'h3A06,4);
TASK_PP(16'h3A07,4);
TASK_PP(16'h3A08,4);
TASK_PP(16'h3A09,4);
TASK_PP(16'h3A0A,4);
TASK_PP(16'h3A0B,4);
TASK_PP(16'h3A0C,4);
TASK_PP(16'h3A0D,4);
TASK_PP(16'h3A0E,4);
TASK_PP(16'h3A0F,4);
TASK_PP(16'h3A10,4);
TASK_PP(16'h3A11,4);
TASK_PP(16'h3A12,4);
TASK_PP(16'h3A13,4);
TASK_PP(16'h3A14,4);
TASK_PP(16'h3A15,4);
TASK_PP(16'h3A16,4);
TASK_PP(16'h3A17,4);
TASK_PP(16'h3A18,4);
TASK_PP(16'h3A19,4);
TASK_PP(16'h3A1A,4);
TASK_PP(16'h3A1B,4);
TASK_PP(16'h3A1C,4);
TASK_PP(16'h3A1D,4);
TASK_PP(16'h3A1E,4);
TASK_PP(16'h3A1F,4);
TASK_PP(16'h3A20,4);
TASK_PP(16'h3A21,4);
TASK_PP(16'h3A22,4);
TASK_PP(16'h3A23,4);
TASK_PP(16'h3A24,4);
TASK_PP(16'h3A25,4);
TASK_PP(16'h3A26,4);
TASK_PP(16'h3A27,4);
TASK_PP(16'h3A28,4);
TASK_PP(16'h3A29,4);
TASK_PP(16'h3A2A,4);
TASK_PP(16'h3A2B,4);
TASK_PP(16'h3A2C,4);
TASK_PP(16'h3A2D,4);
TASK_PP(16'h3A2E,4);
TASK_PP(16'h3A2F,4);
TASK_PP(16'h3A30,4);
TASK_PP(16'h3A31,4);
TASK_PP(16'h3A32,4);
TASK_PP(16'h3A33,4);
TASK_PP(16'h3A34,4);
TASK_PP(16'h3A35,4);
TASK_PP(16'h3A36,4);
TASK_PP(16'h3A37,4);
TASK_PP(16'h3A38,4);
TASK_PP(16'h3A39,4);
TASK_PP(16'h3A3A,4);
TASK_PP(16'h3A3B,4);
TASK_PP(16'h3A3C,4);
TASK_PP(16'h3A3D,4);
TASK_PP(16'h3A3E,4);
TASK_PP(16'h3A3F,4);
TASK_PP(16'h3A40,4);
TASK_PP(16'h3A41,4);
TASK_PP(16'h3A42,4);
TASK_PP(16'h3A43,4);
TASK_PP(16'h3A44,4);
TASK_PP(16'h3A45,4);
TASK_PP(16'h3A46,4);
TASK_PP(16'h3A47,4);
TASK_PP(16'h3A48,4);
TASK_PP(16'h3A49,4);
TASK_PP(16'h3A4A,4);
TASK_PP(16'h3A4B,4);
TASK_PP(16'h3A4C,4);
TASK_PP(16'h3A4D,4);
TASK_PP(16'h3A4E,4);
TASK_PP(16'h3A4F,4);
TASK_PP(16'h3A50,4);
TASK_PP(16'h3A51,4);
TASK_PP(16'h3A52,4);
TASK_PP(16'h3A53,4);
TASK_PP(16'h3A54,4);
TASK_PP(16'h3A55,4);
TASK_PP(16'h3A56,4);
TASK_PP(16'h3A57,4);
TASK_PP(16'h3A58,4);
TASK_PP(16'h3A59,4);
TASK_PP(16'h3A5A,4);
TASK_PP(16'h3A5B,4);
TASK_PP(16'h3A5C,4);
TASK_PP(16'h3A5D,4);
TASK_PP(16'h3A5E,4);
TASK_PP(16'h3A5F,4);
TASK_PP(16'h3A60,4);
TASK_PP(16'h3A61,4);
TASK_PP(16'h3A62,4);
TASK_PP(16'h3A63,4);
TASK_PP(16'h3A64,4);
TASK_PP(16'h3A65,4);
TASK_PP(16'h3A66,4);
TASK_PP(16'h3A67,4);
TASK_PP(16'h3A68,4);
TASK_PP(16'h3A69,4);
TASK_PP(16'h3A6A,4);
TASK_PP(16'h3A6B,4);
TASK_PP(16'h3A6C,4);
TASK_PP(16'h3A6D,4);
TASK_PP(16'h3A6E,4);
TASK_PP(16'h3A6F,4);
TASK_PP(16'h3A70,4);
TASK_PP(16'h3A71,4);
TASK_PP(16'h3A72,4);
TASK_PP(16'h3A73,4);
TASK_PP(16'h3A74,4);
TASK_PP(16'h3A75,4);
TASK_PP(16'h3A76,4);
TASK_PP(16'h3A77,4);
TASK_PP(16'h3A78,4);
TASK_PP(16'h3A79,4);
TASK_PP(16'h3A7A,4);
TASK_PP(16'h3A7B,4);
TASK_PP(16'h3A7C,4);
TASK_PP(16'h3A7D,4);
TASK_PP(16'h3A7E,4);
TASK_PP(16'h3A7F,4);
TASK_PP(16'h3A80,4);
TASK_PP(16'h3A81,4);
TASK_PP(16'h3A82,4);
TASK_PP(16'h3A83,4);
TASK_PP(16'h3A84,4);
TASK_PP(16'h3A85,4);
TASK_PP(16'h3A86,4);
TASK_PP(16'h3A87,4);
TASK_PP(16'h3A88,4);
TASK_PP(16'h3A89,4);
TASK_PP(16'h3A8A,4);
TASK_PP(16'h3A8B,4);
TASK_PP(16'h3A8C,4);
TASK_PP(16'h3A8D,4);
TASK_PP(16'h3A8E,4);
TASK_PP(16'h3A8F,4);
TASK_PP(16'h3A90,4);
TASK_PP(16'h3A91,4);
TASK_PP(16'h3A92,4);
TASK_PP(16'h3A93,4);
TASK_PP(16'h3A94,4);
TASK_PP(16'h3A95,4);
TASK_PP(16'h3A96,4);
TASK_PP(16'h3A97,4);
TASK_PP(16'h3A98,4);
TASK_PP(16'h3A99,4);
TASK_PP(16'h3A9A,4);
TASK_PP(16'h3A9B,4);
TASK_PP(16'h3A9C,4);
TASK_PP(16'h3A9D,4);
TASK_PP(16'h3A9E,4);
TASK_PP(16'h3A9F,4);
TASK_PP(16'h3AA0,4);
TASK_PP(16'h3AA1,4);
TASK_PP(16'h3AA2,4);
TASK_PP(16'h3AA3,4);
TASK_PP(16'h3AA4,4);
TASK_PP(16'h3AA5,4);
TASK_PP(16'h3AA6,4);
TASK_PP(16'h3AA7,4);
TASK_PP(16'h3AA8,4);
TASK_PP(16'h3AA9,4);
TASK_PP(16'h3AAA,4);
TASK_PP(16'h3AAB,4);
TASK_PP(16'h3AAC,4);
TASK_PP(16'h3AAD,4);
TASK_PP(16'h3AAE,4);
TASK_PP(16'h3AAF,4);
TASK_PP(16'h3AB0,4);
TASK_PP(16'h3AB1,4);
TASK_PP(16'h3AB2,4);
TASK_PP(16'h3AB3,4);
TASK_PP(16'h3AB4,4);
TASK_PP(16'h3AB5,4);
TASK_PP(16'h3AB6,4);
TASK_PP(16'h3AB7,4);
TASK_PP(16'h3AB8,4);
TASK_PP(16'h3AB9,4);
TASK_PP(16'h3ABA,4);
TASK_PP(16'h3ABB,4);
TASK_PP(16'h3ABC,4);
TASK_PP(16'h3ABD,4);
TASK_PP(16'h3ABE,4);
TASK_PP(16'h3ABF,4);
TASK_PP(16'h3AC0,4);
TASK_PP(16'h3AC1,4);
TASK_PP(16'h3AC2,4);
TASK_PP(16'h3AC3,4);
TASK_PP(16'h3AC4,4);
TASK_PP(16'h3AC5,4);
TASK_PP(16'h3AC6,4);
TASK_PP(16'h3AC7,4);
TASK_PP(16'h3AC8,4);
TASK_PP(16'h3AC9,4);
TASK_PP(16'h3ACA,4);
TASK_PP(16'h3ACB,4);
TASK_PP(16'h3ACC,4);
TASK_PP(16'h3ACD,4);
TASK_PP(16'h3ACE,4);
TASK_PP(16'h3ACF,4);
TASK_PP(16'h3AD0,4);
TASK_PP(16'h3AD1,4);
TASK_PP(16'h3AD2,4);
TASK_PP(16'h3AD3,4);
TASK_PP(16'h3AD4,4);
TASK_PP(16'h3AD5,4);
TASK_PP(16'h3AD6,4);
TASK_PP(16'h3AD7,4);
TASK_PP(16'h3AD8,4);
TASK_PP(16'h3AD9,4);
TASK_PP(16'h3ADA,4);
TASK_PP(16'h3ADB,4);
TASK_PP(16'h3ADC,4);
TASK_PP(16'h3ADD,4);
TASK_PP(16'h3ADE,4);
TASK_PP(16'h3ADF,4);
TASK_PP(16'h3AE0,4);
TASK_PP(16'h3AE1,4);
TASK_PP(16'h3AE2,4);
TASK_PP(16'h3AE3,4);
TASK_PP(16'h3AE4,4);
TASK_PP(16'h3AE5,4);
TASK_PP(16'h3AE6,4);
TASK_PP(16'h3AE7,4);
TASK_PP(16'h3AE8,4);
TASK_PP(16'h3AE9,4);
TASK_PP(16'h3AEA,4);
TASK_PP(16'h3AEB,4);
TASK_PP(16'h3AEC,4);
TASK_PP(16'h3AED,4);
TASK_PP(16'h3AEE,4);
TASK_PP(16'h3AEF,4);
TASK_PP(16'h3AF0,4);
TASK_PP(16'h3AF1,4);
TASK_PP(16'h3AF2,4);
TASK_PP(16'h3AF3,4);
TASK_PP(16'h3AF4,4);
TASK_PP(16'h3AF5,4);
TASK_PP(16'h3AF6,4);
TASK_PP(16'h3AF7,4);
TASK_PP(16'h3AF8,4);
TASK_PP(16'h3AF9,4);
TASK_PP(16'h3AFA,4);
TASK_PP(16'h3AFB,4);
TASK_PP(16'h3AFC,4);
TASK_PP(16'h3AFD,4);
TASK_PP(16'h3AFE,4);
TASK_PP(16'h3AFF,4);
TASK_PP(16'h3B00,4);
TASK_PP(16'h3B01,4);
TASK_PP(16'h3B02,4);
TASK_PP(16'h3B03,4);
TASK_PP(16'h3B04,4);
TASK_PP(16'h3B05,4);
TASK_PP(16'h3B06,4);
TASK_PP(16'h3B07,4);
TASK_PP(16'h3B08,4);
TASK_PP(16'h3B09,4);
TASK_PP(16'h3B0A,4);
TASK_PP(16'h3B0B,4);
TASK_PP(16'h3B0C,4);
TASK_PP(16'h3B0D,4);
TASK_PP(16'h3B0E,4);
TASK_PP(16'h3B0F,4);
TASK_PP(16'h3B10,4);
TASK_PP(16'h3B11,4);
TASK_PP(16'h3B12,4);
TASK_PP(16'h3B13,4);
TASK_PP(16'h3B14,4);
TASK_PP(16'h3B15,4);
TASK_PP(16'h3B16,4);
TASK_PP(16'h3B17,4);
TASK_PP(16'h3B18,4);
TASK_PP(16'h3B19,4);
TASK_PP(16'h3B1A,4);
TASK_PP(16'h3B1B,4);
TASK_PP(16'h3B1C,4);
TASK_PP(16'h3B1D,4);
TASK_PP(16'h3B1E,4);
TASK_PP(16'h3B1F,4);
TASK_PP(16'h3B20,4);
TASK_PP(16'h3B21,4);
TASK_PP(16'h3B22,4);
TASK_PP(16'h3B23,4);
TASK_PP(16'h3B24,4);
TASK_PP(16'h3B25,4);
TASK_PP(16'h3B26,4);
TASK_PP(16'h3B27,4);
TASK_PP(16'h3B28,4);
TASK_PP(16'h3B29,4);
TASK_PP(16'h3B2A,4);
TASK_PP(16'h3B2B,4);
TASK_PP(16'h3B2C,4);
TASK_PP(16'h3B2D,4);
TASK_PP(16'h3B2E,4);
TASK_PP(16'h3B2F,4);
TASK_PP(16'h3B30,4);
TASK_PP(16'h3B31,4);
TASK_PP(16'h3B32,4);
TASK_PP(16'h3B33,4);
TASK_PP(16'h3B34,4);
TASK_PP(16'h3B35,4);
TASK_PP(16'h3B36,4);
TASK_PP(16'h3B37,4);
TASK_PP(16'h3B38,4);
TASK_PP(16'h3B39,4);
TASK_PP(16'h3B3A,4);
TASK_PP(16'h3B3B,4);
TASK_PP(16'h3B3C,4);
TASK_PP(16'h3B3D,4);
TASK_PP(16'h3B3E,4);
TASK_PP(16'h3B3F,4);
TASK_PP(16'h3B40,4);
TASK_PP(16'h3B41,4);
TASK_PP(16'h3B42,4);
TASK_PP(16'h3B43,4);
TASK_PP(16'h3B44,4);
TASK_PP(16'h3B45,4);
TASK_PP(16'h3B46,4);
TASK_PP(16'h3B47,4);
TASK_PP(16'h3B48,4);
TASK_PP(16'h3B49,4);
TASK_PP(16'h3B4A,4);
TASK_PP(16'h3B4B,4);
TASK_PP(16'h3B4C,4);
TASK_PP(16'h3B4D,4);
TASK_PP(16'h3B4E,4);
TASK_PP(16'h3B4F,4);
TASK_PP(16'h3B50,4);
TASK_PP(16'h3B51,4);
TASK_PP(16'h3B52,4);
TASK_PP(16'h3B53,4);
TASK_PP(16'h3B54,4);
TASK_PP(16'h3B55,4);
TASK_PP(16'h3B56,4);
TASK_PP(16'h3B57,4);
TASK_PP(16'h3B58,4);
TASK_PP(16'h3B59,4);
TASK_PP(16'h3B5A,4);
TASK_PP(16'h3B5B,4);
TASK_PP(16'h3B5C,4);
TASK_PP(16'h3B5D,4);
TASK_PP(16'h3B5E,4);
TASK_PP(16'h3B5F,4);
TASK_PP(16'h3B60,4);
TASK_PP(16'h3B61,4);
TASK_PP(16'h3B62,4);
TASK_PP(16'h3B63,4);
TASK_PP(16'h3B64,4);
TASK_PP(16'h3B65,4);
TASK_PP(16'h3B66,4);
TASK_PP(16'h3B67,4);
TASK_PP(16'h3B68,4);
TASK_PP(16'h3B69,4);
TASK_PP(16'h3B6A,4);
TASK_PP(16'h3B6B,4);
TASK_PP(16'h3B6C,4);
TASK_PP(16'h3B6D,4);
TASK_PP(16'h3B6E,4);
TASK_PP(16'h3B6F,4);
TASK_PP(16'h3B70,4);
TASK_PP(16'h3B71,4);
TASK_PP(16'h3B72,4);
TASK_PP(16'h3B73,4);
TASK_PP(16'h3B74,4);
TASK_PP(16'h3B75,4);
TASK_PP(16'h3B76,4);
TASK_PP(16'h3B77,4);
TASK_PP(16'h3B78,4);
TASK_PP(16'h3B79,4);
TASK_PP(16'h3B7A,4);
TASK_PP(16'h3B7B,4);
TASK_PP(16'h3B7C,4);
TASK_PP(16'h3B7D,4);
TASK_PP(16'h3B7E,4);
TASK_PP(16'h3B7F,4);
TASK_PP(16'h3B80,4);
TASK_PP(16'h3B81,4);
TASK_PP(16'h3B82,4);
TASK_PP(16'h3B83,4);
TASK_PP(16'h3B84,4);
TASK_PP(16'h3B85,4);
TASK_PP(16'h3B86,4);
TASK_PP(16'h3B87,4);
TASK_PP(16'h3B88,4);
TASK_PP(16'h3B89,4);
TASK_PP(16'h3B8A,4);
TASK_PP(16'h3B8B,4);
TASK_PP(16'h3B8C,4);
TASK_PP(16'h3B8D,4);
TASK_PP(16'h3B8E,4);
TASK_PP(16'h3B8F,4);
TASK_PP(16'h3B90,4);
TASK_PP(16'h3B91,4);
TASK_PP(16'h3B92,4);
TASK_PP(16'h3B93,4);
TASK_PP(16'h3B94,4);
TASK_PP(16'h3B95,4);
TASK_PP(16'h3B96,4);
TASK_PP(16'h3B97,4);
TASK_PP(16'h3B98,4);
TASK_PP(16'h3B99,4);
TASK_PP(16'h3B9A,4);
TASK_PP(16'h3B9B,4);
TASK_PP(16'h3B9C,4);
TASK_PP(16'h3B9D,4);
TASK_PP(16'h3B9E,4);
TASK_PP(16'h3B9F,4);
TASK_PP(16'h3BA0,4);
TASK_PP(16'h3BA1,4);
TASK_PP(16'h3BA2,4);
TASK_PP(16'h3BA3,4);
TASK_PP(16'h3BA4,4);
TASK_PP(16'h3BA5,4);
TASK_PP(16'h3BA6,4);
TASK_PP(16'h3BA7,4);
TASK_PP(16'h3BA8,4);
TASK_PP(16'h3BA9,4);
TASK_PP(16'h3BAA,4);
TASK_PP(16'h3BAB,4);
TASK_PP(16'h3BAC,4);
TASK_PP(16'h3BAD,4);
TASK_PP(16'h3BAE,4);
TASK_PP(16'h3BAF,4);
TASK_PP(16'h3BB0,4);
TASK_PP(16'h3BB1,4);
TASK_PP(16'h3BB2,4);
TASK_PP(16'h3BB3,4);
TASK_PP(16'h3BB4,4);
TASK_PP(16'h3BB5,4);
TASK_PP(16'h3BB6,4);
TASK_PP(16'h3BB7,4);
TASK_PP(16'h3BB8,4);
TASK_PP(16'h3BB9,4);
TASK_PP(16'h3BBA,4);
TASK_PP(16'h3BBB,4);
TASK_PP(16'h3BBC,4);
TASK_PP(16'h3BBD,4);
TASK_PP(16'h3BBE,4);
TASK_PP(16'h3BBF,4);
TASK_PP(16'h3BC0,4);
TASK_PP(16'h3BC1,4);
TASK_PP(16'h3BC2,4);
TASK_PP(16'h3BC3,4);
TASK_PP(16'h3BC4,4);
TASK_PP(16'h3BC5,4);
TASK_PP(16'h3BC6,4);
TASK_PP(16'h3BC7,4);
TASK_PP(16'h3BC8,4);
TASK_PP(16'h3BC9,4);
TASK_PP(16'h3BCA,4);
TASK_PP(16'h3BCB,4);
TASK_PP(16'h3BCC,4);
TASK_PP(16'h3BCD,4);
TASK_PP(16'h3BCE,4);
TASK_PP(16'h3BCF,4);
TASK_PP(16'h3BD0,4);
TASK_PP(16'h3BD1,4);
TASK_PP(16'h3BD2,4);
TASK_PP(16'h3BD3,4);
TASK_PP(16'h3BD4,4);
TASK_PP(16'h3BD5,4);
TASK_PP(16'h3BD6,4);
TASK_PP(16'h3BD7,4);
TASK_PP(16'h3BD8,4);
TASK_PP(16'h3BD9,4);
TASK_PP(16'h3BDA,4);
TASK_PP(16'h3BDB,4);
TASK_PP(16'h3BDC,4);
TASK_PP(16'h3BDD,4);
TASK_PP(16'h3BDE,4);
TASK_PP(16'h3BDF,4);
TASK_PP(16'h3BE0,4);
TASK_PP(16'h3BE1,4);
TASK_PP(16'h3BE2,4);
TASK_PP(16'h3BE3,4);
TASK_PP(16'h3BE4,4);
TASK_PP(16'h3BE5,4);
TASK_PP(16'h3BE6,4);
TASK_PP(16'h3BE7,4);
TASK_PP(16'h3BE8,4);
TASK_PP(16'h3BE9,4);
TASK_PP(16'h3BEA,4);
TASK_PP(16'h3BEB,4);
TASK_PP(16'h3BEC,4);
TASK_PP(16'h3BED,4);
TASK_PP(16'h3BEE,4);
TASK_PP(16'h3BEF,4);
TASK_PP(16'h3BF0,4);
TASK_PP(16'h3BF1,4);
TASK_PP(16'h3BF2,4);
TASK_PP(16'h3BF3,4);
TASK_PP(16'h3BF4,4);
TASK_PP(16'h3BF5,4);
TASK_PP(16'h3BF6,4);
TASK_PP(16'h3BF7,4);
TASK_PP(16'h3BF8,4);
TASK_PP(16'h3BF9,4);
TASK_PP(16'h3BFA,4);
TASK_PP(16'h3BFB,4);
TASK_PP(16'h3BFC,4);
TASK_PP(16'h3BFD,4);
TASK_PP(16'h3BFE,4);
TASK_PP(16'h3BFF,4);
TASK_PP(16'h3C00,4);
TASK_PP(16'h3C01,4);
TASK_PP(16'h3C02,4);
TASK_PP(16'h3C03,4);
TASK_PP(16'h3C04,4);
TASK_PP(16'h3C05,4);
TASK_PP(16'h3C06,4);
TASK_PP(16'h3C07,4);
TASK_PP(16'h3C08,4);
TASK_PP(16'h3C09,4);
TASK_PP(16'h3C0A,4);
TASK_PP(16'h3C0B,4);
TASK_PP(16'h3C0C,4);
TASK_PP(16'h3C0D,4);
TASK_PP(16'h3C0E,4);
TASK_PP(16'h3C0F,4);
TASK_PP(16'h3C10,4);
TASK_PP(16'h3C11,4);
TASK_PP(16'h3C12,4);
TASK_PP(16'h3C13,4);
TASK_PP(16'h3C14,4);
TASK_PP(16'h3C15,4);
TASK_PP(16'h3C16,4);
TASK_PP(16'h3C17,4);
TASK_PP(16'h3C18,4);
TASK_PP(16'h3C19,4);
TASK_PP(16'h3C1A,4);
TASK_PP(16'h3C1B,4);
TASK_PP(16'h3C1C,4);
TASK_PP(16'h3C1D,4);
TASK_PP(16'h3C1E,4);
TASK_PP(16'h3C1F,4);
TASK_PP(16'h3C20,4);
TASK_PP(16'h3C21,4);
TASK_PP(16'h3C22,4);
TASK_PP(16'h3C23,4);
TASK_PP(16'h3C24,4);
TASK_PP(16'h3C25,4);
TASK_PP(16'h3C26,4);
TASK_PP(16'h3C27,4);
TASK_PP(16'h3C28,4);
TASK_PP(16'h3C29,4);
TASK_PP(16'h3C2A,4);
TASK_PP(16'h3C2B,4);
TASK_PP(16'h3C2C,4);
TASK_PP(16'h3C2D,4);
TASK_PP(16'h3C2E,4);
TASK_PP(16'h3C2F,4);
TASK_PP(16'h3C30,4);
TASK_PP(16'h3C31,4);
TASK_PP(16'h3C32,4);
TASK_PP(16'h3C33,4);
TASK_PP(16'h3C34,4);
TASK_PP(16'h3C35,4);
TASK_PP(16'h3C36,4);
TASK_PP(16'h3C37,4);
TASK_PP(16'h3C38,4);
TASK_PP(16'h3C39,4);
TASK_PP(16'h3C3A,4);
TASK_PP(16'h3C3B,4);
TASK_PP(16'h3C3C,4);
TASK_PP(16'h3C3D,4);
TASK_PP(16'h3C3E,4);
TASK_PP(16'h3C3F,4);
TASK_PP(16'h3C40,4);
TASK_PP(16'h3C41,4);
TASK_PP(16'h3C42,4);
TASK_PP(16'h3C43,4);
TASK_PP(16'h3C44,4);
TASK_PP(16'h3C45,4);
TASK_PP(16'h3C46,4);
TASK_PP(16'h3C47,4);
TASK_PP(16'h3C48,4);
TASK_PP(16'h3C49,4);
TASK_PP(16'h3C4A,4);
TASK_PP(16'h3C4B,4);
TASK_PP(16'h3C4C,4);
TASK_PP(16'h3C4D,4);
TASK_PP(16'h3C4E,4);
TASK_PP(16'h3C4F,4);
TASK_PP(16'h3C50,4);
TASK_PP(16'h3C51,4);
TASK_PP(16'h3C52,4);
TASK_PP(16'h3C53,4);
TASK_PP(16'h3C54,4);
TASK_PP(16'h3C55,4);
TASK_PP(16'h3C56,4);
TASK_PP(16'h3C57,4);
TASK_PP(16'h3C58,4);
TASK_PP(16'h3C59,4);
TASK_PP(16'h3C5A,4);
TASK_PP(16'h3C5B,4);
TASK_PP(16'h3C5C,4);
TASK_PP(16'h3C5D,4);
TASK_PP(16'h3C5E,4);
TASK_PP(16'h3C5F,4);
TASK_PP(16'h3C60,4);
TASK_PP(16'h3C61,4);
TASK_PP(16'h3C62,4);
TASK_PP(16'h3C63,4);
TASK_PP(16'h3C64,4);
TASK_PP(16'h3C65,4);
TASK_PP(16'h3C66,4);
TASK_PP(16'h3C67,4);
TASK_PP(16'h3C68,4);
TASK_PP(16'h3C69,4);
TASK_PP(16'h3C6A,4);
TASK_PP(16'h3C6B,4);
TASK_PP(16'h3C6C,4);
TASK_PP(16'h3C6D,4);
TASK_PP(16'h3C6E,4);
TASK_PP(16'h3C6F,4);
TASK_PP(16'h3C70,4);
TASK_PP(16'h3C71,4);
TASK_PP(16'h3C72,4);
TASK_PP(16'h3C73,4);
TASK_PP(16'h3C74,4);
TASK_PP(16'h3C75,4);
TASK_PP(16'h3C76,4);
TASK_PP(16'h3C77,4);
TASK_PP(16'h3C78,4);
TASK_PP(16'h3C79,4);
TASK_PP(16'h3C7A,4);
TASK_PP(16'h3C7B,4);
TASK_PP(16'h3C7C,4);
TASK_PP(16'h3C7D,4);
TASK_PP(16'h3C7E,4);
TASK_PP(16'h3C7F,4);
TASK_PP(16'h3C80,4);
TASK_PP(16'h3C81,4);
TASK_PP(16'h3C82,4);
TASK_PP(16'h3C83,4);
TASK_PP(16'h3C84,4);
TASK_PP(16'h3C85,4);
TASK_PP(16'h3C86,4);
TASK_PP(16'h3C87,4);
TASK_PP(16'h3C88,4);
TASK_PP(16'h3C89,4);
TASK_PP(16'h3C8A,4);
TASK_PP(16'h3C8B,4);
TASK_PP(16'h3C8C,4);
TASK_PP(16'h3C8D,4);
TASK_PP(16'h3C8E,4);
TASK_PP(16'h3C8F,4);
TASK_PP(16'h3C90,4);
TASK_PP(16'h3C91,4);
TASK_PP(16'h3C92,4);
TASK_PP(16'h3C93,4);
TASK_PP(16'h3C94,4);
TASK_PP(16'h3C95,4);
TASK_PP(16'h3C96,4);
TASK_PP(16'h3C97,4);
TASK_PP(16'h3C98,4);
TASK_PP(16'h3C99,4);
TASK_PP(16'h3C9A,4);
TASK_PP(16'h3C9B,4);
TASK_PP(16'h3C9C,4);
TASK_PP(16'h3C9D,4);
TASK_PP(16'h3C9E,4);
TASK_PP(16'h3C9F,4);
TASK_PP(16'h3CA0,4);
TASK_PP(16'h3CA1,4);
TASK_PP(16'h3CA2,4);
TASK_PP(16'h3CA3,4);
TASK_PP(16'h3CA4,4);
TASK_PP(16'h3CA5,4);
TASK_PP(16'h3CA6,4);
TASK_PP(16'h3CA7,4);
TASK_PP(16'h3CA8,4);
TASK_PP(16'h3CA9,4);
TASK_PP(16'h3CAA,4);
TASK_PP(16'h3CAB,4);
TASK_PP(16'h3CAC,4);
TASK_PP(16'h3CAD,4);
TASK_PP(16'h3CAE,4);
TASK_PP(16'h3CAF,4);
TASK_PP(16'h3CB0,4);
TASK_PP(16'h3CB1,4);
TASK_PP(16'h3CB2,4);
TASK_PP(16'h3CB3,4);
TASK_PP(16'h3CB4,4);
TASK_PP(16'h3CB5,4);
TASK_PP(16'h3CB6,4);
TASK_PP(16'h3CB7,4);
TASK_PP(16'h3CB8,4);
TASK_PP(16'h3CB9,4);
TASK_PP(16'h3CBA,4);
TASK_PP(16'h3CBB,4);
TASK_PP(16'h3CBC,4);
TASK_PP(16'h3CBD,4);
TASK_PP(16'h3CBE,4);
TASK_PP(16'h3CBF,4);
TASK_PP(16'h3CC0,4);
TASK_PP(16'h3CC1,4);
TASK_PP(16'h3CC2,4);
TASK_PP(16'h3CC3,4);
TASK_PP(16'h3CC4,4);
TASK_PP(16'h3CC5,4);
TASK_PP(16'h3CC6,4);
TASK_PP(16'h3CC7,4);
TASK_PP(16'h3CC8,4);
TASK_PP(16'h3CC9,4);
TASK_PP(16'h3CCA,4);
TASK_PP(16'h3CCB,4);
TASK_PP(16'h3CCC,4);
TASK_PP(16'h3CCD,4);
TASK_PP(16'h3CCE,4);
TASK_PP(16'h3CCF,4);
TASK_PP(16'h3CD0,4);
TASK_PP(16'h3CD1,4);
TASK_PP(16'h3CD2,4);
TASK_PP(16'h3CD3,4);
TASK_PP(16'h3CD4,4);
TASK_PP(16'h3CD5,4);
TASK_PP(16'h3CD6,4);
TASK_PP(16'h3CD7,4);
TASK_PP(16'h3CD8,4);
TASK_PP(16'h3CD9,4);
TASK_PP(16'h3CDA,4);
TASK_PP(16'h3CDB,4);
TASK_PP(16'h3CDC,4);
TASK_PP(16'h3CDD,4);
TASK_PP(16'h3CDE,4);
TASK_PP(16'h3CDF,4);
TASK_PP(16'h3CE0,4);
TASK_PP(16'h3CE1,4);
TASK_PP(16'h3CE2,4);
TASK_PP(16'h3CE3,4);
TASK_PP(16'h3CE4,4);
TASK_PP(16'h3CE5,4);
TASK_PP(16'h3CE6,4);
TASK_PP(16'h3CE7,4);
TASK_PP(16'h3CE8,4);
TASK_PP(16'h3CE9,4);
TASK_PP(16'h3CEA,4);
TASK_PP(16'h3CEB,4);
TASK_PP(16'h3CEC,4);
TASK_PP(16'h3CED,4);
TASK_PP(16'h3CEE,4);
TASK_PP(16'h3CEF,4);
TASK_PP(16'h3CF0,4);
TASK_PP(16'h3CF1,4);
TASK_PP(16'h3CF2,4);
TASK_PP(16'h3CF3,4);
TASK_PP(16'h3CF4,4);
TASK_PP(16'h3CF5,4);
TASK_PP(16'h3CF6,4);
TASK_PP(16'h3CF7,4);
TASK_PP(16'h3CF8,4);
TASK_PP(16'h3CF9,4);
TASK_PP(16'h3CFA,4);
TASK_PP(16'h3CFB,4);
TASK_PP(16'h3CFC,4);
TASK_PP(16'h3CFD,4);
TASK_PP(16'h3CFE,4);
TASK_PP(16'h3CFF,4);
TASK_PP(16'h3D00,4);
TASK_PP(16'h3D01,4);
TASK_PP(16'h3D02,4);
TASK_PP(16'h3D03,4);
TASK_PP(16'h3D04,4);
TASK_PP(16'h3D05,4);
TASK_PP(16'h3D06,4);
TASK_PP(16'h3D07,4);
TASK_PP(16'h3D08,4);
TASK_PP(16'h3D09,4);
TASK_PP(16'h3D0A,4);
TASK_PP(16'h3D0B,4);
TASK_PP(16'h3D0C,4);
TASK_PP(16'h3D0D,4);
TASK_PP(16'h3D0E,4);
TASK_PP(16'h3D0F,4);
TASK_PP(16'h3D10,4);
TASK_PP(16'h3D11,4);
TASK_PP(16'h3D12,4);
TASK_PP(16'h3D13,4);
TASK_PP(16'h3D14,4);
TASK_PP(16'h3D15,4);
TASK_PP(16'h3D16,4);
TASK_PP(16'h3D17,4);
TASK_PP(16'h3D18,4);
TASK_PP(16'h3D19,4);
TASK_PP(16'h3D1A,4);
TASK_PP(16'h3D1B,4);
TASK_PP(16'h3D1C,4);
TASK_PP(16'h3D1D,4);
TASK_PP(16'h3D1E,4);
TASK_PP(16'h3D1F,4);
TASK_PP(16'h3D20,4);
TASK_PP(16'h3D21,4);
TASK_PP(16'h3D22,4);
TASK_PP(16'h3D23,4);
TASK_PP(16'h3D24,4);
TASK_PP(16'h3D25,4);
TASK_PP(16'h3D26,4);
TASK_PP(16'h3D27,4);
TASK_PP(16'h3D28,4);
TASK_PP(16'h3D29,4);
TASK_PP(16'h3D2A,4);
TASK_PP(16'h3D2B,4);
TASK_PP(16'h3D2C,4);
TASK_PP(16'h3D2D,4);
TASK_PP(16'h3D2E,4);
TASK_PP(16'h3D2F,4);
TASK_PP(16'h3D30,4);
TASK_PP(16'h3D31,4);
TASK_PP(16'h3D32,4);
TASK_PP(16'h3D33,4);
TASK_PP(16'h3D34,4);
TASK_PP(16'h3D35,4);
TASK_PP(16'h3D36,4);
TASK_PP(16'h3D37,4);
TASK_PP(16'h3D38,4);
TASK_PP(16'h3D39,4);
TASK_PP(16'h3D3A,4);
TASK_PP(16'h3D3B,4);
TASK_PP(16'h3D3C,4);
TASK_PP(16'h3D3D,4);
TASK_PP(16'h3D3E,4);
TASK_PP(16'h3D3F,4);
TASK_PP(16'h3D40,4);
TASK_PP(16'h3D41,4);
TASK_PP(16'h3D42,4);
TASK_PP(16'h3D43,4);
TASK_PP(16'h3D44,4);
TASK_PP(16'h3D45,4);
TASK_PP(16'h3D46,4);
TASK_PP(16'h3D47,4);
TASK_PP(16'h3D48,4);
TASK_PP(16'h3D49,4);
TASK_PP(16'h3D4A,4);
TASK_PP(16'h3D4B,4);
TASK_PP(16'h3D4C,4);
TASK_PP(16'h3D4D,4);
TASK_PP(16'h3D4E,4);
TASK_PP(16'h3D4F,4);
TASK_PP(16'h3D50,4);
TASK_PP(16'h3D51,4);
TASK_PP(16'h3D52,4);
TASK_PP(16'h3D53,4);
TASK_PP(16'h3D54,4);
TASK_PP(16'h3D55,4);
TASK_PP(16'h3D56,4);
TASK_PP(16'h3D57,4);
TASK_PP(16'h3D58,4);
TASK_PP(16'h3D59,4);
TASK_PP(16'h3D5A,4);
TASK_PP(16'h3D5B,4);
TASK_PP(16'h3D5C,4);
TASK_PP(16'h3D5D,4);
TASK_PP(16'h3D5E,4);
TASK_PP(16'h3D5F,4);
TASK_PP(16'h3D60,4);
TASK_PP(16'h3D61,4);
TASK_PP(16'h3D62,4);
TASK_PP(16'h3D63,4);
TASK_PP(16'h3D64,4);
TASK_PP(16'h3D65,4);
TASK_PP(16'h3D66,4);
TASK_PP(16'h3D67,4);
TASK_PP(16'h3D68,4);
TASK_PP(16'h3D69,4);
TASK_PP(16'h3D6A,4);
TASK_PP(16'h3D6B,4);
TASK_PP(16'h3D6C,4);
TASK_PP(16'h3D6D,4);
TASK_PP(16'h3D6E,4);
TASK_PP(16'h3D6F,4);
TASK_PP(16'h3D70,4);
TASK_PP(16'h3D71,4);
TASK_PP(16'h3D72,4);
TASK_PP(16'h3D73,4);
TASK_PP(16'h3D74,4);
TASK_PP(16'h3D75,4);
TASK_PP(16'h3D76,4);
TASK_PP(16'h3D77,4);
TASK_PP(16'h3D78,4);
TASK_PP(16'h3D79,4);
TASK_PP(16'h3D7A,4);
TASK_PP(16'h3D7B,4);
TASK_PP(16'h3D7C,4);
TASK_PP(16'h3D7D,4);
TASK_PP(16'h3D7E,4);
TASK_PP(16'h3D7F,4);
TASK_PP(16'h3D80,4);
TASK_PP(16'h3D81,4);
TASK_PP(16'h3D82,4);
TASK_PP(16'h3D83,4);
TASK_PP(16'h3D84,4);
TASK_PP(16'h3D85,4);
TASK_PP(16'h3D86,4);
TASK_PP(16'h3D87,4);
TASK_PP(16'h3D88,4);
TASK_PP(16'h3D89,4);
TASK_PP(16'h3D8A,4);
TASK_PP(16'h3D8B,4);
TASK_PP(16'h3D8C,4);
TASK_PP(16'h3D8D,4);
TASK_PP(16'h3D8E,4);
TASK_PP(16'h3D8F,4);
TASK_PP(16'h3D90,4);
TASK_PP(16'h3D91,4);
TASK_PP(16'h3D92,4);
TASK_PP(16'h3D93,4);
TASK_PP(16'h3D94,4);
TASK_PP(16'h3D95,4);
TASK_PP(16'h3D96,4);
TASK_PP(16'h3D97,4);
TASK_PP(16'h3D98,4);
TASK_PP(16'h3D99,4);
TASK_PP(16'h3D9A,4);
TASK_PP(16'h3D9B,4);
TASK_PP(16'h3D9C,4);
TASK_PP(16'h3D9D,4);
TASK_PP(16'h3D9E,4);
TASK_PP(16'h3D9F,4);
TASK_PP(16'h3DA0,4);
TASK_PP(16'h3DA1,4);
TASK_PP(16'h3DA2,4);
TASK_PP(16'h3DA3,4);
TASK_PP(16'h3DA4,4);
TASK_PP(16'h3DA5,4);
TASK_PP(16'h3DA6,4);
TASK_PP(16'h3DA7,4);
TASK_PP(16'h3DA8,4);
TASK_PP(16'h3DA9,4);
TASK_PP(16'h3DAA,4);
TASK_PP(16'h3DAB,4);
TASK_PP(16'h3DAC,4);
TASK_PP(16'h3DAD,4);
TASK_PP(16'h3DAE,4);
TASK_PP(16'h3DAF,4);
TASK_PP(16'h3DB0,4);
TASK_PP(16'h3DB1,4);
TASK_PP(16'h3DB2,4);
TASK_PP(16'h3DB3,4);
TASK_PP(16'h3DB4,4);
TASK_PP(16'h3DB5,4);
TASK_PP(16'h3DB6,4);
TASK_PP(16'h3DB7,4);
TASK_PP(16'h3DB8,4);
TASK_PP(16'h3DB9,4);
TASK_PP(16'h3DBA,4);
TASK_PP(16'h3DBB,4);
TASK_PP(16'h3DBC,4);
TASK_PP(16'h3DBD,4);
TASK_PP(16'h3DBE,4);
TASK_PP(16'h3DBF,4);
TASK_PP(16'h3DC0,4);
TASK_PP(16'h3DC1,4);
TASK_PP(16'h3DC2,4);
TASK_PP(16'h3DC3,4);
TASK_PP(16'h3DC4,4);
TASK_PP(16'h3DC5,4);
TASK_PP(16'h3DC6,4);
TASK_PP(16'h3DC7,4);
TASK_PP(16'h3DC8,4);
TASK_PP(16'h3DC9,4);
TASK_PP(16'h3DCA,4);
TASK_PP(16'h3DCB,4);
TASK_PP(16'h3DCC,4);
TASK_PP(16'h3DCD,4);
TASK_PP(16'h3DCE,4);
TASK_PP(16'h3DCF,4);
TASK_PP(16'h3DD0,4);
TASK_PP(16'h3DD1,4);
TASK_PP(16'h3DD2,4);
TASK_PP(16'h3DD3,4);
TASK_PP(16'h3DD4,4);
TASK_PP(16'h3DD5,4);
TASK_PP(16'h3DD6,4);
TASK_PP(16'h3DD7,4);
TASK_PP(16'h3DD8,4);
TASK_PP(16'h3DD9,4);
TASK_PP(16'h3DDA,4);
TASK_PP(16'h3DDB,4);
TASK_PP(16'h3DDC,4);
TASK_PP(16'h3DDD,4);
TASK_PP(16'h3DDE,4);
TASK_PP(16'h3DDF,4);
TASK_PP(16'h3DE0,4);
TASK_PP(16'h3DE1,4);
TASK_PP(16'h3DE2,4);
TASK_PP(16'h3DE3,4);
TASK_PP(16'h3DE4,4);
TASK_PP(16'h3DE5,4);
TASK_PP(16'h3DE6,4);
TASK_PP(16'h3DE7,4);
TASK_PP(16'h3DE8,4);
TASK_PP(16'h3DE9,4);
TASK_PP(16'h3DEA,4);
TASK_PP(16'h3DEB,4);
TASK_PP(16'h3DEC,4);
TASK_PP(16'h3DED,4);
TASK_PP(16'h3DEE,4);
TASK_PP(16'h3DEF,4);
TASK_PP(16'h3DF0,4);
TASK_PP(16'h3DF1,4);
TASK_PP(16'h3DF2,4);
TASK_PP(16'h3DF3,4);
TASK_PP(16'h3DF4,4);
TASK_PP(16'h3DF5,4);
TASK_PP(16'h3DF6,4);
TASK_PP(16'h3DF7,4);
TASK_PP(16'h3DF8,4);
TASK_PP(16'h3DF9,4);
TASK_PP(16'h3DFA,4);
TASK_PP(16'h3DFB,4);
TASK_PP(16'h3DFC,4);
TASK_PP(16'h3DFD,4);
TASK_PP(16'h3DFE,4);
TASK_PP(16'h3DFF,4);
TASK_PP(16'h3E00,4);
TASK_PP(16'h3E01,4);
TASK_PP(16'h3E02,4);
TASK_PP(16'h3E03,4);
TASK_PP(16'h3E04,4);
TASK_PP(16'h3E05,4);
TASK_PP(16'h3E06,4);
TASK_PP(16'h3E07,4);
TASK_PP(16'h3E08,4);
TASK_PP(16'h3E09,4);
TASK_PP(16'h3E0A,4);
TASK_PP(16'h3E0B,4);
TASK_PP(16'h3E0C,4);
TASK_PP(16'h3E0D,4);
TASK_PP(16'h3E0E,4);
TASK_PP(16'h3E0F,4);
TASK_PP(16'h3E10,4);
TASK_PP(16'h3E11,4);
TASK_PP(16'h3E12,4);
TASK_PP(16'h3E13,4);
TASK_PP(16'h3E14,4);
TASK_PP(16'h3E15,4);
TASK_PP(16'h3E16,4);
TASK_PP(16'h3E17,4);
TASK_PP(16'h3E18,4);
TASK_PP(16'h3E19,4);
TASK_PP(16'h3E1A,4);
TASK_PP(16'h3E1B,4);
TASK_PP(16'h3E1C,4);
TASK_PP(16'h3E1D,4);
TASK_PP(16'h3E1E,4);
TASK_PP(16'h3E1F,4);
TASK_PP(16'h3E20,4);
TASK_PP(16'h3E21,4);
TASK_PP(16'h3E22,4);
TASK_PP(16'h3E23,4);
TASK_PP(16'h3E24,4);
TASK_PP(16'h3E25,4);
TASK_PP(16'h3E26,4);
TASK_PP(16'h3E27,4);
TASK_PP(16'h3E28,4);
TASK_PP(16'h3E29,4);
TASK_PP(16'h3E2A,4);
TASK_PP(16'h3E2B,4);
TASK_PP(16'h3E2C,4);
TASK_PP(16'h3E2D,4);
TASK_PP(16'h3E2E,4);
TASK_PP(16'h3E2F,4);
TASK_PP(16'h3E30,4);
TASK_PP(16'h3E31,4);
TASK_PP(16'h3E32,4);
TASK_PP(16'h3E33,4);
TASK_PP(16'h3E34,4);
TASK_PP(16'h3E35,4);
TASK_PP(16'h3E36,4);
TASK_PP(16'h3E37,4);
TASK_PP(16'h3E38,4);
TASK_PP(16'h3E39,4);
TASK_PP(16'h3E3A,4);
TASK_PP(16'h3E3B,4);
TASK_PP(16'h3E3C,4);
TASK_PP(16'h3E3D,4);
TASK_PP(16'h3E3E,4);
TASK_PP(16'h3E3F,4);
TASK_PP(16'h3E40,4);
TASK_PP(16'h3E41,4);
TASK_PP(16'h3E42,4);
TASK_PP(16'h3E43,4);
TASK_PP(16'h3E44,4);
TASK_PP(16'h3E45,4);
TASK_PP(16'h3E46,4);
TASK_PP(16'h3E47,4);
TASK_PP(16'h3E48,4);
TASK_PP(16'h3E49,4);
TASK_PP(16'h3E4A,4);
TASK_PP(16'h3E4B,4);
TASK_PP(16'h3E4C,4);
TASK_PP(16'h3E4D,4);
TASK_PP(16'h3E4E,4);
TASK_PP(16'h3E4F,4);
TASK_PP(16'h3E50,4);
TASK_PP(16'h3E51,4);
TASK_PP(16'h3E52,4);
TASK_PP(16'h3E53,4);
TASK_PP(16'h3E54,4);
TASK_PP(16'h3E55,4);
TASK_PP(16'h3E56,4);
TASK_PP(16'h3E57,4);
TASK_PP(16'h3E58,4);
TASK_PP(16'h3E59,4);
TASK_PP(16'h3E5A,4);
TASK_PP(16'h3E5B,4);
TASK_PP(16'h3E5C,4);
TASK_PP(16'h3E5D,4);
TASK_PP(16'h3E5E,4);
TASK_PP(16'h3E5F,4);
TASK_PP(16'h3E60,4);
TASK_PP(16'h3E61,4);
TASK_PP(16'h3E62,4);
TASK_PP(16'h3E63,4);
TASK_PP(16'h3E64,4);
TASK_PP(16'h3E65,4);
TASK_PP(16'h3E66,4);
TASK_PP(16'h3E67,4);
TASK_PP(16'h3E68,4);
TASK_PP(16'h3E69,4);
TASK_PP(16'h3E6A,4);
TASK_PP(16'h3E6B,4);
TASK_PP(16'h3E6C,4);
TASK_PP(16'h3E6D,4);
TASK_PP(16'h3E6E,4);
TASK_PP(16'h3E6F,4);
TASK_PP(16'h3E70,4);
TASK_PP(16'h3E71,4);
TASK_PP(16'h3E72,4);
TASK_PP(16'h3E73,4);
TASK_PP(16'h3E74,4);
TASK_PP(16'h3E75,4);
TASK_PP(16'h3E76,4);
TASK_PP(16'h3E77,4);
TASK_PP(16'h3E78,4);
TASK_PP(16'h3E79,4);
TASK_PP(16'h3E7A,4);
TASK_PP(16'h3E7B,4);
TASK_PP(16'h3E7C,4);
TASK_PP(16'h3E7D,4);
TASK_PP(16'h3E7E,4);
TASK_PP(16'h3E7F,4);
TASK_PP(16'h3E80,4);
TASK_PP(16'h3E81,4);
TASK_PP(16'h3E82,4);
TASK_PP(16'h3E83,4);
TASK_PP(16'h3E84,4);
TASK_PP(16'h3E85,4);
TASK_PP(16'h3E86,4);
TASK_PP(16'h3E87,4);
TASK_PP(16'h3E88,4);
TASK_PP(16'h3E89,4);
TASK_PP(16'h3E8A,4);
TASK_PP(16'h3E8B,4);
TASK_PP(16'h3E8C,4);
TASK_PP(16'h3E8D,4);
TASK_PP(16'h3E8E,4);
TASK_PP(16'h3E8F,4);
TASK_PP(16'h3E90,4);
TASK_PP(16'h3E91,4);
TASK_PP(16'h3E92,4);
TASK_PP(16'h3E93,4);
TASK_PP(16'h3E94,4);
TASK_PP(16'h3E95,4);
TASK_PP(16'h3E96,4);
TASK_PP(16'h3E97,4);
TASK_PP(16'h3E98,4);
TASK_PP(16'h3E99,4);
TASK_PP(16'h3E9A,4);
TASK_PP(16'h3E9B,4);
TASK_PP(16'h3E9C,4);
TASK_PP(16'h3E9D,4);
TASK_PP(16'h3E9E,4);
TASK_PP(16'h3E9F,4);
TASK_PP(16'h3EA0,4);
TASK_PP(16'h3EA1,4);
TASK_PP(16'h3EA2,4);
TASK_PP(16'h3EA3,4);
TASK_PP(16'h3EA4,4);
TASK_PP(16'h3EA5,4);
TASK_PP(16'h3EA6,4);
TASK_PP(16'h3EA7,4);
TASK_PP(16'h3EA8,4);
TASK_PP(16'h3EA9,4);
TASK_PP(16'h3EAA,4);
TASK_PP(16'h3EAB,4);
TASK_PP(16'h3EAC,4);
TASK_PP(16'h3EAD,4);
TASK_PP(16'h3EAE,4);
TASK_PP(16'h3EAF,4);
TASK_PP(16'h3EB0,4);
TASK_PP(16'h3EB1,4);
TASK_PP(16'h3EB2,4);
TASK_PP(16'h3EB3,4);
TASK_PP(16'h3EB4,4);
TASK_PP(16'h3EB5,4);
TASK_PP(16'h3EB6,4);
TASK_PP(16'h3EB7,4);
TASK_PP(16'h3EB8,4);
TASK_PP(16'h3EB9,4);
TASK_PP(16'h3EBA,4);
TASK_PP(16'h3EBB,4);
TASK_PP(16'h3EBC,4);
TASK_PP(16'h3EBD,4);
TASK_PP(16'h3EBE,4);
TASK_PP(16'h3EBF,4);
TASK_PP(16'h3EC0,4);
TASK_PP(16'h3EC1,4);
TASK_PP(16'h3EC2,4);
TASK_PP(16'h3EC3,4);
TASK_PP(16'h3EC4,4);
TASK_PP(16'h3EC5,4);
TASK_PP(16'h3EC6,4);
TASK_PP(16'h3EC7,4);
TASK_PP(16'h3EC8,4);
TASK_PP(16'h3EC9,4);
TASK_PP(16'h3ECA,4);
TASK_PP(16'h3ECB,4);
TASK_PP(16'h3ECC,4);
TASK_PP(16'h3ECD,4);
TASK_PP(16'h3ECE,4);
TASK_PP(16'h3ECF,4);
TASK_PP(16'h3ED0,4);
TASK_PP(16'h3ED1,4);
TASK_PP(16'h3ED2,4);
TASK_PP(16'h3ED3,4);
TASK_PP(16'h3ED4,4);
TASK_PP(16'h3ED5,4);
TASK_PP(16'h3ED6,4);
TASK_PP(16'h3ED7,4);
TASK_PP(16'h3ED8,4);
TASK_PP(16'h3ED9,4);
TASK_PP(16'h3EDA,4);
TASK_PP(16'h3EDB,4);
TASK_PP(16'h3EDC,4);
TASK_PP(16'h3EDD,4);
TASK_PP(16'h3EDE,4);
TASK_PP(16'h3EDF,4);
TASK_PP(16'h3EE0,4);
TASK_PP(16'h3EE1,4);
TASK_PP(16'h3EE2,4);
TASK_PP(16'h3EE3,4);
TASK_PP(16'h3EE4,4);
TASK_PP(16'h3EE5,4);
TASK_PP(16'h3EE6,4);
TASK_PP(16'h3EE7,4);
TASK_PP(16'h3EE8,4);
TASK_PP(16'h3EE9,4);
TASK_PP(16'h3EEA,4);
TASK_PP(16'h3EEB,4);
TASK_PP(16'h3EEC,4);
TASK_PP(16'h3EED,4);
TASK_PP(16'h3EEE,4);
TASK_PP(16'h3EEF,4);
TASK_PP(16'h3EF0,4);
TASK_PP(16'h3EF1,4);
TASK_PP(16'h3EF2,4);
TASK_PP(16'h3EF3,4);
TASK_PP(16'h3EF4,4);
TASK_PP(16'h3EF5,4);
TASK_PP(16'h3EF6,4);
TASK_PP(16'h3EF7,4);
TASK_PP(16'h3EF8,4);
TASK_PP(16'h3EF9,4);
TASK_PP(16'h3EFA,4);
TASK_PP(16'h3EFB,4);
TASK_PP(16'h3EFC,4);
TASK_PP(16'h3EFD,4);
TASK_PP(16'h3EFE,4);
TASK_PP(16'h3EFF,4);
TASK_PP(16'h3F00,4);
TASK_PP(16'h3F01,4);
TASK_PP(16'h3F02,4);
TASK_PP(16'h3F03,4);
TASK_PP(16'h3F04,4);
TASK_PP(16'h3F05,4);
TASK_PP(16'h3F06,4);
TASK_PP(16'h3F07,4);
TASK_PP(16'h3F08,4);
TASK_PP(16'h3F09,4);
TASK_PP(16'h3F0A,4);
TASK_PP(16'h3F0B,4);
TASK_PP(16'h3F0C,4);
TASK_PP(16'h3F0D,4);
TASK_PP(16'h3F0E,4);
TASK_PP(16'h3F0F,4);
TASK_PP(16'h3F10,4);
TASK_PP(16'h3F11,4);
TASK_PP(16'h3F12,4);
TASK_PP(16'h3F13,4);
TASK_PP(16'h3F14,4);
TASK_PP(16'h3F15,4);
TASK_PP(16'h3F16,4);
TASK_PP(16'h3F17,4);
TASK_PP(16'h3F18,4);
TASK_PP(16'h3F19,4);
TASK_PP(16'h3F1A,4);
TASK_PP(16'h3F1B,4);
TASK_PP(16'h3F1C,4);
TASK_PP(16'h3F1D,4);
TASK_PP(16'h3F1E,4);
TASK_PP(16'h3F1F,4);
TASK_PP(16'h3F20,4);
TASK_PP(16'h3F21,4);
TASK_PP(16'h3F22,4);
TASK_PP(16'h3F23,4);
TASK_PP(16'h3F24,4);
TASK_PP(16'h3F25,4);
TASK_PP(16'h3F26,4);
TASK_PP(16'h3F27,4);
TASK_PP(16'h3F28,4);
TASK_PP(16'h3F29,4);
TASK_PP(16'h3F2A,4);
TASK_PP(16'h3F2B,4);
TASK_PP(16'h3F2C,4);
TASK_PP(16'h3F2D,4);
TASK_PP(16'h3F2E,4);
TASK_PP(16'h3F2F,4);
TASK_PP(16'h3F30,4);
TASK_PP(16'h3F31,4);
TASK_PP(16'h3F32,4);
TASK_PP(16'h3F33,4);
TASK_PP(16'h3F34,4);
TASK_PP(16'h3F35,4);
TASK_PP(16'h3F36,4);
TASK_PP(16'h3F37,4);
TASK_PP(16'h3F38,4);
TASK_PP(16'h3F39,4);
TASK_PP(16'h3F3A,4);
TASK_PP(16'h3F3B,4);
TASK_PP(16'h3F3C,4);
TASK_PP(16'h3F3D,4);
TASK_PP(16'h3F3E,4);
TASK_PP(16'h3F3F,4);
TASK_PP(16'h3F40,4);
TASK_PP(16'h3F41,4);
TASK_PP(16'h3F42,4);
TASK_PP(16'h3F43,4);
TASK_PP(16'h3F44,4);
TASK_PP(16'h3F45,4);
TASK_PP(16'h3F46,4);
TASK_PP(16'h3F47,4);
TASK_PP(16'h3F48,4);
TASK_PP(16'h3F49,4);
TASK_PP(16'h3F4A,4);
TASK_PP(16'h3F4B,4);
TASK_PP(16'h3F4C,4);
TASK_PP(16'h3F4D,4);
TASK_PP(16'h3F4E,4);
TASK_PP(16'h3F4F,4);
TASK_PP(16'h3F50,4);
TASK_PP(16'h3F51,4);
TASK_PP(16'h3F52,4);
TASK_PP(16'h3F53,4);
TASK_PP(16'h3F54,4);
TASK_PP(16'h3F55,4);
TASK_PP(16'h3F56,4);
TASK_PP(16'h3F57,4);
TASK_PP(16'h3F58,4);
TASK_PP(16'h3F59,4);
TASK_PP(16'h3F5A,4);
TASK_PP(16'h3F5B,4);
TASK_PP(16'h3F5C,4);
TASK_PP(16'h3F5D,4);
TASK_PP(16'h3F5E,4);
TASK_PP(16'h3F5F,4);
TASK_PP(16'h3F60,4);
TASK_PP(16'h3F61,4);
TASK_PP(16'h3F62,4);
TASK_PP(16'h3F63,4);
TASK_PP(16'h3F64,4);
TASK_PP(16'h3F65,4);
TASK_PP(16'h3F66,4);
TASK_PP(16'h3F67,4);
TASK_PP(16'h3F68,4);
TASK_PP(16'h3F69,4);
TASK_PP(16'h3F6A,4);
TASK_PP(16'h3F6B,4);
TASK_PP(16'h3F6C,4);
TASK_PP(16'h3F6D,4);
TASK_PP(16'h3F6E,4);
TASK_PP(16'h3F6F,4);
TASK_PP(16'h3F70,4);
TASK_PP(16'h3F71,4);
TASK_PP(16'h3F72,4);
TASK_PP(16'h3F73,4);
TASK_PP(16'h3F74,4);
TASK_PP(16'h3F75,4);
TASK_PP(16'h3F76,4);
TASK_PP(16'h3F77,4);
TASK_PP(16'h3F78,4);
TASK_PP(16'h3F79,4);
TASK_PP(16'h3F7A,4);
TASK_PP(16'h3F7B,4);
TASK_PP(16'h3F7C,4);
TASK_PP(16'h3F7D,4);
TASK_PP(16'h3F7E,4);
TASK_PP(16'h3F7F,4);
TASK_PP(16'h3F80,4);
TASK_PP(16'h3F81,4);
TASK_PP(16'h3F82,4);
TASK_PP(16'h3F83,4);
TASK_PP(16'h3F84,4);
TASK_PP(16'h3F85,4);
TASK_PP(16'h3F86,4);
TASK_PP(16'h3F87,4);
TASK_PP(16'h3F88,4);
TASK_PP(16'h3F89,4);
TASK_PP(16'h3F8A,4);
TASK_PP(16'h3F8B,4);
TASK_PP(16'h3F8C,4);
TASK_PP(16'h3F8D,4);
TASK_PP(16'h3F8E,4);
TASK_PP(16'h3F8F,4);
TASK_PP(16'h3F90,4);
TASK_PP(16'h3F91,4);
TASK_PP(16'h3F92,4);
TASK_PP(16'h3F93,4);
TASK_PP(16'h3F94,4);
TASK_PP(16'h3F95,4);
TASK_PP(16'h3F96,4);
TASK_PP(16'h3F97,4);
TASK_PP(16'h3F98,4);
TASK_PP(16'h3F99,4);
TASK_PP(16'h3F9A,4);
TASK_PP(16'h3F9B,4);
TASK_PP(16'h3F9C,4);
TASK_PP(16'h3F9D,4);
TASK_PP(16'h3F9E,4);
TASK_PP(16'h3F9F,4);
TASK_PP(16'h3FA0,4);
TASK_PP(16'h3FA1,4);
TASK_PP(16'h3FA2,4);
TASK_PP(16'h3FA3,4);
TASK_PP(16'h3FA4,4);
TASK_PP(16'h3FA5,4);
TASK_PP(16'h3FA6,4);
TASK_PP(16'h3FA7,4);
TASK_PP(16'h3FA8,4);
TASK_PP(16'h3FA9,4);
TASK_PP(16'h3FAA,4);
TASK_PP(16'h3FAB,4);
TASK_PP(16'h3FAC,4);
TASK_PP(16'h3FAD,4);
TASK_PP(16'h3FAE,4);
TASK_PP(16'h3FAF,4);
TASK_PP(16'h3FB0,4);
TASK_PP(16'h3FB1,4);
TASK_PP(16'h3FB2,4);
TASK_PP(16'h3FB3,4);
TASK_PP(16'h3FB4,4);
TASK_PP(16'h3FB5,4);
TASK_PP(16'h3FB6,4);
TASK_PP(16'h3FB7,4);
TASK_PP(16'h3FB8,4);
TASK_PP(16'h3FB9,4);
TASK_PP(16'h3FBA,4);
TASK_PP(16'h3FBB,4);
TASK_PP(16'h3FBC,4);
TASK_PP(16'h3FBD,4);
TASK_PP(16'h3FBE,4);
TASK_PP(16'h3FBF,4);
TASK_PP(16'h3FC0,4);
TASK_PP(16'h3FC1,4);
TASK_PP(16'h3FC2,4);
TASK_PP(16'h3FC3,4);
TASK_PP(16'h3FC4,4);
TASK_PP(16'h3FC5,4);
TASK_PP(16'h3FC6,4);
TASK_PP(16'h3FC7,4);
TASK_PP(16'h3FC8,4);
TASK_PP(16'h3FC9,4);
TASK_PP(16'h3FCA,4);
TASK_PP(16'h3FCB,4);
TASK_PP(16'h3FCC,4);
TASK_PP(16'h3FCD,4);
TASK_PP(16'h3FCE,4);
TASK_PP(16'h3FCF,4);
TASK_PP(16'h3FD0,4);
TASK_PP(16'h3FD1,4);
TASK_PP(16'h3FD2,4);
TASK_PP(16'h3FD3,4);
TASK_PP(16'h3FD4,4);
TASK_PP(16'h3FD5,4);
TASK_PP(16'h3FD6,4);
TASK_PP(16'h3FD7,4);
TASK_PP(16'h3FD8,4);
TASK_PP(16'h3FD9,4);
TASK_PP(16'h3FDA,4);
TASK_PP(16'h3FDB,4);
TASK_PP(16'h3FDC,4);
TASK_PP(16'h3FDD,4);
TASK_PP(16'h3FDE,4);
TASK_PP(16'h3FDF,4);
TASK_PP(16'h3FE0,4);
TASK_PP(16'h3FE1,4);
TASK_PP(16'h3FE2,4);
TASK_PP(16'h3FE3,4);
TASK_PP(16'h3FE4,4);
TASK_PP(16'h3FE5,4);
TASK_PP(16'h3FE6,4);
TASK_PP(16'h3FE7,4);
TASK_PP(16'h3FE8,4);
TASK_PP(16'h3FE9,4);
TASK_PP(16'h3FEA,4);
TASK_PP(16'h3FEB,4);
TASK_PP(16'h3FEC,4);
TASK_PP(16'h3FED,4);
TASK_PP(16'h3FEE,4);
TASK_PP(16'h3FEF,4);
TASK_PP(16'h3FF0,4);
TASK_PP(16'h3FF1,4);
TASK_PP(16'h3FF2,4);
TASK_PP(16'h3FF3,4);
TASK_PP(16'h3FF4,4);
TASK_PP(16'h3FF5,4);
TASK_PP(16'h3FF6,4);
TASK_PP(16'h3FF7,4);
TASK_PP(16'h3FF8,4);
TASK_PP(16'h3FF9,4);
TASK_PP(16'h3FFA,4);
TASK_PP(16'h3FFB,4);
TASK_PP(16'h3FFC,4);
TASK_PP(16'h3FFD,4);
TASK_PP(16'h3FFE,4);
TASK_PP(16'h3FFF,4);
TASK_PP(16'h4000,4);
TASK_PP(16'h4001,4);
TASK_PP(16'h4002,4);
TASK_PP(16'h4003,4);
TASK_PP(16'h4004,4);
TASK_PP(16'h4005,4);
TASK_PP(16'h4006,4);
TASK_PP(16'h4007,4);
TASK_PP(16'h4008,4);
TASK_PP(16'h4009,4);
TASK_PP(16'h400A,4);
TASK_PP(16'h400B,4);
TASK_PP(16'h400C,4);
TASK_PP(16'h400D,4);
TASK_PP(16'h400E,4);
TASK_PP(16'h400F,4);
TASK_PP(16'h4010,4);
TASK_PP(16'h4011,4);
TASK_PP(16'h4012,4);
TASK_PP(16'h4013,4);
TASK_PP(16'h4014,4);
TASK_PP(16'h4015,4);
TASK_PP(16'h4016,4);
TASK_PP(16'h4017,4);
TASK_PP(16'h4018,4);
TASK_PP(16'h4019,4);
TASK_PP(16'h401A,4);
TASK_PP(16'h401B,4);
TASK_PP(16'h401C,4);
TASK_PP(16'h401D,4);
TASK_PP(16'h401E,4);
TASK_PP(16'h401F,4);
TASK_PP(16'h4020,4);
TASK_PP(16'h4021,4);
TASK_PP(16'h4022,4);
TASK_PP(16'h4023,4);
TASK_PP(16'h4024,4);
TASK_PP(16'h4025,4);
TASK_PP(16'h4026,4);
TASK_PP(16'h4027,4);
TASK_PP(16'h4028,4);
TASK_PP(16'h4029,4);
TASK_PP(16'h402A,4);
TASK_PP(16'h402B,4);
TASK_PP(16'h402C,4);
TASK_PP(16'h402D,4);
TASK_PP(16'h402E,4);
TASK_PP(16'h402F,4);
TASK_PP(16'h4030,4);
TASK_PP(16'h4031,4);
TASK_PP(16'h4032,4);
TASK_PP(16'h4033,4);
TASK_PP(16'h4034,4);
TASK_PP(16'h4035,4);
TASK_PP(16'h4036,4);
TASK_PP(16'h4037,4);
TASK_PP(16'h4038,4);
TASK_PP(16'h4039,4);
TASK_PP(16'h403A,4);
TASK_PP(16'h403B,4);
TASK_PP(16'h403C,4);
TASK_PP(16'h403D,4);
TASK_PP(16'h403E,4);
TASK_PP(16'h403F,4);
TASK_PP(16'h4040,4);
TASK_PP(16'h4041,4);
TASK_PP(16'h4042,4);
TASK_PP(16'h4043,4);
TASK_PP(16'h4044,4);
TASK_PP(16'h4045,4);
TASK_PP(16'h4046,4);
TASK_PP(16'h4047,4);
TASK_PP(16'h4048,4);
TASK_PP(16'h4049,4);
TASK_PP(16'h404A,4);
TASK_PP(16'h404B,4);
TASK_PP(16'h404C,4);
TASK_PP(16'h404D,4);
TASK_PP(16'h404E,4);
TASK_PP(16'h404F,4);
TASK_PP(16'h4050,4);
TASK_PP(16'h4051,4);
TASK_PP(16'h4052,4);
TASK_PP(16'h4053,4);
TASK_PP(16'h4054,4);
TASK_PP(16'h4055,4);
TASK_PP(16'h4056,4);
TASK_PP(16'h4057,4);
TASK_PP(16'h4058,4);
TASK_PP(16'h4059,4);
TASK_PP(16'h405A,4);
TASK_PP(16'h405B,4);
TASK_PP(16'h405C,4);
TASK_PP(16'h405D,4);
TASK_PP(16'h405E,4);
TASK_PP(16'h405F,4);
TASK_PP(16'h4060,4);
TASK_PP(16'h4061,4);
TASK_PP(16'h4062,4);
TASK_PP(16'h4063,4);
TASK_PP(16'h4064,4);
TASK_PP(16'h4065,4);
TASK_PP(16'h4066,4);
TASK_PP(16'h4067,4);
TASK_PP(16'h4068,4);
TASK_PP(16'h4069,4);
TASK_PP(16'h406A,4);
TASK_PP(16'h406B,4);
TASK_PP(16'h406C,4);
TASK_PP(16'h406D,4);
TASK_PP(16'h406E,4);
TASK_PP(16'h406F,4);
TASK_PP(16'h4070,4);
TASK_PP(16'h4071,4);
TASK_PP(16'h4072,4);
TASK_PP(16'h4073,4);
TASK_PP(16'h4074,4);
TASK_PP(16'h4075,4);
TASK_PP(16'h4076,4);
TASK_PP(16'h4077,4);
TASK_PP(16'h4078,4);
TASK_PP(16'h4079,4);
TASK_PP(16'h407A,4);
TASK_PP(16'h407B,4);
TASK_PP(16'h407C,4);
TASK_PP(16'h407D,4);
TASK_PP(16'h407E,4);
TASK_PP(16'h407F,4);
TASK_PP(16'h4080,4);
TASK_PP(16'h4081,4);
TASK_PP(16'h4082,4);
TASK_PP(16'h4083,4);
TASK_PP(16'h4084,4);
TASK_PP(16'h4085,4);
TASK_PP(16'h4086,4);
TASK_PP(16'h4087,4);
TASK_PP(16'h4088,4);
TASK_PP(16'h4089,4);
TASK_PP(16'h408A,4);
TASK_PP(16'h408B,4);
TASK_PP(16'h408C,4);
TASK_PP(16'h408D,4);
TASK_PP(16'h408E,4);
TASK_PP(16'h408F,4);
TASK_PP(16'h4090,4);
TASK_PP(16'h4091,4);
TASK_PP(16'h4092,4);
TASK_PP(16'h4093,4);
TASK_PP(16'h4094,4);
TASK_PP(16'h4095,4);
TASK_PP(16'h4096,4);
TASK_PP(16'h4097,4);
TASK_PP(16'h4098,4);
TASK_PP(16'h4099,4);
TASK_PP(16'h409A,4);
TASK_PP(16'h409B,4);
TASK_PP(16'h409C,4);
TASK_PP(16'h409D,4);
TASK_PP(16'h409E,4);
TASK_PP(16'h409F,4);
TASK_PP(16'h40A0,4);
TASK_PP(16'h40A1,4);
TASK_PP(16'h40A2,4);
TASK_PP(16'h40A3,4);
TASK_PP(16'h40A4,4);
TASK_PP(16'h40A5,4);
TASK_PP(16'h40A6,4);
TASK_PP(16'h40A7,4);
TASK_PP(16'h40A8,4);
TASK_PP(16'h40A9,4);
TASK_PP(16'h40AA,4);
TASK_PP(16'h40AB,4);
TASK_PP(16'h40AC,4);
TASK_PP(16'h40AD,4);
TASK_PP(16'h40AE,4);
TASK_PP(16'h40AF,4);
TASK_PP(16'h40B0,4);
TASK_PP(16'h40B1,4);
TASK_PP(16'h40B2,4);
TASK_PP(16'h40B3,4);
TASK_PP(16'h40B4,4);
TASK_PP(16'h40B5,4);
TASK_PP(16'h40B6,4);
TASK_PP(16'h40B7,4);
TASK_PP(16'h40B8,4);
TASK_PP(16'h40B9,4);
TASK_PP(16'h40BA,4);
TASK_PP(16'h40BB,4);
TASK_PP(16'h40BC,4);
TASK_PP(16'h40BD,4);
TASK_PP(16'h40BE,4);
TASK_PP(16'h40BF,4);
TASK_PP(16'h40C0,4);
TASK_PP(16'h40C1,4);
TASK_PP(16'h40C2,4);
TASK_PP(16'h40C3,4);
TASK_PP(16'h40C4,4);
TASK_PP(16'h40C5,4);
TASK_PP(16'h40C6,4);
TASK_PP(16'h40C7,4);
TASK_PP(16'h40C8,4);
TASK_PP(16'h40C9,4);
TASK_PP(16'h40CA,4);
TASK_PP(16'h40CB,4);
TASK_PP(16'h40CC,4);
TASK_PP(16'h40CD,4);
TASK_PP(16'h40CE,4);
TASK_PP(16'h40CF,4);
TASK_PP(16'h40D0,4);
TASK_PP(16'h40D1,4);
TASK_PP(16'h40D2,4);
TASK_PP(16'h40D3,4);
TASK_PP(16'h40D4,4);
TASK_PP(16'h40D5,4);
TASK_PP(16'h40D6,4);
TASK_PP(16'h40D7,4);
TASK_PP(16'h40D8,4);
TASK_PP(16'h40D9,4);
TASK_PP(16'h40DA,4);
TASK_PP(16'h40DB,4);
TASK_PP(16'h40DC,4);
TASK_PP(16'h40DD,4);
TASK_PP(16'h40DE,4);
TASK_PP(16'h40DF,4);
TASK_PP(16'h40E0,4);
TASK_PP(16'h40E1,4);
TASK_PP(16'h40E2,4);
TASK_PP(16'h40E3,4);
TASK_PP(16'h40E4,4);
TASK_PP(16'h40E5,4);
TASK_PP(16'h40E6,4);
TASK_PP(16'h40E7,4);
TASK_PP(16'h40E8,4);
TASK_PP(16'h40E9,4);
TASK_PP(16'h40EA,4);
TASK_PP(16'h40EB,4);
TASK_PP(16'h40EC,4);
TASK_PP(16'h40ED,4);
TASK_PP(16'h40EE,4);
TASK_PP(16'h40EF,4);
TASK_PP(16'h40F0,4);
TASK_PP(16'h40F1,4);
TASK_PP(16'h40F2,4);
TASK_PP(16'h40F3,4);
TASK_PP(16'h40F4,4);
TASK_PP(16'h40F5,4);
TASK_PP(16'h40F6,4);
TASK_PP(16'h40F7,4);
TASK_PP(16'h40F8,4);
TASK_PP(16'h40F9,4);
TASK_PP(16'h40FA,4);
TASK_PP(16'h40FB,4);
TASK_PP(16'h40FC,4);
TASK_PP(16'h40FD,4);
TASK_PP(16'h40FE,4);
TASK_PP(16'h40FF,4);
TASK_PP(16'h4100,4);
TASK_PP(16'h4101,4);
TASK_PP(16'h4102,4);
TASK_PP(16'h4103,4);
TASK_PP(16'h4104,4);
TASK_PP(16'h4105,4);
TASK_PP(16'h4106,4);
TASK_PP(16'h4107,4);
TASK_PP(16'h4108,4);
TASK_PP(16'h4109,4);
TASK_PP(16'h410A,4);
TASK_PP(16'h410B,4);
TASK_PP(16'h410C,4);
TASK_PP(16'h410D,4);
TASK_PP(16'h410E,4);
TASK_PP(16'h410F,4);
TASK_PP(16'h4110,4);
TASK_PP(16'h4111,4);
TASK_PP(16'h4112,4);
TASK_PP(16'h4113,4);
TASK_PP(16'h4114,4);
TASK_PP(16'h4115,4);
TASK_PP(16'h4116,4);
TASK_PP(16'h4117,4);
TASK_PP(16'h4118,4);
TASK_PP(16'h4119,4);
TASK_PP(16'h411A,4);
TASK_PP(16'h411B,4);
TASK_PP(16'h411C,4);
TASK_PP(16'h411D,4);
TASK_PP(16'h411E,4);
TASK_PP(16'h411F,4);
TASK_PP(16'h4120,4);
TASK_PP(16'h4121,4);
TASK_PP(16'h4122,4);
TASK_PP(16'h4123,4);
TASK_PP(16'h4124,4);
TASK_PP(16'h4125,4);
TASK_PP(16'h4126,4);
TASK_PP(16'h4127,4);
TASK_PP(16'h4128,4);
TASK_PP(16'h4129,4);
TASK_PP(16'h412A,4);
TASK_PP(16'h412B,4);
TASK_PP(16'h412C,4);
TASK_PP(16'h412D,4);
TASK_PP(16'h412E,4);
TASK_PP(16'h412F,4);
TASK_PP(16'h4130,4);
TASK_PP(16'h4131,4);
TASK_PP(16'h4132,4);
TASK_PP(16'h4133,4);
TASK_PP(16'h4134,4);
TASK_PP(16'h4135,4);
TASK_PP(16'h4136,4);
TASK_PP(16'h4137,4);
TASK_PP(16'h4138,4);
TASK_PP(16'h4139,4);
TASK_PP(16'h413A,4);
TASK_PP(16'h413B,4);
TASK_PP(16'h413C,4);
TASK_PP(16'h413D,4);
TASK_PP(16'h413E,4);
TASK_PP(16'h413F,4);
TASK_PP(16'h4140,4);
TASK_PP(16'h4141,4);
TASK_PP(16'h4142,4);
TASK_PP(16'h4143,4);
TASK_PP(16'h4144,4);
TASK_PP(16'h4145,4);
TASK_PP(16'h4146,4);
TASK_PP(16'h4147,4);
TASK_PP(16'h4148,4);
TASK_PP(16'h4149,4);
TASK_PP(16'h414A,4);
TASK_PP(16'h414B,4);
TASK_PP(16'h414C,4);
TASK_PP(16'h414D,4);
TASK_PP(16'h414E,4);
TASK_PP(16'h414F,4);
TASK_PP(16'h4150,4);
TASK_PP(16'h4151,4);
TASK_PP(16'h4152,4);
TASK_PP(16'h4153,4);
TASK_PP(16'h4154,4);
TASK_PP(16'h4155,4);
TASK_PP(16'h4156,4);
TASK_PP(16'h4157,4);
TASK_PP(16'h4158,4);
TASK_PP(16'h4159,4);
TASK_PP(16'h415A,4);
TASK_PP(16'h415B,4);
TASK_PP(16'h415C,4);
TASK_PP(16'h415D,4);
TASK_PP(16'h415E,4);
TASK_PP(16'h415F,4);
TASK_PP(16'h4160,4);
TASK_PP(16'h4161,4);
TASK_PP(16'h4162,4);
TASK_PP(16'h4163,4);
TASK_PP(16'h4164,4);
TASK_PP(16'h4165,4);
TASK_PP(16'h4166,4);
TASK_PP(16'h4167,4);
TASK_PP(16'h4168,4);
TASK_PP(16'h4169,4);
TASK_PP(16'h416A,4);
TASK_PP(16'h416B,4);
TASK_PP(16'h416C,4);
TASK_PP(16'h416D,4);
TASK_PP(16'h416E,4);
TASK_PP(16'h416F,4);
TASK_PP(16'h4170,4);
TASK_PP(16'h4171,4);
TASK_PP(16'h4172,4);
TASK_PP(16'h4173,4);
TASK_PP(16'h4174,4);
TASK_PP(16'h4175,4);
TASK_PP(16'h4176,4);
TASK_PP(16'h4177,4);
TASK_PP(16'h4178,4);
TASK_PP(16'h4179,4);
TASK_PP(16'h417A,4);
TASK_PP(16'h417B,4);
TASK_PP(16'h417C,4);
TASK_PP(16'h417D,4);
TASK_PP(16'h417E,4);
TASK_PP(16'h417F,4);
TASK_PP(16'h4180,4);
TASK_PP(16'h4181,4);
TASK_PP(16'h4182,4);
TASK_PP(16'h4183,4);
TASK_PP(16'h4184,4);
TASK_PP(16'h4185,4);
TASK_PP(16'h4186,4);
TASK_PP(16'h4187,4);
TASK_PP(16'h4188,4);
TASK_PP(16'h4189,4);
TASK_PP(16'h418A,4);
TASK_PP(16'h418B,4);
TASK_PP(16'h418C,4);
TASK_PP(16'h418D,4);
TASK_PP(16'h418E,4);
TASK_PP(16'h418F,4);
TASK_PP(16'h4190,4);
TASK_PP(16'h4191,4);
TASK_PP(16'h4192,4);
TASK_PP(16'h4193,4);
TASK_PP(16'h4194,4);
TASK_PP(16'h4195,4);
TASK_PP(16'h4196,4);
TASK_PP(16'h4197,4);
TASK_PP(16'h4198,4);
TASK_PP(16'h4199,4);
TASK_PP(16'h419A,4);
TASK_PP(16'h419B,4);
TASK_PP(16'h419C,4);
TASK_PP(16'h419D,4);
TASK_PP(16'h419E,4);
TASK_PP(16'h419F,4);
TASK_PP(16'h41A0,4);
TASK_PP(16'h41A1,4);
TASK_PP(16'h41A2,4);
TASK_PP(16'h41A3,4);
TASK_PP(16'h41A4,4);
TASK_PP(16'h41A5,4);
TASK_PP(16'h41A6,4);
TASK_PP(16'h41A7,4);
TASK_PP(16'h41A8,4);
TASK_PP(16'h41A9,4);
TASK_PP(16'h41AA,4);
TASK_PP(16'h41AB,4);
TASK_PP(16'h41AC,4);
TASK_PP(16'h41AD,4);
TASK_PP(16'h41AE,4);
TASK_PP(16'h41AF,4);
TASK_PP(16'h41B0,4);
TASK_PP(16'h41B1,4);
TASK_PP(16'h41B2,4);
TASK_PP(16'h41B3,4);
TASK_PP(16'h41B4,4);
TASK_PP(16'h41B5,4);
TASK_PP(16'h41B6,4);
TASK_PP(16'h41B7,4);
TASK_PP(16'h41B8,4);
TASK_PP(16'h41B9,4);
TASK_PP(16'h41BA,4);
TASK_PP(16'h41BB,4);
TASK_PP(16'h41BC,4);
TASK_PP(16'h41BD,4);
TASK_PP(16'h41BE,4);
TASK_PP(16'h41BF,4);
TASK_PP(16'h41C0,4);
TASK_PP(16'h41C1,4);
TASK_PP(16'h41C2,4);
TASK_PP(16'h41C3,4);
TASK_PP(16'h41C4,4);
TASK_PP(16'h41C5,4);
TASK_PP(16'h41C6,4);
TASK_PP(16'h41C7,4);
TASK_PP(16'h41C8,4);
TASK_PP(16'h41C9,4);
TASK_PP(16'h41CA,4);
TASK_PP(16'h41CB,4);
TASK_PP(16'h41CC,4);
TASK_PP(16'h41CD,4);
TASK_PP(16'h41CE,4);
TASK_PP(16'h41CF,4);
TASK_PP(16'h41D0,4);
TASK_PP(16'h41D1,4);
TASK_PP(16'h41D2,4);
TASK_PP(16'h41D3,4);
TASK_PP(16'h41D4,4);
TASK_PP(16'h41D5,4);
TASK_PP(16'h41D6,4);
TASK_PP(16'h41D7,4);
TASK_PP(16'h41D8,4);
TASK_PP(16'h41D9,4);
TASK_PP(16'h41DA,4);
TASK_PP(16'h41DB,4);
TASK_PP(16'h41DC,4);
TASK_PP(16'h41DD,4);
TASK_PP(16'h41DE,4);
TASK_PP(16'h41DF,4);
TASK_PP(16'h41E0,4);
TASK_PP(16'h41E1,4);
TASK_PP(16'h41E2,4);
TASK_PP(16'h41E3,4);
TASK_PP(16'h41E4,4);
TASK_PP(16'h41E5,4);
TASK_PP(16'h41E6,4);
TASK_PP(16'h41E7,4);
TASK_PP(16'h41E8,4);
TASK_PP(16'h41E9,4);
TASK_PP(16'h41EA,4);
TASK_PP(16'h41EB,4);
TASK_PP(16'h41EC,4);
TASK_PP(16'h41ED,4);
TASK_PP(16'h41EE,4);
TASK_PP(16'h41EF,4);
TASK_PP(16'h41F0,4);
TASK_PP(16'h41F1,4);
TASK_PP(16'h41F2,4);
TASK_PP(16'h41F3,4);
TASK_PP(16'h41F4,4);
TASK_PP(16'h41F5,4);
TASK_PP(16'h41F6,4);
TASK_PP(16'h41F7,4);
TASK_PP(16'h41F8,4);
TASK_PP(16'h41F9,4);
TASK_PP(16'h41FA,4);
TASK_PP(16'h41FB,4);
TASK_PP(16'h41FC,4);
TASK_PP(16'h41FD,4);
TASK_PP(16'h41FE,4);
TASK_PP(16'h41FF,4);
TASK_PP(16'h4200,4);
TASK_PP(16'h4201,4);
TASK_PP(16'h4202,4);
TASK_PP(16'h4203,4);
TASK_PP(16'h4204,4);
TASK_PP(16'h4205,4);
TASK_PP(16'h4206,4);
TASK_PP(16'h4207,4);
TASK_PP(16'h4208,4);
TASK_PP(16'h4209,4);
TASK_PP(16'h420A,4);
TASK_PP(16'h420B,4);
TASK_PP(16'h420C,4);
TASK_PP(16'h420D,4);
TASK_PP(16'h420E,4);
TASK_PP(16'h420F,4);
TASK_PP(16'h4210,4);
TASK_PP(16'h4211,4);
TASK_PP(16'h4212,4);
TASK_PP(16'h4213,4);
TASK_PP(16'h4214,4);
TASK_PP(16'h4215,4);
TASK_PP(16'h4216,4);
TASK_PP(16'h4217,4);
TASK_PP(16'h4218,4);
TASK_PP(16'h4219,4);
TASK_PP(16'h421A,4);
TASK_PP(16'h421B,4);
TASK_PP(16'h421C,4);
TASK_PP(16'h421D,4);
TASK_PP(16'h421E,4);
TASK_PP(16'h421F,4);
TASK_PP(16'h4220,4);
TASK_PP(16'h4221,4);
TASK_PP(16'h4222,4);
TASK_PP(16'h4223,4);
TASK_PP(16'h4224,4);
TASK_PP(16'h4225,4);
TASK_PP(16'h4226,4);
TASK_PP(16'h4227,4);
TASK_PP(16'h4228,4);
TASK_PP(16'h4229,4);
TASK_PP(16'h422A,4);
TASK_PP(16'h422B,4);
TASK_PP(16'h422C,4);
TASK_PP(16'h422D,4);
TASK_PP(16'h422E,4);
TASK_PP(16'h422F,4);
TASK_PP(16'h4230,4);
TASK_PP(16'h4231,4);
TASK_PP(16'h4232,4);
TASK_PP(16'h4233,4);
TASK_PP(16'h4234,4);
TASK_PP(16'h4235,4);
TASK_PP(16'h4236,4);
TASK_PP(16'h4237,4);
TASK_PP(16'h4238,4);
TASK_PP(16'h4239,4);
TASK_PP(16'h423A,4);
TASK_PP(16'h423B,4);
TASK_PP(16'h423C,4);
TASK_PP(16'h423D,4);
TASK_PP(16'h423E,4);
TASK_PP(16'h423F,4);
TASK_PP(16'h4240,4);
TASK_PP(16'h4241,4);
TASK_PP(16'h4242,4);
TASK_PP(16'h4243,4);
TASK_PP(16'h4244,4);
TASK_PP(16'h4245,4);
TASK_PP(16'h4246,4);
TASK_PP(16'h4247,4);
TASK_PP(16'h4248,4);
TASK_PP(16'h4249,4);
TASK_PP(16'h424A,4);
TASK_PP(16'h424B,4);
TASK_PP(16'h424C,4);
TASK_PP(16'h424D,4);
TASK_PP(16'h424E,4);
TASK_PP(16'h424F,4);
TASK_PP(16'h4250,4);
TASK_PP(16'h4251,4);
TASK_PP(16'h4252,4);
TASK_PP(16'h4253,4);
TASK_PP(16'h4254,4);
TASK_PP(16'h4255,4);
TASK_PP(16'h4256,4);
TASK_PP(16'h4257,4);
TASK_PP(16'h4258,4);
TASK_PP(16'h4259,4);
TASK_PP(16'h425A,4);
TASK_PP(16'h425B,4);
TASK_PP(16'h425C,4);
TASK_PP(16'h425D,4);
TASK_PP(16'h425E,4);
TASK_PP(16'h425F,4);
TASK_PP(16'h4260,4);
TASK_PP(16'h4261,4);
TASK_PP(16'h4262,4);
TASK_PP(16'h4263,4);
TASK_PP(16'h4264,4);
TASK_PP(16'h4265,4);
TASK_PP(16'h4266,4);
TASK_PP(16'h4267,4);
TASK_PP(16'h4268,4);
TASK_PP(16'h4269,4);
TASK_PP(16'h426A,4);
TASK_PP(16'h426B,4);
TASK_PP(16'h426C,4);
TASK_PP(16'h426D,4);
TASK_PP(16'h426E,4);
TASK_PP(16'h426F,4);
TASK_PP(16'h4270,4);
TASK_PP(16'h4271,4);
TASK_PP(16'h4272,4);
TASK_PP(16'h4273,4);
TASK_PP(16'h4274,4);
TASK_PP(16'h4275,4);
TASK_PP(16'h4276,4);
TASK_PP(16'h4277,4);
TASK_PP(16'h4278,4);
TASK_PP(16'h4279,4);
TASK_PP(16'h427A,4);
TASK_PP(16'h427B,4);
TASK_PP(16'h427C,4);
TASK_PP(16'h427D,4);
TASK_PP(16'h427E,4);
TASK_PP(16'h427F,4);
TASK_PP(16'h4280,4);
TASK_PP(16'h4281,4);
TASK_PP(16'h4282,4);
TASK_PP(16'h4283,4);
TASK_PP(16'h4284,4);
TASK_PP(16'h4285,4);
TASK_PP(16'h4286,4);
TASK_PP(16'h4287,4);
TASK_PP(16'h4288,4);
TASK_PP(16'h4289,4);
TASK_PP(16'h428A,4);
TASK_PP(16'h428B,4);
TASK_PP(16'h428C,4);
TASK_PP(16'h428D,4);
TASK_PP(16'h428E,4);
TASK_PP(16'h428F,4);
TASK_PP(16'h4290,4);
TASK_PP(16'h4291,4);
TASK_PP(16'h4292,4);
TASK_PP(16'h4293,4);
TASK_PP(16'h4294,4);
TASK_PP(16'h4295,4);
TASK_PP(16'h4296,4);
TASK_PP(16'h4297,4);
TASK_PP(16'h4298,4);
TASK_PP(16'h4299,4);
TASK_PP(16'h429A,4);
TASK_PP(16'h429B,4);
TASK_PP(16'h429C,4);
TASK_PP(16'h429D,4);
TASK_PP(16'h429E,4);
TASK_PP(16'h429F,4);
TASK_PP(16'h42A0,4);
TASK_PP(16'h42A1,4);
TASK_PP(16'h42A2,4);
TASK_PP(16'h42A3,4);
TASK_PP(16'h42A4,4);
TASK_PP(16'h42A5,4);
TASK_PP(16'h42A6,4);
TASK_PP(16'h42A7,4);
TASK_PP(16'h42A8,4);
TASK_PP(16'h42A9,4);
TASK_PP(16'h42AA,4);
TASK_PP(16'h42AB,4);
TASK_PP(16'h42AC,4);
TASK_PP(16'h42AD,4);
TASK_PP(16'h42AE,4);
TASK_PP(16'h42AF,4);
TASK_PP(16'h42B0,4);
TASK_PP(16'h42B1,4);
TASK_PP(16'h42B2,4);
TASK_PP(16'h42B3,4);
TASK_PP(16'h42B4,4);
TASK_PP(16'h42B5,4);
TASK_PP(16'h42B6,4);
TASK_PP(16'h42B7,4);
TASK_PP(16'h42B8,4);
TASK_PP(16'h42B9,4);
TASK_PP(16'h42BA,4);
TASK_PP(16'h42BB,4);
TASK_PP(16'h42BC,4);
TASK_PP(16'h42BD,4);
TASK_PP(16'h42BE,4);
TASK_PP(16'h42BF,4);
TASK_PP(16'h42C0,4);
TASK_PP(16'h42C1,4);
TASK_PP(16'h42C2,4);
TASK_PP(16'h42C3,4);
TASK_PP(16'h42C4,4);
TASK_PP(16'h42C5,4);
TASK_PP(16'h42C6,4);
TASK_PP(16'h42C7,4);
TASK_PP(16'h42C8,4);
TASK_PP(16'h42C9,4);
TASK_PP(16'h42CA,4);
TASK_PP(16'h42CB,4);
TASK_PP(16'h42CC,4);
TASK_PP(16'h42CD,4);
TASK_PP(16'h42CE,4);
TASK_PP(16'h42CF,4);
TASK_PP(16'h42D0,4);
TASK_PP(16'h42D1,4);
TASK_PP(16'h42D2,4);
TASK_PP(16'h42D3,4);
TASK_PP(16'h42D4,4);
TASK_PP(16'h42D5,4);
TASK_PP(16'h42D6,4);
TASK_PP(16'h42D7,4);
TASK_PP(16'h42D8,4);
TASK_PP(16'h42D9,4);
TASK_PP(16'h42DA,4);
TASK_PP(16'h42DB,4);
TASK_PP(16'h42DC,4);
TASK_PP(16'h42DD,4);
TASK_PP(16'h42DE,4);
TASK_PP(16'h42DF,4);
TASK_PP(16'h42E0,4);
TASK_PP(16'h42E1,4);
TASK_PP(16'h42E2,4);
TASK_PP(16'h42E3,4);
TASK_PP(16'h42E4,4);
TASK_PP(16'h42E5,4);
TASK_PP(16'h42E6,4);
TASK_PP(16'h42E7,4);
TASK_PP(16'h42E8,4);
TASK_PP(16'h42E9,4);
TASK_PP(16'h42EA,4);
TASK_PP(16'h42EB,4);
TASK_PP(16'h42EC,4);
TASK_PP(16'h42ED,4);
TASK_PP(16'h42EE,4);
TASK_PP(16'h42EF,4);
TASK_PP(16'h42F0,4);
TASK_PP(16'h42F1,4);
TASK_PP(16'h42F2,4);
TASK_PP(16'h42F3,4);
TASK_PP(16'h42F4,4);
TASK_PP(16'h42F5,4);
TASK_PP(16'h42F6,4);
TASK_PP(16'h42F7,4);
TASK_PP(16'h42F8,4);
TASK_PP(16'h42F9,4);
TASK_PP(16'h42FA,4);
TASK_PP(16'h42FB,4);
TASK_PP(16'h42FC,4);
TASK_PP(16'h42FD,4);
TASK_PP(16'h42FE,4);
TASK_PP(16'h42FF,4);
TASK_PP(16'h4300,4);
TASK_PP(16'h4301,4);
TASK_PP(16'h4302,4);
TASK_PP(16'h4303,4);
TASK_PP(16'h4304,4);
TASK_PP(16'h4305,4);
TASK_PP(16'h4306,4);
TASK_PP(16'h4307,4);
TASK_PP(16'h4308,4);
TASK_PP(16'h4309,4);
TASK_PP(16'h430A,4);
TASK_PP(16'h430B,4);
TASK_PP(16'h430C,4);
TASK_PP(16'h430D,4);
TASK_PP(16'h430E,4);
TASK_PP(16'h430F,4);
TASK_PP(16'h4310,4);
TASK_PP(16'h4311,4);
TASK_PP(16'h4312,4);
TASK_PP(16'h4313,4);
TASK_PP(16'h4314,4);
TASK_PP(16'h4315,4);
TASK_PP(16'h4316,4);
TASK_PP(16'h4317,4);
TASK_PP(16'h4318,4);
TASK_PP(16'h4319,4);
TASK_PP(16'h431A,4);
TASK_PP(16'h431B,4);
TASK_PP(16'h431C,4);
TASK_PP(16'h431D,4);
TASK_PP(16'h431E,4);
TASK_PP(16'h431F,4);
TASK_PP(16'h4320,4);
TASK_PP(16'h4321,4);
TASK_PP(16'h4322,4);
TASK_PP(16'h4323,4);
TASK_PP(16'h4324,4);
TASK_PP(16'h4325,4);
TASK_PP(16'h4326,4);
TASK_PP(16'h4327,4);
TASK_PP(16'h4328,4);
TASK_PP(16'h4329,4);
TASK_PP(16'h432A,4);
TASK_PP(16'h432B,4);
TASK_PP(16'h432C,4);
TASK_PP(16'h432D,4);
TASK_PP(16'h432E,4);
TASK_PP(16'h432F,4);
TASK_PP(16'h4330,4);
TASK_PP(16'h4331,4);
TASK_PP(16'h4332,4);
TASK_PP(16'h4333,4);
TASK_PP(16'h4334,4);
TASK_PP(16'h4335,4);
TASK_PP(16'h4336,4);
TASK_PP(16'h4337,4);
TASK_PP(16'h4338,4);
TASK_PP(16'h4339,4);
TASK_PP(16'h433A,4);
TASK_PP(16'h433B,4);
TASK_PP(16'h433C,4);
TASK_PP(16'h433D,4);
TASK_PP(16'h433E,4);
TASK_PP(16'h433F,4);
TASK_PP(16'h4340,4);
TASK_PP(16'h4341,4);
TASK_PP(16'h4342,4);
TASK_PP(16'h4343,4);
TASK_PP(16'h4344,4);
TASK_PP(16'h4345,4);
TASK_PP(16'h4346,4);
TASK_PP(16'h4347,4);
TASK_PP(16'h4348,4);
TASK_PP(16'h4349,4);
TASK_PP(16'h434A,4);
TASK_PP(16'h434B,4);
TASK_PP(16'h434C,4);
TASK_PP(16'h434D,4);
TASK_PP(16'h434E,4);
TASK_PP(16'h434F,4);
TASK_PP(16'h4350,4);
TASK_PP(16'h4351,4);
TASK_PP(16'h4352,4);
TASK_PP(16'h4353,4);
TASK_PP(16'h4354,4);
TASK_PP(16'h4355,4);
TASK_PP(16'h4356,4);
TASK_PP(16'h4357,4);
TASK_PP(16'h4358,4);
TASK_PP(16'h4359,4);
TASK_PP(16'h435A,4);
TASK_PP(16'h435B,4);
TASK_PP(16'h435C,4);
TASK_PP(16'h435D,4);
TASK_PP(16'h435E,4);
TASK_PP(16'h435F,4);
TASK_PP(16'h4360,4);
TASK_PP(16'h4361,4);
TASK_PP(16'h4362,4);
TASK_PP(16'h4363,4);
TASK_PP(16'h4364,4);
TASK_PP(16'h4365,4);
TASK_PP(16'h4366,4);
TASK_PP(16'h4367,4);
TASK_PP(16'h4368,4);
TASK_PP(16'h4369,4);
TASK_PP(16'h436A,4);
TASK_PP(16'h436B,4);
TASK_PP(16'h436C,4);
TASK_PP(16'h436D,4);
TASK_PP(16'h436E,4);
TASK_PP(16'h436F,4);
TASK_PP(16'h4370,4);
TASK_PP(16'h4371,4);
TASK_PP(16'h4372,4);
TASK_PP(16'h4373,4);
TASK_PP(16'h4374,4);
TASK_PP(16'h4375,4);
TASK_PP(16'h4376,4);
TASK_PP(16'h4377,4);
TASK_PP(16'h4378,4);
TASK_PP(16'h4379,4);
TASK_PP(16'h437A,4);
TASK_PP(16'h437B,4);
TASK_PP(16'h437C,4);
TASK_PP(16'h437D,4);
TASK_PP(16'h437E,4);
TASK_PP(16'h437F,4);
TASK_PP(16'h4380,4);
TASK_PP(16'h4381,4);
TASK_PP(16'h4382,4);
TASK_PP(16'h4383,4);
TASK_PP(16'h4384,4);
TASK_PP(16'h4385,4);
TASK_PP(16'h4386,4);
TASK_PP(16'h4387,4);
TASK_PP(16'h4388,4);
TASK_PP(16'h4389,4);
TASK_PP(16'h438A,4);
TASK_PP(16'h438B,4);
TASK_PP(16'h438C,4);
TASK_PP(16'h438D,4);
TASK_PP(16'h438E,4);
TASK_PP(16'h438F,4);
TASK_PP(16'h4390,4);
TASK_PP(16'h4391,4);
TASK_PP(16'h4392,4);
TASK_PP(16'h4393,4);
TASK_PP(16'h4394,4);
TASK_PP(16'h4395,4);
TASK_PP(16'h4396,4);
TASK_PP(16'h4397,4);
TASK_PP(16'h4398,4);
TASK_PP(16'h4399,4);
TASK_PP(16'h439A,4);
TASK_PP(16'h439B,4);
TASK_PP(16'h439C,4);
TASK_PP(16'h439D,4);
TASK_PP(16'h439E,4);
TASK_PP(16'h439F,4);
TASK_PP(16'h43A0,4);
TASK_PP(16'h43A1,4);
TASK_PP(16'h43A2,4);
TASK_PP(16'h43A3,4);
TASK_PP(16'h43A4,4);
TASK_PP(16'h43A5,4);
TASK_PP(16'h43A6,4);
TASK_PP(16'h43A7,4);
TASK_PP(16'h43A8,4);
TASK_PP(16'h43A9,4);
TASK_PP(16'h43AA,4);
TASK_PP(16'h43AB,4);
TASK_PP(16'h43AC,4);
TASK_PP(16'h43AD,4);
TASK_PP(16'h43AE,4);
TASK_PP(16'h43AF,4);
TASK_PP(16'h43B0,4);
TASK_PP(16'h43B1,4);
TASK_PP(16'h43B2,4);
TASK_PP(16'h43B3,4);
TASK_PP(16'h43B4,4);
TASK_PP(16'h43B5,4);
TASK_PP(16'h43B6,4);
TASK_PP(16'h43B7,4);
TASK_PP(16'h43B8,4);
TASK_PP(16'h43B9,4);
TASK_PP(16'h43BA,4);
TASK_PP(16'h43BB,4);
TASK_PP(16'h43BC,4);
TASK_PP(16'h43BD,4);
TASK_PP(16'h43BE,4);
TASK_PP(16'h43BF,4);
TASK_PP(16'h43C0,4);
TASK_PP(16'h43C1,4);
TASK_PP(16'h43C2,4);
TASK_PP(16'h43C3,4);
TASK_PP(16'h43C4,4);
TASK_PP(16'h43C5,4);
TASK_PP(16'h43C6,4);
TASK_PP(16'h43C7,4);
TASK_PP(16'h43C8,4);
TASK_PP(16'h43C9,4);
TASK_PP(16'h43CA,4);
TASK_PP(16'h43CB,4);
TASK_PP(16'h43CC,4);
TASK_PP(16'h43CD,4);
TASK_PP(16'h43CE,4);
TASK_PP(16'h43CF,4);
TASK_PP(16'h43D0,4);
TASK_PP(16'h43D1,4);
TASK_PP(16'h43D2,4);
TASK_PP(16'h43D3,4);
TASK_PP(16'h43D4,4);
TASK_PP(16'h43D5,4);
TASK_PP(16'h43D6,4);
TASK_PP(16'h43D7,4);
TASK_PP(16'h43D8,4);
TASK_PP(16'h43D9,4);
TASK_PP(16'h43DA,4);
TASK_PP(16'h43DB,4);
TASK_PP(16'h43DC,4);
TASK_PP(16'h43DD,4);
TASK_PP(16'h43DE,4);
TASK_PP(16'h43DF,4);
TASK_PP(16'h43E0,4);
TASK_PP(16'h43E1,4);
TASK_PP(16'h43E2,4);
TASK_PP(16'h43E3,4);
TASK_PP(16'h43E4,4);
TASK_PP(16'h43E5,4);
TASK_PP(16'h43E6,4);
TASK_PP(16'h43E7,4);
TASK_PP(16'h43E8,4);
TASK_PP(16'h43E9,4);
TASK_PP(16'h43EA,4);
TASK_PP(16'h43EB,4);
TASK_PP(16'h43EC,4);
TASK_PP(16'h43ED,4);
TASK_PP(16'h43EE,4);
TASK_PP(16'h43EF,4);
TASK_PP(16'h43F0,4);
TASK_PP(16'h43F1,4);
TASK_PP(16'h43F2,4);
TASK_PP(16'h43F3,4);
TASK_PP(16'h43F4,4);
TASK_PP(16'h43F5,4);
TASK_PP(16'h43F6,4);
TASK_PP(16'h43F7,4);
TASK_PP(16'h43F8,4);
TASK_PP(16'h43F9,4);
TASK_PP(16'h43FA,4);
TASK_PP(16'h43FB,4);
TASK_PP(16'h43FC,4);
TASK_PP(16'h43FD,4);
TASK_PP(16'h43FE,4);
TASK_PP(16'h43FF,4);
TASK_PP(16'h4400,4);
TASK_PP(16'h4401,4);
TASK_PP(16'h4402,4);
TASK_PP(16'h4403,4);
TASK_PP(16'h4404,4);
TASK_PP(16'h4405,4);
TASK_PP(16'h4406,4);
TASK_PP(16'h4407,4);
TASK_PP(16'h4408,4);
TASK_PP(16'h4409,4);
TASK_PP(16'h440A,4);
TASK_PP(16'h440B,4);
TASK_PP(16'h440C,4);
TASK_PP(16'h440D,4);
TASK_PP(16'h440E,4);
TASK_PP(16'h440F,4);
TASK_PP(16'h4410,4);
TASK_PP(16'h4411,4);
TASK_PP(16'h4412,4);
TASK_PP(16'h4413,4);
TASK_PP(16'h4414,4);
TASK_PP(16'h4415,4);
TASK_PP(16'h4416,4);
TASK_PP(16'h4417,4);
TASK_PP(16'h4418,4);
TASK_PP(16'h4419,4);
TASK_PP(16'h441A,4);
TASK_PP(16'h441B,4);
TASK_PP(16'h441C,4);
TASK_PP(16'h441D,4);
TASK_PP(16'h441E,4);
TASK_PP(16'h441F,4);
TASK_PP(16'h4420,4);
TASK_PP(16'h4421,4);
TASK_PP(16'h4422,4);
TASK_PP(16'h4423,4);
TASK_PP(16'h4424,4);
TASK_PP(16'h4425,4);
TASK_PP(16'h4426,4);
TASK_PP(16'h4427,4);
TASK_PP(16'h4428,4);
TASK_PP(16'h4429,4);
TASK_PP(16'h442A,4);
TASK_PP(16'h442B,4);
TASK_PP(16'h442C,4);
TASK_PP(16'h442D,4);
TASK_PP(16'h442E,4);
TASK_PP(16'h442F,4);
TASK_PP(16'h4430,4);
TASK_PP(16'h4431,4);
TASK_PP(16'h4432,4);
TASK_PP(16'h4433,4);
TASK_PP(16'h4434,4);
TASK_PP(16'h4435,4);
TASK_PP(16'h4436,4);
TASK_PP(16'h4437,4);
TASK_PP(16'h4438,4);
TASK_PP(16'h4439,4);
TASK_PP(16'h443A,4);
TASK_PP(16'h443B,4);
TASK_PP(16'h443C,4);
TASK_PP(16'h443D,4);
TASK_PP(16'h443E,4);
TASK_PP(16'h443F,4);
TASK_PP(16'h4440,4);
TASK_PP(16'h4441,4);
TASK_PP(16'h4442,4);
TASK_PP(16'h4443,4);
TASK_PP(16'h4444,4);
TASK_PP(16'h4445,4);
TASK_PP(16'h4446,4);
TASK_PP(16'h4447,4);
TASK_PP(16'h4448,4);
TASK_PP(16'h4449,4);
TASK_PP(16'h444A,4);
TASK_PP(16'h444B,4);
TASK_PP(16'h444C,4);
TASK_PP(16'h444D,4);
TASK_PP(16'h444E,4);
TASK_PP(16'h444F,4);
TASK_PP(16'h4450,4);
TASK_PP(16'h4451,4);
TASK_PP(16'h4452,4);
TASK_PP(16'h4453,4);
TASK_PP(16'h4454,4);
TASK_PP(16'h4455,4);
TASK_PP(16'h4456,4);
TASK_PP(16'h4457,4);
TASK_PP(16'h4458,4);
TASK_PP(16'h4459,4);
TASK_PP(16'h445A,4);
TASK_PP(16'h445B,4);
TASK_PP(16'h445C,4);
TASK_PP(16'h445D,4);
TASK_PP(16'h445E,4);
TASK_PP(16'h445F,4);
TASK_PP(16'h4460,4);
TASK_PP(16'h4461,4);
TASK_PP(16'h4462,4);
TASK_PP(16'h4463,4);
TASK_PP(16'h4464,4);
TASK_PP(16'h4465,4);
TASK_PP(16'h4466,4);
TASK_PP(16'h4467,4);
TASK_PP(16'h4468,4);
TASK_PP(16'h4469,4);
TASK_PP(16'h446A,4);
TASK_PP(16'h446B,4);
TASK_PP(16'h446C,4);
TASK_PP(16'h446D,4);
TASK_PP(16'h446E,4);
TASK_PP(16'h446F,4);
TASK_PP(16'h4470,4);
TASK_PP(16'h4471,4);
TASK_PP(16'h4472,4);
TASK_PP(16'h4473,4);
TASK_PP(16'h4474,4);
TASK_PP(16'h4475,4);
TASK_PP(16'h4476,4);
TASK_PP(16'h4477,4);
TASK_PP(16'h4478,4);
TASK_PP(16'h4479,4);
TASK_PP(16'h447A,4);
TASK_PP(16'h447B,4);
TASK_PP(16'h447C,4);
TASK_PP(16'h447D,4);
TASK_PP(16'h447E,4);
TASK_PP(16'h447F,4);
TASK_PP(16'h4480,4);
TASK_PP(16'h4481,4);
TASK_PP(16'h4482,4);
TASK_PP(16'h4483,4);
TASK_PP(16'h4484,4);
TASK_PP(16'h4485,4);
TASK_PP(16'h4486,4);
TASK_PP(16'h4487,4);
TASK_PP(16'h4488,4);
TASK_PP(16'h4489,4);
TASK_PP(16'h448A,4);
TASK_PP(16'h448B,4);
TASK_PP(16'h448C,4);
TASK_PP(16'h448D,4);
TASK_PP(16'h448E,4);
TASK_PP(16'h448F,4);
TASK_PP(16'h4490,4);
TASK_PP(16'h4491,4);
TASK_PP(16'h4492,4);
TASK_PP(16'h4493,4);
TASK_PP(16'h4494,4);
TASK_PP(16'h4495,4);
TASK_PP(16'h4496,4);
TASK_PP(16'h4497,4);
TASK_PP(16'h4498,4);
TASK_PP(16'h4499,4);
TASK_PP(16'h449A,4);
TASK_PP(16'h449B,4);
TASK_PP(16'h449C,4);
TASK_PP(16'h449D,4);
TASK_PP(16'h449E,4);
TASK_PP(16'h449F,4);
TASK_PP(16'h44A0,4);
TASK_PP(16'h44A1,4);
TASK_PP(16'h44A2,4);
TASK_PP(16'h44A3,4);
TASK_PP(16'h44A4,4);
TASK_PP(16'h44A5,4);
TASK_PP(16'h44A6,4);
TASK_PP(16'h44A7,4);
TASK_PP(16'h44A8,4);
TASK_PP(16'h44A9,4);
TASK_PP(16'h44AA,4);
TASK_PP(16'h44AB,4);
TASK_PP(16'h44AC,4);
TASK_PP(16'h44AD,4);
TASK_PP(16'h44AE,4);
TASK_PP(16'h44AF,4);
TASK_PP(16'h44B0,4);
TASK_PP(16'h44B1,4);
TASK_PP(16'h44B2,4);
TASK_PP(16'h44B3,4);
TASK_PP(16'h44B4,4);
TASK_PP(16'h44B5,4);
TASK_PP(16'h44B6,4);
TASK_PP(16'h44B7,4);
TASK_PP(16'h44B8,4);
TASK_PP(16'h44B9,4);
TASK_PP(16'h44BA,4);
TASK_PP(16'h44BB,4);
TASK_PP(16'h44BC,4);
TASK_PP(16'h44BD,4);
TASK_PP(16'h44BE,4);
TASK_PP(16'h44BF,4);
TASK_PP(16'h44C0,4);
TASK_PP(16'h44C1,4);
TASK_PP(16'h44C2,4);
TASK_PP(16'h44C3,4);
TASK_PP(16'h44C4,4);
TASK_PP(16'h44C5,4);
TASK_PP(16'h44C6,4);
TASK_PP(16'h44C7,4);
TASK_PP(16'h44C8,4);
TASK_PP(16'h44C9,4);
TASK_PP(16'h44CA,4);
TASK_PP(16'h44CB,4);
TASK_PP(16'h44CC,4);
TASK_PP(16'h44CD,4);
TASK_PP(16'h44CE,4);
TASK_PP(16'h44CF,4);
TASK_PP(16'h44D0,4);
TASK_PP(16'h44D1,4);
TASK_PP(16'h44D2,4);
TASK_PP(16'h44D3,4);
TASK_PP(16'h44D4,4);
TASK_PP(16'h44D5,4);
TASK_PP(16'h44D6,4);
TASK_PP(16'h44D7,4);
TASK_PP(16'h44D8,4);
TASK_PP(16'h44D9,4);
TASK_PP(16'h44DA,4);
TASK_PP(16'h44DB,4);
TASK_PP(16'h44DC,4);
TASK_PP(16'h44DD,4);
TASK_PP(16'h44DE,4);
TASK_PP(16'h44DF,4);
TASK_PP(16'h44E0,4);
TASK_PP(16'h44E1,4);
TASK_PP(16'h44E2,4);
TASK_PP(16'h44E3,4);
TASK_PP(16'h44E4,4);
TASK_PP(16'h44E5,4);
TASK_PP(16'h44E6,4);
TASK_PP(16'h44E7,4);
TASK_PP(16'h44E8,4);
TASK_PP(16'h44E9,4);
TASK_PP(16'h44EA,4);
TASK_PP(16'h44EB,4);
TASK_PP(16'h44EC,4);
TASK_PP(16'h44ED,4);
TASK_PP(16'h44EE,4);
TASK_PP(16'h44EF,4);
TASK_PP(16'h44F0,4);
TASK_PP(16'h44F1,4);
TASK_PP(16'h44F2,4);
TASK_PP(16'h44F3,4);
TASK_PP(16'h44F4,4);
TASK_PP(16'h44F5,4);
TASK_PP(16'h44F6,4);
TASK_PP(16'h44F7,4);
TASK_PP(16'h44F8,4);
TASK_PP(16'h44F9,4);
TASK_PP(16'h44FA,4);
TASK_PP(16'h44FB,4);
TASK_PP(16'h44FC,4);
TASK_PP(16'h44FD,4);
TASK_PP(16'h44FE,4);
TASK_PP(16'h44FF,4);
TASK_PP(16'h4500,4);
TASK_PP(16'h4501,4);
TASK_PP(16'h4502,4);
TASK_PP(16'h4503,4);
TASK_PP(16'h4504,4);
TASK_PP(16'h4505,4);
TASK_PP(16'h4506,4);
TASK_PP(16'h4507,4);
TASK_PP(16'h4508,4);
TASK_PP(16'h4509,4);
TASK_PP(16'h450A,4);
TASK_PP(16'h450B,4);
TASK_PP(16'h450C,4);
TASK_PP(16'h450D,4);
TASK_PP(16'h450E,4);
TASK_PP(16'h450F,4);
TASK_PP(16'h4510,4);
TASK_PP(16'h4511,4);
TASK_PP(16'h4512,4);
TASK_PP(16'h4513,4);
TASK_PP(16'h4514,4);
TASK_PP(16'h4515,4);
TASK_PP(16'h4516,4);
TASK_PP(16'h4517,4);
TASK_PP(16'h4518,4);
TASK_PP(16'h4519,4);
TASK_PP(16'h451A,4);
TASK_PP(16'h451B,4);
TASK_PP(16'h451C,4);
TASK_PP(16'h451D,4);
TASK_PP(16'h451E,4);
TASK_PP(16'h451F,4);
TASK_PP(16'h4520,4);
TASK_PP(16'h4521,4);
TASK_PP(16'h4522,4);
TASK_PP(16'h4523,4);
TASK_PP(16'h4524,4);
TASK_PP(16'h4525,4);
TASK_PP(16'h4526,4);
TASK_PP(16'h4527,4);
TASK_PP(16'h4528,4);
TASK_PP(16'h4529,4);
TASK_PP(16'h452A,4);
TASK_PP(16'h452B,4);
TASK_PP(16'h452C,4);
TASK_PP(16'h452D,4);
TASK_PP(16'h452E,4);
TASK_PP(16'h452F,4);
TASK_PP(16'h4530,4);
TASK_PP(16'h4531,4);
TASK_PP(16'h4532,4);
TASK_PP(16'h4533,4);
TASK_PP(16'h4534,4);
TASK_PP(16'h4535,4);
TASK_PP(16'h4536,4);
TASK_PP(16'h4537,4);
TASK_PP(16'h4538,4);
TASK_PP(16'h4539,4);
TASK_PP(16'h453A,4);
TASK_PP(16'h453B,4);
TASK_PP(16'h453C,4);
TASK_PP(16'h453D,4);
TASK_PP(16'h453E,4);
TASK_PP(16'h453F,4);
TASK_PP(16'h4540,4);
TASK_PP(16'h4541,4);
TASK_PP(16'h4542,4);
TASK_PP(16'h4543,4);
TASK_PP(16'h4544,4);
TASK_PP(16'h4545,4);
TASK_PP(16'h4546,4);
TASK_PP(16'h4547,4);
TASK_PP(16'h4548,4);
TASK_PP(16'h4549,4);
TASK_PP(16'h454A,4);
TASK_PP(16'h454B,4);
TASK_PP(16'h454C,4);
TASK_PP(16'h454D,4);
TASK_PP(16'h454E,4);
TASK_PP(16'h454F,4);
TASK_PP(16'h4550,4);
TASK_PP(16'h4551,4);
TASK_PP(16'h4552,4);
TASK_PP(16'h4553,4);
TASK_PP(16'h4554,4);
TASK_PP(16'h4555,4);
TASK_PP(16'h4556,4);
TASK_PP(16'h4557,4);
TASK_PP(16'h4558,4);
TASK_PP(16'h4559,4);
TASK_PP(16'h455A,4);
TASK_PP(16'h455B,4);
TASK_PP(16'h455C,4);
TASK_PP(16'h455D,4);
TASK_PP(16'h455E,4);
TASK_PP(16'h455F,4);
TASK_PP(16'h4560,4);
TASK_PP(16'h4561,4);
TASK_PP(16'h4562,4);
TASK_PP(16'h4563,4);
TASK_PP(16'h4564,4);
TASK_PP(16'h4565,4);
TASK_PP(16'h4566,4);
TASK_PP(16'h4567,4);
TASK_PP(16'h4568,4);
TASK_PP(16'h4569,4);
TASK_PP(16'h456A,4);
TASK_PP(16'h456B,4);
TASK_PP(16'h456C,4);
TASK_PP(16'h456D,4);
TASK_PP(16'h456E,4);
TASK_PP(16'h456F,4);
TASK_PP(16'h4570,4);
TASK_PP(16'h4571,4);
TASK_PP(16'h4572,4);
TASK_PP(16'h4573,4);
TASK_PP(16'h4574,4);
TASK_PP(16'h4575,4);
TASK_PP(16'h4576,4);
TASK_PP(16'h4577,4);
TASK_PP(16'h4578,4);
TASK_PP(16'h4579,4);
TASK_PP(16'h457A,4);
TASK_PP(16'h457B,4);
TASK_PP(16'h457C,4);
TASK_PP(16'h457D,4);
TASK_PP(16'h457E,4);
TASK_PP(16'h457F,4);
TASK_PP(16'h4580,4);
TASK_PP(16'h4581,4);
TASK_PP(16'h4582,4);
TASK_PP(16'h4583,4);
TASK_PP(16'h4584,4);
TASK_PP(16'h4585,4);
TASK_PP(16'h4586,4);
TASK_PP(16'h4587,4);
TASK_PP(16'h4588,4);
TASK_PP(16'h4589,4);
TASK_PP(16'h458A,4);
TASK_PP(16'h458B,4);
TASK_PP(16'h458C,4);
TASK_PP(16'h458D,4);
TASK_PP(16'h458E,4);
TASK_PP(16'h458F,4);
TASK_PP(16'h4590,4);
TASK_PP(16'h4591,4);
TASK_PP(16'h4592,4);
TASK_PP(16'h4593,4);
TASK_PP(16'h4594,4);
TASK_PP(16'h4595,4);
TASK_PP(16'h4596,4);
TASK_PP(16'h4597,4);
TASK_PP(16'h4598,4);
TASK_PP(16'h4599,4);
TASK_PP(16'h459A,4);
TASK_PP(16'h459B,4);
TASK_PP(16'h459C,4);
TASK_PP(16'h459D,4);
TASK_PP(16'h459E,4);
TASK_PP(16'h459F,4);
TASK_PP(16'h45A0,4);
TASK_PP(16'h45A1,4);
TASK_PP(16'h45A2,4);
TASK_PP(16'h45A3,4);
TASK_PP(16'h45A4,4);
TASK_PP(16'h45A5,4);
TASK_PP(16'h45A6,4);
TASK_PP(16'h45A7,4);
TASK_PP(16'h45A8,4);
TASK_PP(16'h45A9,4);
TASK_PP(16'h45AA,4);
TASK_PP(16'h45AB,4);
TASK_PP(16'h45AC,4);
TASK_PP(16'h45AD,4);
TASK_PP(16'h45AE,4);
TASK_PP(16'h45AF,4);
TASK_PP(16'h45B0,4);
TASK_PP(16'h45B1,4);
TASK_PP(16'h45B2,4);
TASK_PP(16'h45B3,4);
TASK_PP(16'h45B4,4);
TASK_PP(16'h45B5,4);
TASK_PP(16'h45B6,4);
TASK_PP(16'h45B7,4);
TASK_PP(16'h45B8,4);
TASK_PP(16'h45B9,4);
TASK_PP(16'h45BA,4);
TASK_PP(16'h45BB,4);
TASK_PP(16'h45BC,4);
TASK_PP(16'h45BD,4);
TASK_PP(16'h45BE,4);
TASK_PP(16'h45BF,4);
TASK_PP(16'h45C0,4);
TASK_PP(16'h45C1,4);
TASK_PP(16'h45C2,4);
TASK_PP(16'h45C3,4);
TASK_PP(16'h45C4,4);
TASK_PP(16'h45C5,4);
TASK_PP(16'h45C6,4);
TASK_PP(16'h45C7,4);
TASK_PP(16'h45C8,4);
TASK_PP(16'h45C9,4);
TASK_PP(16'h45CA,4);
TASK_PP(16'h45CB,4);
TASK_PP(16'h45CC,4);
TASK_PP(16'h45CD,4);
TASK_PP(16'h45CE,4);
TASK_PP(16'h45CF,4);
TASK_PP(16'h45D0,4);
TASK_PP(16'h45D1,4);
TASK_PP(16'h45D2,4);
TASK_PP(16'h45D3,4);
TASK_PP(16'h45D4,4);
TASK_PP(16'h45D5,4);
TASK_PP(16'h45D6,4);
TASK_PP(16'h45D7,4);
TASK_PP(16'h45D8,4);
TASK_PP(16'h45D9,4);
TASK_PP(16'h45DA,4);
TASK_PP(16'h45DB,4);
TASK_PP(16'h45DC,4);
TASK_PP(16'h45DD,4);
TASK_PP(16'h45DE,4);
TASK_PP(16'h45DF,4);
TASK_PP(16'h45E0,4);
TASK_PP(16'h45E1,4);
TASK_PP(16'h45E2,4);
TASK_PP(16'h45E3,4);
TASK_PP(16'h45E4,4);
TASK_PP(16'h45E5,4);
TASK_PP(16'h45E6,4);
TASK_PP(16'h45E7,4);
TASK_PP(16'h45E8,4);
TASK_PP(16'h45E9,4);
TASK_PP(16'h45EA,4);
TASK_PP(16'h45EB,4);
TASK_PP(16'h45EC,4);
TASK_PP(16'h45ED,4);
TASK_PP(16'h45EE,4);
TASK_PP(16'h45EF,4);
TASK_PP(16'h45F0,4);
TASK_PP(16'h45F1,4);
TASK_PP(16'h45F2,4);
TASK_PP(16'h45F3,4);
TASK_PP(16'h45F4,4);
TASK_PP(16'h45F5,4);
TASK_PP(16'h45F6,4);
TASK_PP(16'h45F7,4);
TASK_PP(16'h45F8,4);
TASK_PP(16'h45F9,4);
TASK_PP(16'h45FA,4);
TASK_PP(16'h45FB,4);
TASK_PP(16'h45FC,4);
TASK_PP(16'h45FD,4);
TASK_PP(16'h45FE,4);
TASK_PP(16'h45FF,4);
TASK_PP(16'h4600,4);
TASK_PP(16'h4601,4);
TASK_PP(16'h4602,4);
TASK_PP(16'h4603,4);
TASK_PP(16'h4604,4);
TASK_PP(16'h4605,4);
TASK_PP(16'h4606,4);
TASK_PP(16'h4607,4);
TASK_PP(16'h4608,4);
TASK_PP(16'h4609,4);
TASK_PP(16'h460A,4);
TASK_PP(16'h460B,4);
TASK_PP(16'h460C,4);
TASK_PP(16'h460D,4);
TASK_PP(16'h460E,4);
TASK_PP(16'h460F,4);
TASK_PP(16'h4610,4);
TASK_PP(16'h4611,4);
TASK_PP(16'h4612,4);
TASK_PP(16'h4613,4);
TASK_PP(16'h4614,4);
TASK_PP(16'h4615,4);
TASK_PP(16'h4616,4);
TASK_PP(16'h4617,4);
TASK_PP(16'h4618,4);
TASK_PP(16'h4619,4);
TASK_PP(16'h461A,4);
TASK_PP(16'h461B,4);
TASK_PP(16'h461C,4);
TASK_PP(16'h461D,4);
TASK_PP(16'h461E,4);
TASK_PP(16'h461F,4);
TASK_PP(16'h4620,4);
TASK_PP(16'h4621,4);
TASK_PP(16'h4622,4);
TASK_PP(16'h4623,4);
TASK_PP(16'h4624,4);
TASK_PP(16'h4625,4);
TASK_PP(16'h4626,4);
TASK_PP(16'h4627,4);
TASK_PP(16'h4628,4);
TASK_PP(16'h4629,4);
TASK_PP(16'h462A,4);
TASK_PP(16'h462B,4);
TASK_PP(16'h462C,4);
TASK_PP(16'h462D,4);
TASK_PP(16'h462E,4);
TASK_PP(16'h462F,4);
TASK_PP(16'h4630,4);
TASK_PP(16'h4631,4);
TASK_PP(16'h4632,4);
TASK_PP(16'h4633,4);
TASK_PP(16'h4634,4);
TASK_PP(16'h4635,4);
TASK_PP(16'h4636,4);
TASK_PP(16'h4637,4);
TASK_PP(16'h4638,4);
TASK_PP(16'h4639,4);
TASK_PP(16'h463A,4);
TASK_PP(16'h463B,4);
TASK_PP(16'h463C,4);
TASK_PP(16'h463D,4);
TASK_PP(16'h463E,4);
TASK_PP(16'h463F,4);
TASK_PP(16'h4640,4);
TASK_PP(16'h4641,4);
TASK_PP(16'h4642,4);
TASK_PP(16'h4643,4);
TASK_PP(16'h4644,4);
TASK_PP(16'h4645,4);
TASK_PP(16'h4646,4);
TASK_PP(16'h4647,4);
TASK_PP(16'h4648,4);
TASK_PP(16'h4649,4);
TASK_PP(16'h464A,4);
TASK_PP(16'h464B,4);
TASK_PP(16'h464C,4);
TASK_PP(16'h464D,4);
TASK_PP(16'h464E,4);
TASK_PP(16'h464F,4);
TASK_PP(16'h4650,4);
TASK_PP(16'h4651,4);
TASK_PP(16'h4652,4);
TASK_PP(16'h4653,4);
TASK_PP(16'h4654,4);
TASK_PP(16'h4655,4);
TASK_PP(16'h4656,4);
TASK_PP(16'h4657,4);
TASK_PP(16'h4658,4);
TASK_PP(16'h4659,4);
TASK_PP(16'h465A,4);
TASK_PP(16'h465B,4);
TASK_PP(16'h465C,4);
TASK_PP(16'h465D,4);
TASK_PP(16'h465E,4);
TASK_PP(16'h465F,4);
TASK_PP(16'h4660,4);
TASK_PP(16'h4661,4);
TASK_PP(16'h4662,4);
TASK_PP(16'h4663,4);
TASK_PP(16'h4664,4);
TASK_PP(16'h4665,4);
TASK_PP(16'h4666,4);
TASK_PP(16'h4667,4);
TASK_PP(16'h4668,4);
TASK_PP(16'h4669,4);
TASK_PP(16'h466A,4);
TASK_PP(16'h466B,4);
TASK_PP(16'h466C,4);
TASK_PP(16'h466D,4);
TASK_PP(16'h466E,4);
TASK_PP(16'h466F,4);
TASK_PP(16'h4670,4);
TASK_PP(16'h4671,4);
TASK_PP(16'h4672,4);
TASK_PP(16'h4673,4);
TASK_PP(16'h4674,4);
TASK_PP(16'h4675,4);
TASK_PP(16'h4676,4);
TASK_PP(16'h4677,4);
TASK_PP(16'h4678,4);
TASK_PP(16'h4679,4);
TASK_PP(16'h467A,4);
TASK_PP(16'h467B,4);
TASK_PP(16'h467C,4);
TASK_PP(16'h467D,4);
TASK_PP(16'h467E,4);
TASK_PP(16'h467F,4);
TASK_PP(16'h4680,4);
TASK_PP(16'h4681,4);
TASK_PP(16'h4682,4);
TASK_PP(16'h4683,4);
TASK_PP(16'h4684,4);
TASK_PP(16'h4685,4);
TASK_PP(16'h4686,4);
TASK_PP(16'h4687,4);
TASK_PP(16'h4688,4);
TASK_PP(16'h4689,4);
TASK_PP(16'h468A,4);
TASK_PP(16'h468B,4);
TASK_PP(16'h468C,4);
TASK_PP(16'h468D,4);
TASK_PP(16'h468E,4);
TASK_PP(16'h468F,4);
TASK_PP(16'h4690,4);
TASK_PP(16'h4691,4);
TASK_PP(16'h4692,4);
TASK_PP(16'h4693,4);
TASK_PP(16'h4694,4);
TASK_PP(16'h4695,4);
TASK_PP(16'h4696,4);
TASK_PP(16'h4697,4);
TASK_PP(16'h4698,4);
TASK_PP(16'h4699,4);
TASK_PP(16'h469A,4);
TASK_PP(16'h469B,4);
TASK_PP(16'h469C,4);
TASK_PP(16'h469D,4);
TASK_PP(16'h469E,4);
TASK_PP(16'h469F,4);
TASK_PP(16'h46A0,4);
TASK_PP(16'h46A1,4);
TASK_PP(16'h46A2,4);
TASK_PP(16'h46A3,4);
TASK_PP(16'h46A4,4);
TASK_PP(16'h46A5,4);
TASK_PP(16'h46A6,4);
TASK_PP(16'h46A7,4);
TASK_PP(16'h46A8,4);
TASK_PP(16'h46A9,4);
TASK_PP(16'h46AA,4);
TASK_PP(16'h46AB,4);
TASK_PP(16'h46AC,4);
TASK_PP(16'h46AD,4);
TASK_PP(16'h46AE,4);
TASK_PP(16'h46AF,4);
TASK_PP(16'h46B0,4);
TASK_PP(16'h46B1,4);
TASK_PP(16'h46B2,4);
TASK_PP(16'h46B3,4);
TASK_PP(16'h46B4,4);
TASK_PP(16'h46B5,4);
TASK_PP(16'h46B6,4);
TASK_PP(16'h46B7,4);
TASK_PP(16'h46B8,4);
TASK_PP(16'h46B9,4);
TASK_PP(16'h46BA,4);
TASK_PP(16'h46BB,4);
TASK_PP(16'h46BC,4);
TASK_PP(16'h46BD,4);
TASK_PP(16'h46BE,4);
TASK_PP(16'h46BF,4);
TASK_PP(16'h46C0,4);
TASK_PP(16'h46C1,4);
TASK_PP(16'h46C2,4);
TASK_PP(16'h46C3,4);
TASK_PP(16'h46C4,4);
TASK_PP(16'h46C5,4);
TASK_PP(16'h46C6,4);
TASK_PP(16'h46C7,4);
TASK_PP(16'h46C8,4);
TASK_PP(16'h46C9,4);
TASK_PP(16'h46CA,4);
TASK_PP(16'h46CB,4);
TASK_PP(16'h46CC,4);
TASK_PP(16'h46CD,4);
TASK_PP(16'h46CE,4);
TASK_PP(16'h46CF,4);
TASK_PP(16'h46D0,4);
TASK_PP(16'h46D1,4);
TASK_PP(16'h46D2,4);
TASK_PP(16'h46D3,4);
TASK_PP(16'h46D4,4);
TASK_PP(16'h46D5,4);
TASK_PP(16'h46D6,4);
TASK_PP(16'h46D7,4);
TASK_PP(16'h46D8,4);
TASK_PP(16'h46D9,4);
TASK_PP(16'h46DA,4);
TASK_PP(16'h46DB,4);
TASK_PP(16'h46DC,4);
TASK_PP(16'h46DD,4);
TASK_PP(16'h46DE,4);
TASK_PP(16'h46DF,4);
TASK_PP(16'h46E0,4);
TASK_PP(16'h46E1,4);
TASK_PP(16'h46E2,4);
TASK_PP(16'h46E3,4);
TASK_PP(16'h46E4,4);
TASK_PP(16'h46E5,4);
TASK_PP(16'h46E6,4);
TASK_PP(16'h46E7,4);
TASK_PP(16'h46E8,4);
TASK_PP(16'h46E9,4);
TASK_PP(16'h46EA,4);
TASK_PP(16'h46EB,4);
TASK_PP(16'h46EC,4);
TASK_PP(16'h46ED,4);
TASK_PP(16'h46EE,4);
TASK_PP(16'h46EF,4);
TASK_PP(16'h46F0,4);
TASK_PP(16'h46F1,4);
TASK_PP(16'h46F2,4);
TASK_PP(16'h46F3,4);
TASK_PP(16'h46F4,4);
TASK_PP(16'h46F5,4);
TASK_PP(16'h46F6,4);
TASK_PP(16'h46F7,4);
TASK_PP(16'h46F8,4);
TASK_PP(16'h46F9,4);
TASK_PP(16'h46FA,4);
TASK_PP(16'h46FB,4);
TASK_PP(16'h46FC,4);
TASK_PP(16'h46FD,4);
TASK_PP(16'h46FE,4);
TASK_PP(16'h46FF,4);
TASK_PP(16'h4700,4);
TASK_PP(16'h4701,4);
TASK_PP(16'h4702,4);
TASK_PP(16'h4703,4);
TASK_PP(16'h4704,4);
TASK_PP(16'h4705,4);
TASK_PP(16'h4706,4);
TASK_PP(16'h4707,4);
TASK_PP(16'h4708,4);
TASK_PP(16'h4709,4);
TASK_PP(16'h470A,4);
TASK_PP(16'h470B,4);
TASK_PP(16'h470C,4);
TASK_PP(16'h470D,4);
TASK_PP(16'h470E,4);
TASK_PP(16'h470F,4);
TASK_PP(16'h4710,4);
TASK_PP(16'h4711,4);
TASK_PP(16'h4712,4);
TASK_PP(16'h4713,4);
TASK_PP(16'h4714,4);
TASK_PP(16'h4715,4);
TASK_PP(16'h4716,4);
TASK_PP(16'h4717,4);
TASK_PP(16'h4718,4);
TASK_PP(16'h4719,4);
TASK_PP(16'h471A,4);
TASK_PP(16'h471B,4);
TASK_PP(16'h471C,4);
TASK_PP(16'h471D,4);
TASK_PP(16'h471E,4);
TASK_PP(16'h471F,4);
TASK_PP(16'h4720,4);
TASK_PP(16'h4721,4);
TASK_PP(16'h4722,4);
TASK_PP(16'h4723,4);
TASK_PP(16'h4724,4);
TASK_PP(16'h4725,4);
TASK_PP(16'h4726,4);
TASK_PP(16'h4727,4);
TASK_PP(16'h4728,4);
TASK_PP(16'h4729,4);
TASK_PP(16'h472A,4);
TASK_PP(16'h472B,4);
TASK_PP(16'h472C,4);
TASK_PP(16'h472D,4);
TASK_PP(16'h472E,4);
TASK_PP(16'h472F,4);
TASK_PP(16'h4730,4);
TASK_PP(16'h4731,4);
TASK_PP(16'h4732,4);
TASK_PP(16'h4733,4);
TASK_PP(16'h4734,4);
TASK_PP(16'h4735,4);
TASK_PP(16'h4736,4);
TASK_PP(16'h4737,4);
TASK_PP(16'h4738,4);
TASK_PP(16'h4739,4);
TASK_PP(16'h473A,4);
TASK_PP(16'h473B,4);
TASK_PP(16'h473C,4);
TASK_PP(16'h473D,4);
TASK_PP(16'h473E,4);
TASK_PP(16'h473F,4);
TASK_PP(16'h4740,4);
TASK_PP(16'h4741,4);
TASK_PP(16'h4742,4);
TASK_PP(16'h4743,4);
TASK_PP(16'h4744,4);
TASK_PP(16'h4745,4);
TASK_PP(16'h4746,4);
TASK_PP(16'h4747,4);
TASK_PP(16'h4748,4);
TASK_PP(16'h4749,4);
TASK_PP(16'h474A,4);
TASK_PP(16'h474B,4);
TASK_PP(16'h474C,4);
TASK_PP(16'h474D,4);
TASK_PP(16'h474E,4);
TASK_PP(16'h474F,4);
TASK_PP(16'h4750,4);
TASK_PP(16'h4751,4);
TASK_PP(16'h4752,4);
TASK_PP(16'h4753,4);
TASK_PP(16'h4754,4);
TASK_PP(16'h4755,4);
TASK_PP(16'h4756,4);
TASK_PP(16'h4757,4);
TASK_PP(16'h4758,4);
TASK_PP(16'h4759,4);
TASK_PP(16'h475A,4);
TASK_PP(16'h475B,4);
TASK_PP(16'h475C,4);
TASK_PP(16'h475D,4);
TASK_PP(16'h475E,4);
TASK_PP(16'h475F,4);
TASK_PP(16'h4760,4);
TASK_PP(16'h4761,4);
TASK_PP(16'h4762,4);
TASK_PP(16'h4763,4);
TASK_PP(16'h4764,4);
TASK_PP(16'h4765,4);
TASK_PP(16'h4766,4);
TASK_PP(16'h4767,4);
TASK_PP(16'h4768,4);
TASK_PP(16'h4769,4);
TASK_PP(16'h476A,4);
TASK_PP(16'h476B,4);
TASK_PP(16'h476C,4);
TASK_PP(16'h476D,4);
TASK_PP(16'h476E,4);
TASK_PP(16'h476F,4);
TASK_PP(16'h4770,4);
TASK_PP(16'h4771,4);
TASK_PP(16'h4772,4);
TASK_PP(16'h4773,4);
TASK_PP(16'h4774,4);
TASK_PP(16'h4775,4);
TASK_PP(16'h4776,4);
TASK_PP(16'h4777,4);
TASK_PP(16'h4778,4);
TASK_PP(16'h4779,4);
TASK_PP(16'h477A,4);
TASK_PP(16'h477B,4);
TASK_PP(16'h477C,4);
TASK_PP(16'h477D,4);
TASK_PP(16'h477E,4);
TASK_PP(16'h477F,4);
TASK_PP(16'h4780,4);
TASK_PP(16'h4781,4);
TASK_PP(16'h4782,4);
TASK_PP(16'h4783,4);
TASK_PP(16'h4784,4);
TASK_PP(16'h4785,4);
TASK_PP(16'h4786,4);
TASK_PP(16'h4787,4);
TASK_PP(16'h4788,4);
TASK_PP(16'h4789,4);
TASK_PP(16'h478A,4);
TASK_PP(16'h478B,4);
TASK_PP(16'h478C,4);
TASK_PP(16'h478D,4);
TASK_PP(16'h478E,4);
TASK_PP(16'h478F,4);
TASK_PP(16'h4790,4);
TASK_PP(16'h4791,4);
TASK_PP(16'h4792,4);
TASK_PP(16'h4793,4);
TASK_PP(16'h4794,4);
TASK_PP(16'h4795,4);
TASK_PP(16'h4796,4);
TASK_PP(16'h4797,4);
TASK_PP(16'h4798,4);
TASK_PP(16'h4799,4);
TASK_PP(16'h479A,4);
TASK_PP(16'h479B,4);
TASK_PP(16'h479C,4);
TASK_PP(16'h479D,4);
TASK_PP(16'h479E,4);
TASK_PP(16'h479F,4);
TASK_PP(16'h47A0,4);
TASK_PP(16'h47A1,4);
TASK_PP(16'h47A2,4);
TASK_PP(16'h47A3,4);
TASK_PP(16'h47A4,4);
TASK_PP(16'h47A5,4);
TASK_PP(16'h47A6,4);
TASK_PP(16'h47A7,4);
TASK_PP(16'h47A8,4);
TASK_PP(16'h47A9,4);
TASK_PP(16'h47AA,4);
TASK_PP(16'h47AB,4);
TASK_PP(16'h47AC,4);
TASK_PP(16'h47AD,4);
TASK_PP(16'h47AE,4);
TASK_PP(16'h47AF,4);
TASK_PP(16'h47B0,4);
TASK_PP(16'h47B1,4);
TASK_PP(16'h47B2,4);
TASK_PP(16'h47B3,4);
TASK_PP(16'h47B4,4);
TASK_PP(16'h47B5,4);
TASK_PP(16'h47B6,4);
TASK_PP(16'h47B7,4);
TASK_PP(16'h47B8,4);
TASK_PP(16'h47B9,4);
TASK_PP(16'h47BA,4);
TASK_PP(16'h47BB,4);
TASK_PP(16'h47BC,4);
TASK_PP(16'h47BD,4);
TASK_PP(16'h47BE,4);
TASK_PP(16'h47BF,4);
TASK_PP(16'h47C0,4);
TASK_PP(16'h47C1,4);
TASK_PP(16'h47C2,4);
TASK_PP(16'h47C3,4);
TASK_PP(16'h47C4,4);
TASK_PP(16'h47C5,4);
TASK_PP(16'h47C6,4);
TASK_PP(16'h47C7,4);
TASK_PP(16'h47C8,4);
TASK_PP(16'h47C9,4);
TASK_PP(16'h47CA,4);
TASK_PP(16'h47CB,4);
TASK_PP(16'h47CC,4);
TASK_PP(16'h47CD,4);
TASK_PP(16'h47CE,4);
TASK_PP(16'h47CF,4);
TASK_PP(16'h47D0,4);
TASK_PP(16'h47D1,4);
TASK_PP(16'h47D2,4);
TASK_PP(16'h47D3,4);
TASK_PP(16'h47D4,4);
TASK_PP(16'h47D5,4);
TASK_PP(16'h47D6,4);
TASK_PP(16'h47D7,4);
TASK_PP(16'h47D8,4);
TASK_PP(16'h47D9,4);
TASK_PP(16'h47DA,4);
TASK_PP(16'h47DB,4);
TASK_PP(16'h47DC,4);
TASK_PP(16'h47DD,4);
TASK_PP(16'h47DE,4);
TASK_PP(16'h47DF,4);
TASK_PP(16'h47E0,4);
TASK_PP(16'h47E1,4);
TASK_PP(16'h47E2,4);
TASK_PP(16'h47E3,4);
TASK_PP(16'h47E4,4);
TASK_PP(16'h47E5,4);
TASK_PP(16'h47E6,4);
TASK_PP(16'h47E7,4);
TASK_PP(16'h47E8,4);
TASK_PP(16'h47E9,4);
TASK_PP(16'h47EA,4);
TASK_PP(16'h47EB,4);
TASK_PP(16'h47EC,4);
TASK_PP(16'h47ED,4);
TASK_PP(16'h47EE,4);
TASK_PP(16'h47EF,4);
TASK_PP(16'h47F0,4);
TASK_PP(16'h47F1,4);
TASK_PP(16'h47F2,4);
TASK_PP(16'h47F3,4);
TASK_PP(16'h47F4,4);
TASK_PP(16'h47F5,4);
TASK_PP(16'h47F6,4);
TASK_PP(16'h47F7,4);
TASK_PP(16'h47F8,4);
TASK_PP(16'h47F9,4);
TASK_PP(16'h47FA,4);
TASK_PP(16'h47FB,4);
TASK_PP(16'h47FC,4);
TASK_PP(16'h47FD,4);
TASK_PP(16'h47FE,4);
TASK_PP(16'h47FF,4);
TASK_PP(16'h4800,4);
TASK_PP(16'h4801,4);
TASK_PP(16'h4802,4);
TASK_PP(16'h4803,4);
TASK_PP(16'h4804,4);
TASK_PP(16'h4805,4);
TASK_PP(16'h4806,4);
TASK_PP(16'h4807,4);
TASK_PP(16'h4808,4);
TASK_PP(16'h4809,4);
TASK_PP(16'h480A,4);
TASK_PP(16'h480B,4);
TASK_PP(16'h480C,4);
TASK_PP(16'h480D,4);
TASK_PP(16'h480E,4);
TASK_PP(16'h480F,4);
TASK_PP(16'h4810,4);
TASK_PP(16'h4811,4);
TASK_PP(16'h4812,4);
TASK_PP(16'h4813,4);
TASK_PP(16'h4814,4);
TASK_PP(16'h4815,4);
TASK_PP(16'h4816,4);
TASK_PP(16'h4817,4);
TASK_PP(16'h4818,4);
TASK_PP(16'h4819,4);
TASK_PP(16'h481A,4);
TASK_PP(16'h481B,4);
TASK_PP(16'h481C,4);
TASK_PP(16'h481D,4);
TASK_PP(16'h481E,4);
TASK_PP(16'h481F,4);
TASK_PP(16'h4820,4);
TASK_PP(16'h4821,4);
TASK_PP(16'h4822,4);
TASK_PP(16'h4823,4);
TASK_PP(16'h4824,4);
TASK_PP(16'h4825,4);
TASK_PP(16'h4826,4);
TASK_PP(16'h4827,4);
TASK_PP(16'h4828,4);
TASK_PP(16'h4829,4);
TASK_PP(16'h482A,4);
TASK_PP(16'h482B,4);
TASK_PP(16'h482C,4);
TASK_PP(16'h482D,4);
TASK_PP(16'h482E,4);
TASK_PP(16'h482F,4);
TASK_PP(16'h4830,4);
TASK_PP(16'h4831,4);
TASK_PP(16'h4832,4);
TASK_PP(16'h4833,4);
TASK_PP(16'h4834,4);
TASK_PP(16'h4835,4);
TASK_PP(16'h4836,4);
TASK_PP(16'h4837,4);
TASK_PP(16'h4838,4);
TASK_PP(16'h4839,4);
TASK_PP(16'h483A,4);
TASK_PP(16'h483B,4);
TASK_PP(16'h483C,4);
TASK_PP(16'h483D,4);
TASK_PP(16'h483E,4);
TASK_PP(16'h483F,4);
TASK_PP(16'h4840,4);
TASK_PP(16'h4841,4);
TASK_PP(16'h4842,4);
TASK_PP(16'h4843,4);
TASK_PP(16'h4844,4);
TASK_PP(16'h4845,4);
TASK_PP(16'h4846,4);
TASK_PP(16'h4847,4);
TASK_PP(16'h4848,4);
TASK_PP(16'h4849,4);
TASK_PP(16'h484A,4);
TASK_PP(16'h484B,4);
TASK_PP(16'h484C,4);
TASK_PP(16'h484D,4);
TASK_PP(16'h484E,4);
TASK_PP(16'h484F,4);
TASK_PP(16'h4850,4);
TASK_PP(16'h4851,4);
TASK_PP(16'h4852,4);
TASK_PP(16'h4853,4);
TASK_PP(16'h4854,4);
TASK_PP(16'h4855,4);
TASK_PP(16'h4856,4);
TASK_PP(16'h4857,4);
TASK_PP(16'h4858,4);
TASK_PP(16'h4859,4);
TASK_PP(16'h485A,4);
TASK_PP(16'h485B,4);
TASK_PP(16'h485C,4);
TASK_PP(16'h485D,4);
TASK_PP(16'h485E,4);
TASK_PP(16'h485F,4);
TASK_PP(16'h4860,4);
TASK_PP(16'h4861,4);
TASK_PP(16'h4862,4);
TASK_PP(16'h4863,4);
TASK_PP(16'h4864,4);
TASK_PP(16'h4865,4);
TASK_PP(16'h4866,4);
TASK_PP(16'h4867,4);
TASK_PP(16'h4868,4);
TASK_PP(16'h4869,4);
TASK_PP(16'h486A,4);
TASK_PP(16'h486B,4);
TASK_PP(16'h486C,4);
TASK_PP(16'h486D,4);
TASK_PP(16'h486E,4);
TASK_PP(16'h486F,4);
TASK_PP(16'h4870,4);
TASK_PP(16'h4871,4);
TASK_PP(16'h4872,4);
TASK_PP(16'h4873,4);
TASK_PP(16'h4874,4);
TASK_PP(16'h4875,4);
TASK_PP(16'h4876,4);
TASK_PP(16'h4877,4);
TASK_PP(16'h4878,4);
TASK_PP(16'h4879,4);
TASK_PP(16'h487A,4);
TASK_PP(16'h487B,4);
TASK_PP(16'h487C,4);
TASK_PP(16'h487D,4);
TASK_PP(16'h487E,4);
TASK_PP(16'h487F,4);
TASK_PP(16'h4880,4);
TASK_PP(16'h4881,4);
TASK_PP(16'h4882,4);
TASK_PP(16'h4883,4);
TASK_PP(16'h4884,4);
TASK_PP(16'h4885,4);
TASK_PP(16'h4886,4);
TASK_PP(16'h4887,4);
TASK_PP(16'h4888,4);
TASK_PP(16'h4889,4);
TASK_PP(16'h488A,4);
TASK_PP(16'h488B,4);
TASK_PP(16'h488C,4);
TASK_PP(16'h488D,4);
TASK_PP(16'h488E,4);
TASK_PP(16'h488F,4);
TASK_PP(16'h4890,4);
TASK_PP(16'h4891,4);
TASK_PP(16'h4892,4);
TASK_PP(16'h4893,4);
TASK_PP(16'h4894,4);
TASK_PP(16'h4895,4);
TASK_PP(16'h4896,4);
TASK_PP(16'h4897,4);
TASK_PP(16'h4898,4);
TASK_PP(16'h4899,4);
TASK_PP(16'h489A,4);
TASK_PP(16'h489B,4);
TASK_PP(16'h489C,4);
TASK_PP(16'h489D,4);
TASK_PP(16'h489E,4);
TASK_PP(16'h489F,4);
TASK_PP(16'h48A0,4);
TASK_PP(16'h48A1,4);
TASK_PP(16'h48A2,4);
TASK_PP(16'h48A3,4);
TASK_PP(16'h48A4,4);
TASK_PP(16'h48A5,4);
TASK_PP(16'h48A6,4);
TASK_PP(16'h48A7,4);
TASK_PP(16'h48A8,4);
TASK_PP(16'h48A9,4);
TASK_PP(16'h48AA,4);
TASK_PP(16'h48AB,4);
TASK_PP(16'h48AC,4);
TASK_PP(16'h48AD,4);
TASK_PP(16'h48AE,4);
TASK_PP(16'h48AF,4);
TASK_PP(16'h48B0,4);
TASK_PP(16'h48B1,4);
TASK_PP(16'h48B2,4);
TASK_PP(16'h48B3,4);
TASK_PP(16'h48B4,4);
TASK_PP(16'h48B5,4);
TASK_PP(16'h48B6,4);
TASK_PP(16'h48B7,4);
TASK_PP(16'h48B8,4);
TASK_PP(16'h48B9,4);
TASK_PP(16'h48BA,4);
TASK_PP(16'h48BB,4);
TASK_PP(16'h48BC,4);
TASK_PP(16'h48BD,4);
TASK_PP(16'h48BE,4);
TASK_PP(16'h48BF,4);
TASK_PP(16'h48C0,4);
TASK_PP(16'h48C1,4);
TASK_PP(16'h48C2,4);
TASK_PP(16'h48C3,4);
TASK_PP(16'h48C4,4);
TASK_PP(16'h48C5,4);
TASK_PP(16'h48C6,4);
TASK_PP(16'h48C7,4);
TASK_PP(16'h48C8,4);
TASK_PP(16'h48C9,4);
TASK_PP(16'h48CA,4);
TASK_PP(16'h48CB,4);
TASK_PP(16'h48CC,4);
TASK_PP(16'h48CD,4);
TASK_PP(16'h48CE,4);
TASK_PP(16'h48CF,4);
TASK_PP(16'h48D0,4);
TASK_PP(16'h48D1,4);
TASK_PP(16'h48D2,4);
TASK_PP(16'h48D3,4);
TASK_PP(16'h48D4,4);
TASK_PP(16'h48D5,4);
TASK_PP(16'h48D6,4);
TASK_PP(16'h48D7,4);
TASK_PP(16'h48D8,4);
TASK_PP(16'h48D9,4);
TASK_PP(16'h48DA,4);
TASK_PP(16'h48DB,4);
TASK_PP(16'h48DC,4);
TASK_PP(16'h48DD,4);
TASK_PP(16'h48DE,4);
TASK_PP(16'h48DF,4);
TASK_PP(16'h48E0,4);
TASK_PP(16'h48E1,4);
TASK_PP(16'h48E2,4);
TASK_PP(16'h48E3,4);
TASK_PP(16'h48E4,4);
TASK_PP(16'h48E5,4);
TASK_PP(16'h48E6,4);
TASK_PP(16'h48E7,4);
TASK_PP(16'h48E8,4);
TASK_PP(16'h48E9,4);
TASK_PP(16'h48EA,4);
TASK_PP(16'h48EB,4);
TASK_PP(16'h48EC,4);
TASK_PP(16'h48ED,4);
TASK_PP(16'h48EE,4);
TASK_PP(16'h48EF,4);
TASK_PP(16'h48F0,4);
TASK_PP(16'h48F1,4);
TASK_PP(16'h48F2,4);
TASK_PP(16'h48F3,4);
TASK_PP(16'h48F4,4);
TASK_PP(16'h48F5,4);
TASK_PP(16'h48F6,4);
TASK_PP(16'h48F7,4);
TASK_PP(16'h48F8,4);
TASK_PP(16'h48F9,4);
TASK_PP(16'h48FA,4);
TASK_PP(16'h48FB,4);
TASK_PP(16'h48FC,4);
TASK_PP(16'h48FD,4);
TASK_PP(16'h48FE,4);
TASK_PP(16'h48FF,4);
TASK_PP(16'h4900,4);
TASK_PP(16'h4901,4);
TASK_PP(16'h4902,4);
TASK_PP(16'h4903,4);
TASK_PP(16'h4904,4);
TASK_PP(16'h4905,4);
TASK_PP(16'h4906,4);
TASK_PP(16'h4907,4);
TASK_PP(16'h4908,4);
TASK_PP(16'h4909,4);
TASK_PP(16'h490A,4);
TASK_PP(16'h490B,4);
TASK_PP(16'h490C,4);
TASK_PP(16'h490D,4);
TASK_PP(16'h490E,4);
TASK_PP(16'h490F,4);
TASK_PP(16'h4910,4);
TASK_PP(16'h4911,4);
TASK_PP(16'h4912,4);
TASK_PP(16'h4913,4);
TASK_PP(16'h4914,4);
TASK_PP(16'h4915,4);
TASK_PP(16'h4916,4);
TASK_PP(16'h4917,4);
TASK_PP(16'h4918,4);
TASK_PP(16'h4919,4);
TASK_PP(16'h491A,4);
TASK_PP(16'h491B,4);
TASK_PP(16'h491C,4);
TASK_PP(16'h491D,4);
TASK_PP(16'h491E,4);
TASK_PP(16'h491F,4);
TASK_PP(16'h4920,4);
TASK_PP(16'h4921,4);
TASK_PP(16'h4922,4);
TASK_PP(16'h4923,4);
TASK_PP(16'h4924,4);
TASK_PP(16'h4925,4);
TASK_PP(16'h4926,4);
TASK_PP(16'h4927,4);
TASK_PP(16'h4928,4);
TASK_PP(16'h4929,4);
TASK_PP(16'h492A,4);
TASK_PP(16'h492B,4);
TASK_PP(16'h492C,4);
TASK_PP(16'h492D,4);
TASK_PP(16'h492E,4);
TASK_PP(16'h492F,4);
TASK_PP(16'h4930,4);
TASK_PP(16'h4931,4);
TASK_PP(16'h4932,4);
TASK_PP(16'h4933,4);
TASK_PP(16'h4934,4);
TASK_PP(16'h4935,4);
TASK_PP(16'h4936,4);
TASK_PP(16'h4937,4);
TASK_PP(16'h4938,4);
TASK_PP(16'h4939,4);
TASK_PP(16'h493A,4);
TASK_PP(16'h493B,4);
TASK_PP(16'h493C,4);
TASK_PP(16'h493D,4);
TASK_PP(16'h493E,4);
TASK_PP(16'h493F,4);
TASK_PP(16'h4940,4);
TASK_PP(16'h4941,4);
TASK_PP(16'h4942,4);
TASK_PP(16'h4943,4);
TASK_PP(16'h4944,4);
TASK_PP(16'h4945,4);
TASK_PP(16'h4946,4);
TASK_PP(16'h4947,4);
TASK_PP(16'h4948,4);
TASK_PP(16'h4949,4);
TASK_PP(16'h494A,4);
TASK_PP(16'h494B,4);
TASK_PP(16'h494C,4);
TASK_PP(16'h494D,4);
TASK_PP(16'h494E,4);
TASK_PP(16'h494F,4);
TASK_PP(16'h4950,4);
TASK_PP(16'h4951,4);
TASK_PP(16'h4952,4);
TASK_PP(16'h4953,4);
TASK_PP(16'h4954,4);
TASK_PP(16'h4955,4);
TASK_PP(16'h4956,4);
TASK_PP(16'h4957,4);
TASK_PP(16'h4958,4);
TASK_PP(16'h4959,4);
TASK_PP(16'h495A,4);
TASK_PP(16'h495B,4);
TASK_PP(16'h495C,4);
TASK_PP(16'h495D,4);
TASK_PP(16'h495E,4);
TASK_PP(16'h495F,4);
TASK_PP(16'h4960,4);
TASK_PP(16'h4961,4);
TASK_PP(16'h4962,4);
TASK_PP(16'h4963,4);
TASK_PP(16'h4964,4);
TASK_PP(16'h4965,4);
TASK_PP(16'h4966,4);
TASK_PP(16'h4967,4);
TASK_PP(16'h4968,4);
TASK_PP(16'h4969,4);
TASK_PP(16'h496A,4);
TASK_PP(16'h496B,4);
TASK_PP(16'h496C,4);
TASK_PP(16'h496D,4);
TASK_PP(16'h496E,4);
TASK_PP(16'h496F,4);
TASK_PP(16'h4970,4);
TASK_PP(16'h4971,4);
TASK_PP(16'h4972,4);
TASK_PP(16'h4973,4);
TASK_PP(16'h4974,4);
TASK_PP(16'h4975,4);
TASK_PP(16'h4976,4);
TASK_PP(16'h4977,4);
TASK_PP(16'h4978,4);
TASK_PP(16'h4979,4);
TASK_PP(16'h497A,4);
TASK_PP(16'h497B,4);
TASK_PP(16'h497C,4);
TASK_PP(16'h497D,4);
TASK_PP(16'h497E,4);
TASK_PP(16'h497F,4);
TASK_PP(16'h4980,4);
TASK_PP(16'h4981,4);
TASK_PP(16'h4982,4);
TASK_PP(16'h4983,4);
TASK_PP(16'h4984,4);
TASK_PP(16'h4985,4);
TASK_PP(16'h4986,4);
TASK_PP(16'h4987,4);
TASK_PP(16'h4988,4);
TASK_PP(16'h4989,4);
TASK_PP(16'h498A,4);
TASK_PP(16'h498B,4);
TASK_PP(16'h498C,4);
TASK_PP(16'h498D,4);
TASK_PP(16'h498E,4);
TASK_PP(16'h498F,4);
TASK_PP(16'h4990,4);
TASK_PP(16'h4991,4);
TASK_PP(16'h4992,4);
TASK_PP(16'h4993,4);
TASK_PP(16'h4994,4);
TASK_PP(16'h4995,4);
TASK_PP(16'h4996,4);
TASK_PP(16'h4997,4);
TASK_PP(16'h4998,4);
TASK_PP(16'h4999,4);
TASK_PP(16'h499A,4);
TASK_PP(16'h499B,4);
TASK_PP(16'h499C,4);
TASK_PP(16'h499D,4);
TASK_PP(16'h499E,4);
TASK_PP(16'h499F,4);
TASK_PP(16'h49A0,4);
TASK_PP(16'h49A1,4);
TASK_PP(16'h49A2,4);
TASK_PP(16'h49A3,4);
TASK_PP(16'h49A4,4);
TASK_PP(16'h49A5,4);
TASK_PP(16'h49A6,4);
TASK_PP(16'h49A7,4);
TASK_PP(16'h49A8,4);
TASK_PP(16'h49A9,4);
TASK_PP(16'h49AA,4);
TASK_PP(16'h49AB,4);
TASK_PP(16'h49AC,4);
TASK_PP(16'h49AD,4);
TASK_PP(16'h49AE,4);
TASK_PP(16'h49AF,4);
TASK_PP(16'h49B0,4);
TASK_PP(16'h49B1,4);
TASK_PP(16'h49B2,4);
TASK_PP(16'h49B3,4);
TASK_PP(16'h49B4,4);
TASK_PP(16'h49B5,4);
TASK_PP(16'h49B6,4);
TASK_PP(16'h49B7,4);
TASK_PP(16'h49B8,4);
TASK_PP(16'h49B9,4);
TASK_PP(16'h49BA,4);
TASK_PP(16'h49BB,4);
TASK_PP(16'h49BC,4);
TASK_PP(16'h49BD,4);
TASK_PP(16'h49BE,4);
TASK_PP(16'h49BF,4);
TASK_PP(16'h49C0,4);
TASK_PP(16'h49C1,4);
TASK_PP(16'h49C2,4);
TASK_PP(16'h49C3,4);
TASK_PP(16'h49C4,4);
TASK_PP(16'h49C5,4);
TASK_PP(16'h49C6,4);
TASK_PP(16'h49C7,4);
TASK_PP(16'h49C8,4);
TASK_PP(16'h49C9,4);
TASK_PP(16'h49CA,4);
TASK_PP(16'h49CB,4);
TASK_PP(16'h49CC,4);
TASK_PP(16'h49CD,4);
TASK_PP(16'h49CE,4);
TASK_PP(16'h49CF,4);
TASK_PP(16'h49D0,4);
TASK_PP(16'h49D1,4);
TASK_PP(16'h49D2,4);
TASK_PP(16'h49D3,4);
TASK_PP(16'h49D4,4);
TASK_PP(16'h49D5,4);
TASK_PP(16'h49D6,4);
TASK_PP(16'h49D7,4);
TASK_PP(16'h49D8,4);
TASK_PP(16'h49D9,4);
TASK_PP(16'h49DA,4);
TASK_PP(16'h49DB,4);
TASK_PP(16'h49DC,4);
TASK_PP(16'h49DD,4);
TASK_PP(16'h49DE,4);
TASK_PP(16'h49DF,4);
TASK_PP(16'h49E0,4);
TASK_PP(16'h49E1,4);
TASK_PP(16'h49E2,4);
TASK_PP(16'h49E3,4);
TASK_PP(16'h49E4,4);
TASK_PP(16'h49E5,4);
TASK_PP(16'h49E6,4);
TASK_PP(16'h49E7,4);
TASK_PP(16'h49E8,4);
TASK_PP(16'h49E9,4);
TASK_PP(16'h49EA,4);
TASK_PP(16'h49EB,4);
TASK_PP(16'h49EC,4);
TASK_PP(16'h49ED,4);
TASK_PP(16'h49EE,4);
TASK_PP(16'h49EF,4);
TASK_PP(16'h49F0,4);
TASK_PP(16'h49F1,4);
TASK_PP(16'h49F2,4);
TASK_PP(16'h49F3,4);
TASK_PP(16'h49F4,4);
TASK_PP(16'h49F5,4);
TASK_PP(16'h49F6,4);
TASK_PP(16'h49F7,4);
TASK_PP(16'h49F8,4);
TASK_PP(16'h49F9,4);
TASK_PP(16'h49FA,4);
TASK_PP(16'h49FB,4);
TASK_PP(16'h49FC,4);
TASK_PP(16'h49FD,4);
TASK_PP(16'h49FE,4);
TASK_PP(16'h49FF,4);
TASK_PP(16'h4A00,4);
TASK_PP(16'h4A01,4);
TASK_PP(16'h4A02,4);
TASK_PP(16'h4A03,4);
TASK_PP(16'h4A04,4);
TASK_PP(16'h4A05,4);
TASK_PP(16'h4A06,4);
TASK_PP(16'h4A07,4);
TASK_PP(16'h4A08,4);
TASK_PP(16'h4A09,4);
TASK_PP(16'h4A0A,4);
TASK_PP(16'h4A0B,4);
TASK_PP(16'h4A0C,4);
TASK_PP(16'h4A0D,4);
TASK_PP(16'h4A0E,4);
TASK_PP(16'h4A0F,4);
TASK_PP(16'h4A10,4);
TASK_PP(16'h4A11,4);
TASK_PP(16'h4A12,4);
TASK_PP(16'h4A13,4);
TASK_PP(16'h4A14,4);
TASK_PP(16'h4A15,4);
TASK_PP(16'h4A16,4);
TASK_PP(16'h4A17,4);
TASK_PP(16'h4A18,4);
TASK_PP(16'h4A19,4);
TASK_PP(16'h4A1A,4);
TASK_PP(16'h4A1B,4);
TASK_PP(16'h4A1C,4);
TASK_PP(16'h4A1D,4);
TASK_PP(16'h4A1E,4);
TASK_PP(16'h4A1F,4);
TASK_PP(16'h4A20,4);
TASK_PP(16'h4A21,4);
TASK_PP(16'h4A22,4);
TASK_PP(16'h4A23,4);
TASK_PP(16'h4A24,4);
TASK_PP(16'h4A25,4);
TASK_PP(16'h4A26,4);
TASK_PP(16'h4A27,4);
TASK_PP(16'h4A28,4);
TASK_PP(16'h4A29,4);
TASK_PP(16'h4A2A,4);
TASK_PP(16'h4A2B,4);
TASK_PP(16'h4A2C,4);
TASK_PP(16'h4A2D,4);
TASK_PP(16'h4A2E,4);
TASK_PP(16'h4A2F,4);
TASK_PP(16'h4A30,4);
TASK_PP(16'h4A31,4);
TASK_PP(16'h4A32,4);
TASK_PP(16'h4A33,4);
TASK_PP(16'h4A34,4);
TASK_PP(16'h4A35,4);
TASK_PP(16'h4A36,4);
TASK_PP(16'h4A37,4);
TASK_PP(16'h4A38,4);
TASK_PP(16'h4A39,4);
TASK_PP(16'h4A3A,4);
TASK_PP(16'h4A3B,4);
TASK_PP(16'h4A3C,4);
TASK_PP(16'h4A3D,4);
TASK_PP(16'h4A3E,4);
TASK_PP(16'h4A3F,4);
TASK_PP(16'h4A40,4);
TASK_PP(16'h4A41,4);
TASK_PP(16'h4A42,4);
TASK_PP(16'h4A43,4);
TASK_PP(16'h4A44,4);
TASK_PP(16'h4A45,4);
TASK_PP(16'h4A46,4);
TASK_PP(16'h4A47,4);
TASK_PP(16'h4A48,4);
TASK_PP(16'h4A49,4);
TASK_PP(16'h4A4A,4);
TASK_PP(16'h4A4B,4);
TASK_PP(16'h4A4C,4);
TASK_PP(16'h4A4D,4);
TASK_PP(16'h4A4E,4);
TASK_PP(16'h4A4F,4);
TASK_PP(16'h4A50,4);
TASK_PP(16'h4A51,4);
TASK_PP(16'h4A52,4);
TASK_PP(16'h4A53,4);
TASK_PP(16'h4A54,4);
TASK_PP(16'h4A55,4);
TASK_PP(16'h4A56,4);
TASK_PP(16'h4A57,4);
TASK_PP(16'h4A58,4);
TASK_PP(16'h4A59,4);
TASK_PP(16'h4A5A,4);
TASK_PP(16'h4A5B,4);
TASK_PP(16'h4A5C,4);
TASK_PP(16'h4A5D,4);
TASK_PP(16'h4A5E,4);
TASK_PP(16'h4A5F,4);
TASK_PP(16'h4A60,4);
TASK_PP(16'h4A61,4);
TASK_PP(16'h4A62,4);
TASK_PP(16'h4A63,4);
TASK_PP(16'h4A64,4);
TASK_PP(16'h4A65,4);
TASK_PP(16'h4A66,4);
TASK_PP(16'h4A67,4);
TASK_PP(16'h4A68,4);
TASK_PP(16'h4A69,4);
TASK_PP(16'h4A6A,4);
TASK_PP(16'h4A6B,4);
TASK_PP(16'h4A6C,4);
TASK_PP(16'h4A6D,4);
TASK_PP(16'h4A6E,4);
TASK_PP(16'h4A6F,4);
TASK_PP(16'h4A70,4);
TASK_PP(16'h4A71,4);
TASK_PP(16'h4A72,4);
TASK_PP(16'h4A73,4);
TASK_PP(16'h4A74,4);
TASK_PP(16'h4A75,4);
TASK_PP(16'h4A76,4);
TASK_PP(16'h4A77,4);
TASK_PP(16'h4A78,4);
TASK_PP(16'h4A79,4);
TASK_PP(16'h4A7A,4);
TASK_PP(16'h4A7B,4);
TASK_PP(16'h4A7C,4);
TASK_PP(16'h4A7D,4);
TASK_PP(16'h4A7E,4);
TASK_PP(16'h4A7F,4);
TASK_PP(16'h4A80,4);
TASK_PP(16'h4A81,4);
TASK_PP(16'h4A82,4);
TASK_PP(16'h4A83,4);
TASK_PP(16'h4A84,4);
TASK_PP(16'h4A85,4);
TASK_PP(16'h4A86,4);
TASK_PP(16'h4A87,4);
TASK_PP(16'h4A88,4);
TASK_PP(16'h4A89,4);
TASK_PP(16'h4A8A,4);
TASK_PP(16'h4A8B,4);
TASK_PP(16'h4A8C,4);
TASK_PP(16'h4A8D,4);
TASK_PP(16'h4A8E,4);
TASK_PP(16'h4A8F,4);
TASK_PP(16'h4A90,4);
TASK_PP(16'h4A91,4);
TASK_PP(16'h4A92,4);
TASK_PP(16'h4A93,4);
TASK_PP(16'h4A94,4);
TASK_PP(16'h4A95,4);
TASK_PP(16'h4A96,4);
TASK_PP(16'h4A97,4);
TASK_PP(16'h4A98,4);
TASK_PP(16'h4A99,4);
TASK_PP(16'h4A9A,4);
TASK_PP(16'h4A9B,4);
TASK_PP(16'h4A9C,4);
TASK_PP(16'h4A9D,4);
TASK_PP(16'h4A9E,4);
TASK_PP(16'h4A9F,4);
TASK_PP(16'h4AA0,4);
TASK_PP(16'h4AA1,4);
TASK_PP(16'h4AA2,4);
TASK_PP(16'h4AA3,4);
TASK_PP(16'h4AA4,4);
TASK_PP(16'h4AA5,4);
TASK_PP(16'h4AA6,4);
TASK_PP(16'h4AA7,4);
TASK_PP(16'h4AA8,4);
TASK_PP(16'h4AA9,4);
TASK_PP(16'h4AAA,4);
TASK_PP(16'h4AAB,4);
TASK_PP(16'h4AAC,4);
TASK_PP(16'h4AAD,4);
TASK_PP(16'h4AAE,4);
TASK_PP(16'h4AAF,4);
TASK_PP(16'h4AB0,4);
TASK_PP(16'h4AB1,4);
TASK_PP(16'h4AB2,4);
TASK_PP(16'h4AB3,4);
TASK_PP(16'h4AB4,4);
TASK_PP(16'h4AB5,4);
TASK_PP(16'h4AB6,4);
TASK_PP(16'h4AB7,4);
TASK_PP(16'h4AB8,4);
TASK_PP(16'h4AB9,4);
TASK_PP(16'h4ABA,4);
TASK_PP(16'h4ABB,4);
TASK_PP(16'h4ABC,4);
TASK_PP(16'h4ABD,4);
TASK_PP(16'h4ABE,4);
TASK_PP(16'h4ABF,4);
TASK_PP(16'h4AC0,4);
TASK_PP(16'h4AC1,4);
TASK_PP(16'h4AC2,4);
TASK_PP(16'h4AC3,4);
TASK_PP(16'h4AC4,4);
TASK_PP(16'h4AC5,4);
TASK_PP(16'h4AC6,4);
TASK_PP(16'h4AC7,4);
TASK_PP(16'h4AC8,4);
TASK_PP(16'h4AC9,4);
TASK_PP(16'h4ACA,4);
TASK_PP(16'h4ACB,4);
TASK_PP(16'h4ACC,4);
TASK_PP(16'h4ACD,4);
TASK_PP(16'h4ACE,4);
TASK_PP(16'h4ACF,4);
TASK_PP(16'h4AD0,4);
TASK_PP(16'h4AD1,4);
TASK_PP(16'h4AD2,4);
TASK_PP(16'h4AD3,4);
TASK_PP(16'h4AD4,4);
TASK_PP(16'h4AD5,4);
TASK_PP(16'h4AD6,4);
TASK_PP(16'h4AD7,4);
TASK_PP(16'h4AD8,4);
TASK_PP(16'h4AD9,4);
TASK_PP(16'h4ADA,4);
TASK_PP(16'h4ADB,4);
TASK_PP(16'h4ADC,4);
TASK_PP(16'h4ADD,4);
TASK_PP(16'h4ADE,4);
TASK_PP(16'h4ADF,4);
TASK_PP(16'h4AE0,4);
TASK_PP(16'h4AE1,4);
TASK_PP(16'h4AE2,4);
TASK_PP(16'h4AE3,4);
TASK_PP(16'h4AE4,4);
TASK_PP(16'h4AE5,4);
TASK_PP(16'h4AE6,4);
TASK_PP(16'h4AE7,4);
TASK_PP(16'h4AE8,4);
TASK_PP(16'h4AE9,4);
TASK_PP(16'h4AEA,4);
TASK_PP(16'h4AEB,4);
TASK_PP(16'h4AEC,4);
TASK_PP(16'h4AED,4);
TASK_PP(16'h4AEE,4);
TASK_PP(16'h4AEF,4);
TASK_PP(16'h4AF0,4);
TASK_PP(16'h4AF1,4);
TASK_PP(16'h4AF2,4);
TASK_PP(16'h4AF3,4);
TASK_PP(16'h4AF4,4);
TASK_PP(16'h4AF5,4);
TASK_PP(16'h4AF6,4);
TASK_PP(16'h4AF7,4);
TASK_PP(16'h4AF8,4);
TASK_PP(16'h4AF9,4);
TASK_PP(16'h4AFA,4);
TASK_PP(16'h4AFB,4);
TASK_PP(16'h4AFC,4);
TASK_PP(16'h4AFD,4);
TASK_PP(16'h4AFE,4);
TASK_PP(16'h4AFF,4);
TASK_PP(16'h4B00,4);
TASK_PP(16'h4B01,4);
TASK_PP(16'h4B02,4);
TASK_PP(16'h4B03,4);
TASK_PP(16'h4B04,4);
TASK_PP(16'h4B05,4);
TASK_PP(16'h4B06,4);
TASK_PP(16'h4B07,4);
TASK_PP(16'h4B08,4);
TASK_PP(16'h4B09,4);
TASK_PP(16'h4B0A,4);
TASK_PP(16'h4B0B,4);
TASK_PP(16'h4B0C,4);
TASK_PP(16'h4B0D,4);
TASK_PP(16'h4B0E,4);
TASK_PP(16'h4B0F,4);
TASK_PP(16'h4B10,4);
TASK_PP(16'h4B11,4);
TASK_PP(16'h4B12,4);
TASK_PP(16'h4B13,4);
TASK_PP(16'h4B14,4);
TASK_PP(16'h4B15,4);
TASK_PP(16'h4B16,4);
TASK_PP(16'h4B17,4);
TASK_PP(16'h4B18,4);
TASK_PP(16'h4B19,4);
TASK_PP(16'h4B1A,4);
TASK_PP(16'h4B1B,4);
TASK_PP(16'h4B1C,4);
TASK_PP(16'h4B1D,4);
TASK_PP(16'h4B1E,4);
TASK_PP(16'h4B1F,4);
TASK_PP(16'h4B20,4);
TASK_PP(16'h4B21,4);
TASK_PP(16'h4B22,4);
TASK_PP(16'h4B23,4);
TASK_PP(16'h4B24,4);
TASK_PP(16'h4B25,4);
TASK_PP(16'h4B26,4);
TASK_PP(16'h4B27,4);
TASK_PP(16'h4B28,4);
TASK_PP(16'h4B29,4);
TASK_PP(16'h4B2A,4);
TASK_PP(16'h4B2B,4);
TASK_PP(16'h4B2C,4);
TASK_PP(16'h4B2D,4);
TASK_PP(16'h4B2E,4);
TASK_PP(16'h4B2F,4);
TASK_PP(16'h4B30,4);
TASK_PP(16'h4B31,4);
TASK_PP(16'h4B32,4);
TASK_PP(16'h4B33,4);
TASK_PP(16'h4B34,4);
TASK_PP(16'h4B35,4);
TASK_PP(16'h4B36,4);
TASK_PP(16'h4B37,4);
TASK_PP(16'h4B38,4);
TASK_PP(16'h4B39,4);
TASK_PP(16'h4B3A,4);
TASK_PP(16'h4B3B,4);
TASK_PP(16'h4B3C,4);
TASK_PP(16'h4B3D,4);
TASK_PP(16'h4B3E,4);
TASK_PP(16'h4B3F,4);
TASK_PP(16'h4B40,4);
TASK_PP(16'h4B41,4);
TASK_PP(16'h4B42,4);
TASK_PP(16'h4B43,4);
TASK_PP(16'h4B44,4);
TASK_PP(16'h4B45,4);
TASK_PP(16'h4B46,4);
TASK_PP(16'h4B47,4);
TASK_PP(16'h4B48,4);
TASK_PP(16'h4B49,4);
TASK_PP(16'h4B4A,4);
TASK_PP(16'h4B4B,4);
TASK_PP(16'h4B4C,4);
TASK_PP(16'h4B4D,4);
TASK_PP(16'h4B4E,4);
TASK_PP(16'h4B4F,4);
TASK_PP(16'h4B50,4);
TASK_PP(16'h4B51,4);
TASK_PP(16'h4B52,4);
TASK_PP(16'h4B53,4);
TASK_PP(16'h4B54,4);
TASK_PP(16'h4B55,4);
TASK_PP(16'h4B56,4);
TASK_PP(16'h4B57,4);
TASK_PP(16'h4B58,4);
TASK_PP(16'h4B59,4);
TASK_PP(16'h4B5A,4);
TASK_PP(16'h4B5B,4);
TASK_PP(16'h4B5C,4);
TASK_PP(16'h4B5D,4);
TASK_PP(16'h4B5E,4);
TASK_PP(16'h4B5F,4);
TASK_PP(16'h4B60,4);
TASK_PP(16'h4B61,4);
TASK_PP(16'h4B62,4);
TASK_PP(16'h4B63,4);
TASK_PP(16'h4B64,4);
TASK_PP(16'h4B65,4);
TASK_PP(16'h4B66,4);
TASK_PP(16'h4B67,4);
TASK_PP(16'h4B68,4);
TASK_PP(16'h4B69,4);
TASK_PP(16'h4B6A,4);
TASK_PP(16'h4B6B,4);
TASK_PP(16'h4B6C,4);
TASK_PP(16'h4B6D,4);
TASK_PP(16'h4B6E,4);
TASK_PP(16'h4B6F,4);
TASK_PP(16'h4B70,4);
TASK_PP(16'h4B71,4);
TASK_PP(16'h4B72,4);
TASK_PP(16'h4B73,4);
TASK_PP(16'h4B74,4);
TASK_PP(16'h4B75,4);
TASK_PP(16'h4B76,4);
TASK_PP(16'h4B77,4);
TASK_PP(16'h4B78,4);
TASK_PP(16'h4B79,4);
TASK_PP(16'h4B7A,4);
TASK_PP(16'h4B7B,4);
TASK_PP(16'h4B7C,4);
TASK_PP(16'h4B7D,4);
TASK_PP(16'h4B7E,4);
TASK_PP(16'h4B7F,4);
TASK_PP(16'h4B80,4);
TASK_PP(16'h4B81,4);
TASK_PP(16'h4B82,4);
TASK_PP(16'h4B83,4);
TASK_PP(16'h4B84,4);
TASK_PP(16'h4B85,4);
TASK_PP(16'h4B86,4);
TASK_PP(16'h4B87,4);
TASK_PP(16'h4B88,4);
TASK_PP(16'h4B89,4);
TASK_PP(16'h4B8A,4);
TASK_PP(16'h4B8B,4);
TASK_PP(16'h4B8C,4);
TASK_PP(16'h4B8D,4);
TASK_PP(16'h4B8E,4);
TASK_PP(16'h4B8F,4);
TASK_PP(16'h4B90,4);
TASK_PP(16'h4B91,4);
TASK_PP(16'h4B92,4);
TASK_PP(16'h4B93,4);
TASK_PP(16'h4B94,4);
TASK_PP(16'h4B95,4);
TASK_PP(16'h4B96,4);
TASK_PP(16'h4B97,4);
TASK_PP(16'h4B98,4);
TASK_PP(16'h4B99,4);
TASK_PP(16'h4B9A,4);
TASK_PP(16'h4B9B,4);
TASK_PP(16'h4B9C,4);
TASK_PP(16'h4B9D,4);
TASK_PP(16'h4B9E,4);
TASK_PP(16'h4B9F,4);
TASK_PP(16'h4BA0,4);
TASK_PP(16'h4BA1,4);
TASK_PP(16'h4BA2,4);
TASK_PP(16'h4BA3,4);
TASK_PP(16'h4BA4,4);
TASK_PP(16'h4BA5,4);
TASK_PP(16'h4BA6,4);
TASK_PP(16'h4BA7,4);
TASK_PP(16'h4BA8,4);
TASK_PP(16'h4BA9,4);
TASK_PP(16'h4BAA,4);
TASK_PP(16'h4BAB,4);
TASK_PP(16'h4BAC,4);
TASK_PP(16'h4BAD,4);
TASK_PP(16'h4BAE,4);
TASK_PP(16'h4BAF,4);
TASK_PP(16'h4BB0,4);
TASK_PP(16'h4BB1,4);
TASK_PP(16'h4BB2,4);
TASK_PP(16'h4BB3,4);
TASK_PP(16'h4BB4,4);
TASK_PP(16'h4BB5,4);
TASK_PP(16'h4BB6,4);
TASK_PP(16'h4BB7,4);
TASK_PP(16'h4BB8,4);
TASK_PP(16'h4BB9,4);
TASK_PP(16'h4BBA,4);
TASK_PP(16'h4BBB,4);
TASK_PP(16'h4BBC,4);
TASK_PP(16'h4BBD,4);
TASK_PP(16'h4BBE,4);
TASK_PP(16'h4BBF,4);
TASK_PP(16'h4BC0,4);
TASK_PP(16'h4BC1,4);
TASK_PP(16'h4BC2,4);
TASK_PP(16'h4BC3,4);
TASK_PP(16'h4BC4,4);
TASK_PP(16'h4BC5,4);
TASK_PP(16'h4BC6,4);
TASK_PP(16'h4BC7,4);
TASK_PP(16'h4BC8,4);
TASK_PP(16'h4BC9,4);
TASK_PP(16'h4BCA,4);
TASK_PP(16'h4BCB,4);
TASK_PP(16'h4BCC,4);
TASK_PP(16'h4BCD,4);
TASK_PP(16'h4BCE,4);
TASK_PP(16'h4BCF,4);
TASK_PP(16'h4BD0,4);
TASK_PP(16'h4BD1,4);
TASK_PP(16'h4BD2,4);
TASK_PP(16'h4BD3,4);
TASK_PP(16'h4BD4,4);
TASK_PP(16'h4BD5,4);
TASK_PP(16'h4BD6,4);
TASK_PP(16'h4BD7,4);
TASK_PP(16'h4BD8,4);
TASK_PP(16'h4BD9,4);
TASK_PP(16'h4BDA,4);
TASK_PP(16'h4BDB,4);
TASK_PP(16'h4BDC,4);
TASK_PP(16'h4BDD,4);
TASK_PP(16'h4BDE,4);
TASK_PP(16'h4BDF,4);
TASK_PP(16'h4BE0,4);
TASK_PP(16'h4BE1,4);
TASK_PP(16'h4BE2,4);
TASK_PP(16'h4BE3,4);
TASK_PP(16'h4BE4,4);
TASK_PP(16'h4BE5,4);
TASK_PP(16'h4BE6,4);
TASK_PP(16'h4BE7,4);
TASK_PP(16'h4BE8,4);
TASK_PP(16'h4BE9,4);
TASK_PP(16'h4BEA,4);
TASK_PP(16'h4BEB,4);
TASK_PP(16'h4BEC,4);
TASK_PP(16'h4BED,4);
TASK_PP(16'h4BEE,4);
TASK_PP(16'h4BEF,4);
TASK_PP(16'h4BF0,4);
TASK_PP(16'h4BF1,4);
TASK_PP(16'h4BF2,4);
TASK_PP(16'h4BF3,4);
TASK_PP(16'h4BF4,4);
TASK_PP(16'h4BF5,4);
TASK_PP(16'h4BF6,4);
TASK_PP(16'h4BF7,4);
TASK_PP(16'h4BF8,4);
TASK_PP(16'h4BF9,4);
TASK_PP(16'h4BFA,4);
TASK_PP(16'h4BFB,4);
TASK_PP(16'h4BFC,4);
TASK_PP(16'h4BFD,4);
TASK_PP(16'h4BFE,4);
TASK_PP(16'h4BFF,4);
TASK_PP(16'h4C00,4);
TASK_PP(16'h4C01,4);
TASK_PP(16'h4C02,4);
TASK_PP(16'h4C03,4);
TASK_PP(16'h4C04,4);
TASK_PP(16'h4C05,4);
TASK_PP(16'h4C06,4);
TASK_PP(16'h4C07,4);
TASK_PP(16'h4C08,4);
TASK_PP(16'h4C09,4);
TASK_PP(16'h4C0A,4);
TASK_PP(16'h4C0B,4);
TASK_PP(16'h4C0C,4);
TASK_PP(16'h4C0D,4);
TASK_PP(16'h4C0E,4);
TASK_PP(16'h4C0F,4);
TASK_PP(16'h4C10,4);
TASK_PP(16'h4C11,4);
TASK_PP(16'h4C12,4);
TASK_PP(16'h4C13,4);
TASK_PP(16'h4C14,4);
TASK_PP(16'h4C15,4);
TASK_PP(16'h4C16,4);
TASK_PP(16'h4C17,4);
TASK_PP(16'h4C18,4);
TASK_PP(16'h4C19,4);
TASK_PP(16'h4C1A,4);
TASK_PP(16'h4C1B,4);
TASK_PP(16'h4C1C,4);
TASK_PP(16'h4C1D,4);
TASK_PP(16'h4C1E,4);
TASK_PP(16'h4C1F,4);
TASK_PP(16'h4C20,4);
TASK_PP(16'h4C21,4);
TASK_PP(16'h4C22,4);
TASK_PP(16'h4C23,4);
TASK_PP(16'h4C24,4);
TASK_PP(16'h4C25,4);
TASK_PP(16'h4C26,4);
TASK_PP(16'h4C27,4);
TASK_PP(16'h4C28,4);
TASK_PP(16'h4C29,4);
TASK_PP(16'h4C2A,4);
TASK_PP(16'h4C2B,4);
TASK_PP(16'h4C2C,4);
TASK_PP(16'h4C2D,4);
TASK_PP(16'h4C2E,4);
TASK_PP(16'h4C2F,4);
TASK_PP(16'h4C30,4);
TASK_PP(16'h4C31,4);
TASK_PP(16'h4C32,4);
TASK_PP(16'h4C33,4);
TASK_PP(16'h4C34,4);
TASK_PP(16'h4C35,4);
TASK_PP(16'h4C36,4);
TASK_PP(16'h4C37,4);
TASK_PP(16'h4C38,4);
TASK_PP(16'h4C39,4);
TASK_PP(16'h4C3A,4);
TASK_PP(16'h4C3B,4);
TASK_PP(16'h4C3C,4);
TASK_PP(16'h4C3D,4);
TASK_PP(16'h4C3E,4);
TASK_PP(16'h4C3F,4);
TASK_PP(16'h4C40,4);
TASK_PP(16'h4C41,4);
TASK_PP(16'h4C42,4);
TASK_PP(16'h4C43,4);
TASK_PP(16'h4C44,4);
TASK_PP(16'h4C45,4);
TASK_PP(16'h4C46,4);
TASK_PP(16'h4C47,4);
TASK_PP(16'h4C48,4);
TASK_PP(16'h4C49,4);
TASK_PP(16'h4C4A,4);
TASK_PP(16'h4C4B,4);
TASK_PP(16'h4C4C,4);
TASK_PP(16'h4C4D,4);
TASK_PP(16'h4C4E,4);
TASK_PP(16'h4C4F,4);
TASK_PP(16'h4C50,4);
TASK_PP(16'h4C51,4);
TASK_PP(16'h4C52,4);
TASK_PP(16'h4C53,4);
TASK_PP(16'h4C54,4);
TASK_PP(16'h4C55,4);
TASK_PP(16'h4C56,4);
TASK_PP(16'h4C57,4);
TASK_PP(16'h4C58,4);
TASK_PP(16'h4C59,4);
TASK_PP(16'h4C5A,4);
TASK_PP(16'h4C5B,4);
TASK_PP(16'h4C5C,4);
TASK_PP(16'h4C5D,4);
TASK_PP(16'h4C5E,4);
TASK_PP(16'h4C5F,4);
TASK_PP(16'h4C60,4);
TASK_PP(16'h4C61,4);
TASK_PP(16'h4C62,4);
TASK_PP(16'h4C63,4);
TASK_PP(16'h4C64,4);
TASK_PP(16'h4C65,4);
TASK_PP(16'h4C66,4);
TASK_PP(16'h4C67,4);
TASK_PP(16'h4C68,4);
TASK_PP(16'h4C69,4);
TASK_PP(16'h4C6A,4);
TASK_PP(16'h4C6B,4);
TASK_PP(16'h4C6C,4);
TASK_PP(16'h4C6D,4);
TASK_PP(16'h4C6E,4);
TASK_PP(16'h4C6F,4);
TASK_PP(16'h4C70,4);
TASK_PP(16'h4C71,4);
TASK_PP(16'h4C72,4);
TASK_PP(16'h4C73,4);
TASK_PP(16'h4C74,4);
TASK_PP(16'h4C75,4);
TASK_PP(16'h4C76,4);
TASK_PP(16'h4C77,4);
TASK_PP(16'h4C78,4);
TASK_PP(16'h4C79,4);
TASK_PP(16'h4C7A,4);
TASK_PP(16'h4C7B,4);
TASK_PP(16'h4C7C,4);
TASK_PP(16'h4C7D,4);
TASK_PP(16'h4C7E,4);
TASK_PP(16'h4C7F,4);
TASK_PP(16'h4C80,4);
TASK_PP(16'h4C81,4);
TASK_PP(16'h4C82,4);
TASK_PP(16'h4C83,4);
TASK_PP(16'h4C84,4);
TASK_PP(16'h4C85,4);
TASK_PP(16'h4C86,4);
TASK_PP(16'h4C87,4);
TASK_PP(16'h4C88,4);
TASK_PP(16'h4C89,4);
TASK_PP(16'h4C8A,4);
TASK_PP(16'h4C8B,4);
TASK_PP(16'h4C8C,4);
TASK_PP(16'h4C8D,4);
TASK_PP(16'h4C8E,4);
TASK_PP(16'h4C8F,4);
TASK_PP(16'h4C90,4);
TASK_PP(16'h4C91,4);
TASK_PP(16'h4C92,4);
TASK_PP(16'h4C93,4);
TASK_PP(16'h4C94,4);
TASK_PP(16'h4C95,4);
TASK_PP(16'h4C96,4);
TASK_PP(16'h4C97,4);
TASK_PP(16'h4C98,4);
TASK_PP(16'h4C99,4);
TASK_PP(16'h4C9A,4);
TASK_PP(16'h4C9B,4);
TASK_PP(16'h4C9C,4);
TASK_PP(16'h4C9D,4);
TASK_PP(16'h4C9E,4);
TASK_PP(16'h4C9F,4);
TASK_PP(16'h4CA0,4);
TASK_PP(16'h4CA1,4);
TASK_PP(16'h4CA2,4);
TASK_PP(16'h4CA3,4);
TASK_PP(16'h4CA4,4);
TASK_PP(16'h4CA5,4);
TASK_PP(16'h4CA6,4);
TASK_PP(16'h4CA7,4);
TASK_PP(16'h4CA8,4);
TASK_PP(16'h4CA9,4);
TASK_PP(16'h4CAA,4);
TASK_PP(16'h4CAB,4);
TASK_PP(16'h4CAC,4);
TASK_PP(16'h4CAD,4);
TASK_PP(16'h4CAE,4);
TASK_PP(16'h4CAF,4);
TASK_PP(16'h4CB0,4);
TASK_PP(16'h4CB1,4);
TASK_PP(16'h4CB2,4);
TASK_PP(16'h4CB3,4);
TASK_PP(16'h4CB4,4);
TASK_PP(16'h4CB5,4);
TASK_PP(16'h4CB6,4);
TASK_PP(16'h4CB7,4);
TASK_PP(16'h4CB8,4);
TASK_PP(16'h4CB9,4);
TASK_PP(16'h4CBA,4);
TASK_PP(16'h4CBB,4);
TASK_PP(16'h4CBC,4);
TASK_PP(16'h4CBD,4);
TASK_PP(16'h4CBE,4);
TASK_PP(16'h4CBF,4);
TASK_PP(16'h4CC0,4);
TASK_PP(16'h4CC1,4);
TASK_PP(16'h4CC2,4);
TASK_PP(16'h4CC3,4);
TASK_PP(16'h4CC4,4);
TASK_PP(16'h4CC5,4);
TASK_PP(16'h4CC6,4);
TASK_PP(16'h4CC7,4);
TASK_PP(16'h4CC8,4);
TASK_PP(16'h4CC9,4);
TASK_PP(16'h4CCA,4);
TASK_PP(16'h4CCB,4);
TASK_PP(16'h4CCC,4);
TASK_PP(16'h4CCD,4);
TASK_PP(16'h4CCE,4);
TASK_PP(16'h4CCF,4);
TASK_PP(16'h4CD0,4);
TASK_PP(16'h4CD1,4);
TASK_PP(16'h4CD2,4);
TASK_PP(16'h4CD3,4);
TASK_PP(16'h4CD4,4);
TASK_PP(16'h4CD5,4);
TASK_PP(16'h4CD6,4);
TASK_PP(16'h4CD7,4);
TASK_PP(16'h4CD8,4);
TASK_PP(16'h4CD9,4);
TASK_PP(16'h4CDA,4);
TASK_PP(16'h4CDB,4);
TASK_PP(16'h4CDC,4);
TASK_PP(16'h4CDD,4);
TASK_PP(16'h4CDE,4);
TASK_PP(16'h4CDF,4);
TASK_PP(16'h4CE0,4);
TASK_PP(16'h4CE1,4);
TASK_PP(16'h4CE2,4);
TASK_PP(16'h4CE3,4);
TASK_PP(16'h4CE4,4);
TASK_PP(16'h4CE5,4);
TASK_PP(16'h4CE6,4);
TASK_PP(16'h4CE7,4);
TASK_PP(16'h4CE8,4);
TASK_PP(16'h4CE9,4);
TASK_PP(16'h4CEA,4);
TASK_PP(16'h4CEB,4);
TASK_PP(16'h4CEC,4);
TASK_PP(16'h4CED,4);
TASK_PP(16'h4CEE,4);
TASK_PP(16'h4CEF,4);
TASK_PP(16'h4CF0,4);
TASK_PP(16'h4CF1,4);
TASK_PP(16'h4CF2,4);
TASK_PP(16'h4CF3,4);
TASK_PP(16'h4CF4,4);
TASK_PP(16'h4CF5,4);
TASK_PP(16'h4CF6,4);
TASK_PP(16'h4CF7,4);
TASK_PP(16'h4CF8,4);
TASK_PP(16'h4CF9,4);
TASK_PP(16'h4CFA,4);
TASK_PP(16'h4CFB,4);
TASK_PP(16'h4CFC,4);
TASK_PP(16'h4CFD,4);
TASK_PP(16'h4CFE,4);
TASK_PP(16'h4CFF,4);
TASK_PP(16'h4D00,4);
TASK_PP(16'h4D01,4);
TASK_PP(16'h4D02,4);
TASK_PP(16'h4D03,4);
TASK_PP(16'h4D04,4);
TASK_PP(16'h4D05,4);
TASK_PP(16'h4D06,4);
TASK_PP(16'h4D07,4);
TASK_PP(16'h4D08,4);
TASK_PP(16'h4D09,4);
TASK_PP(16'h4D0A,4);
TASK_PP(16'h4D0B,4);
TASK_PP(16'h4D0C,4);
TASK_PP(16'h4D0D,4);
TASK_PP(16'h4D0E,4);
TASK_PP(16'h4D0F,4);
TASK_PP(16'h4D10,4);
TASK_PP(16'h4D11,4);
TASK_PP(16'h4D12,4);
TASK_PP(16'h4D13,4);
TASK_PP(16'h4D14,4);
TASK_PP(16'h4D15,4);
TASK_PP(16'h4D16,4);
TASK_PP(16'h4D17,4);
TASK_PP(16'h4D18,4);
TASK_PP(16'h4D19,4);
TASK_PP(16'h4D1A,4);
TASK_PP(16'h4D1B,4);
TASK_PP(16'h4D1C,4);
TASK_PP(16'h4D1D,4);
TASK_PP(16'h4D1E,4);
TASK_PP(16'h4D1F,4);
TASK_PP(16'h4D20,4);
TASK_PP(16'h4D21,4);
TASK_PP(16'h4D22,4);
TASK_PP(16'h4D23,4);
TASK_PP(16'h4D24,4);
TASK_PP(16'h4D25,4);
TASK_PP(16'h4D26,4);
TASK_PP(16'h4D27,4);
TASK_PP(16'h4D28,4);
TASK_PP(16'h4D29,4);
TASK_PP(16'h4D2A,4);
TASK_PP(16'h4D2B,4);
TASK_PP(16'h4D2C,4);
TASK_PP(16'h4D2D,4);
TASK_PP(16'h4D2E,4);
TASK_PP(16'h4D2F,4);
TASK_PP(16'h4D30,4);
TASK_PP(16'h4D31,4);
TASK_PP(16'h4D32,4);
TASK_PP(16'h4D33,4);
TASK_PP(16'h4D34,4);
TASK_PP(16'h4D35,4);
TASK_PP(16'h4D36,4);
TASK_PP(16'h4D37,4);
TASK_PP(16'h4D38,4);
TASK_PP(16'h4D39,4);
TASK_PP(16'h4D3A,4);
TASK_PP(16'h4D3B,4);
TASK_PP(16'h4D3C,4);
TASK_PP(16'h4D3D,4);
TASK_PP(16'h4D3E,4);
TASK_PP(16'h4D3F,4);
TASK_PP(16'h4D40,4);
TASK_PP(16'h4D41,4);
TASK_PP(16'h4D42,4);
TASK_PP(16'h4D43,4);
TASK_PP(16'h4D44,4);
TASK_PP(16'h4D45,4);
TASK_PP(16'h4D46,4);
TASK_PP(16'h4D47,4);
TASK_PP(16'h4D48,4);
TASK_PP(16'h4D49,4);
TASK_PP(16'h4D4A,4);
TASK_PP(16'h4D4B,4);
TASK_PP(16'h4D4C,4);
TASK_PP(16'h4D4D,4);
TASK_PP(16'h4D4E,4);
TASK_PP(16'h4D4F,4);
TASK_PP(16'h4D50,4);
TASK_PP(16'h4D51,4);
TASK_PP(16'h4D52,4);
TASK_PP(16'h4D53,4);
TASK_PP(16'h4D54,4);
TASK_PP(16'h4D55,4);
TASK_PP(16'h4D56,4);
TASK_PP(16'h4D57,4);
TASK_PP(16'h4D58,4);
TASK_PP(16'h4D59,4);
TASK_PP(16'h4D5A,4);
TASK_PP(16'h4D5B,4);
TASK_PP(16'h4D5C,4);
TASK_PP(16'h4D5D,4);
TASK_PP(16'h4D5E,4);
TASK_PP(16'h4D5F,4);
TASK_PP(16'h4D60,4);
TASK_PP(16'h4D61,4);
TASK_PP(16'h4D62,4);
TASK_PP(16'h4D63,4);
TASK_PP(16'h4D64,4);
TASK_PP(16'h4D65,4);
TASK_PP(16'h4D66,4);
TASK_PP(16'h4D67,4);
TASK_PP(16'h4D68,4);
TASK_PP(16'h4D69,4);
TASK_PP(16'h4D6A,4);
TASK_PP(16'h4D6B,4);
TASK_PP(16'h4D6C,4);
TASK_PP(16'h4D6D,4);
TASK_PP(16'h4D6E,4);
TASK_PP(16'h4D6F,4);
TASK_PP(16'h4D70,4);
TASK_PP(16'h4D71,4);
TASK_PP(16'h4D72,4);
TASK_PP(16'h4D73,4);
TASK_PP(16'h4D74,4);
TASK_PP(16'h4D75,4);
TASK_PP(16'h4D76,4);
TASK_PP(16'h4D77,4);
TASK_PP(16'h4D78,4);
TASK_PP(16'h4D79,4);
TASK_PP(16'h4D7A,4);
TASK_PP(16'h4D7B,4);
TASK_PP(16'h4D7C,4);
TASK_PP(16'h4D7D,4);
TASK_PP(16'h4D7E,4);
TASK_PP(16'h4D7F,4);
TASK_PP(16'h4D80,4);
TASK_PP(16'h4D81,4);
TASK_PP(16'h4D82,4);
TASK_PP(16'h4D83,4);
TASK_PP(16'h4D84,4);
TASK_PP(16'h4D85,4);
TASK_PP(16'h4D86,4);
TASK_PP(16'h4D87,4);
TASK_PP(16'h4D88,4);
TASK_PP(16'h4D89,4);
TASK_PP(16'h4D8A,4);
TASK_PP(16'h4D8B,4);
TASK_PP(16'h4D8C,4);
TASK_PP(16'h4D8D,4);
TASK_PP(16'h4D8E,4);
TASK_PP(16'h4D8F,4);
TASK_PP(16'h4D90,4);
TASK_PP(16'h4D91,4);
TASK_PP(16'h4D92,4);
TASK_PP(16'h4D93,4);
TASK_PP(16'h4D94,4);
TASK_PP(16'h4D95,4);
TASK_PP(16'h4D96,4);
TASK_PP(16'h4D97,4);
TASK_PP(16'h4D98,4);
TASK_PP(16'h4D99,4);
TASK_PP(16'h4D9A,4);
TASK_PP(16'h4D9B,4);
TASK_PP(16'h4D9C,4);
TASK_PP(16'h4D9D,4);
TASK_PP(16'h4D9E,4);
TASK_PP(16'h4D9F,4);
TASK_PP(16'h4DA0,4);
TASK_PP(16'h4DA1,4);
TASK_PP(16'h4DA2,4);
TASK_PP(16'h4DA3,4);
TASK_PP(16'h4DA4,4);
TASK_PP(16'h4DA5,4);
TASK_PP(16'h4DA6,4);
TASK_PP(16'h4DA7,4);
TASK_PP(16'h4DA8,4);
TASK_PP(16'h4DA9,4);
TASK_PP(16'h4DAA,4);
TASK_PP(16'h4DAB,4);
TASK_PP(16'h4DAC,4);
TASK_PP(16'h4DAD,4);
TASK_PP(16'h4DAE,4);
TASK_PP(16'h4DAF,4);
TASK_PP(16'h4DB0,4);
TASK_PP(16'h4DB1,4);
TASK_PP(16'h4DB2,4);
TASK_PP(16'h4DB3,4);
TASK_PP(16'h4DB4,4);
TASK_PP(16'h4DB5,4);
TASK_PP(16'h4DB6,4);
TASK_PP(16'h4DB7,4);
TASK_PP(16'h4DB8,4);
TASK_PP(16'h4DB9,4);
TASK_PP(16'h4DBA,4);
TASK_PP(16'h4DBB,4);
TASK_PP(16'h4DBC,4);
TASK_PP(16'h4DBD,4);
TASK_PP(16'h4DBE,4);
TASK_PP(16'h4DBF,4);
TASK_PP(16'h4DC0,4);
TASK_PP(16'h4DC1,4);
TASK_PP(16'h4DC2,4);
TASK_PP(16'h4DC3,4);
TASK_PP(16'h4DC4,4);
TASK_PP(16'h4DC5,4);
TASK_PP(16'h4DC6,4);
TASK_PP(16'h4DC7,4);
TASK_PP(16'h4DC8,4);
TASK_PP(16'h4DC9,4);
TASK_PP(16'h4DCA,4);
TASK_PP(16'h4DCB,4);
TASK_PP(16'h4DCC,4);
TASK_PP(16'h4DCD,4);
TASK_PP(16'h4DCE,4);
TASK_PP(16'h4DCF,4);
TASK_PP(16'h4DD0,4);
TASK_PP(16'h4DD1,4);
TASK_PP(16'h4DD2,4);
TASK_PP(16'h4DD3,4);
TASK_PP(16'h4DD4,4);
TASK_PP(16'h4DD5,4);
TASK_PP(16'h4DD6,4);
TASK_PP(16'h4DD7,4);
TASK_PP(16'h4DD8,4);
TASK_PP(16'h4DD9,4);
TASK_PP(16'h4DDA,4);
TASK_PP(16'h4DDB,4);
TASK_PP(16'h4DDC,4);
TASK_PP(16'h4DDD,4);
TASK_PP(16'h4DDE,4);
TASK_PP(16'h4DDF,4);
TASK_PP(16'h4DE0,4);
TASK_PP(16'h4DE1,4);
TASK_PP(16'h4DE2,4);
TASK_PP(16'h4DE3,4);
TASK_PP(16'h4DE4,4);
TASK_PP(16'h4DE5,4);
TASK_PP(16'h4DE6,4);
TASK_PP(16'h4DE7,4);
TASK_PP(16'h4DE8,4);
TASK_PP(16'h4DE9,4);
TASK_PP(16'h4DEA,4);
TASK_PP(16'h4DEB,4);
TASK_PP(16'h4DEC,4);
TASK_PP(16'h4DED,4);
TASK_PP(16'h4DEE,4);
TASK_PP(16'h4DEF,4);
TASK_PP(16'h4DF0,4);
TASK_PP(16'h4DF1,4);
TASK_PP(16'h4DF2,4);
TASK_PP(16'h4DF3,4);
TASK_PP(16'h4DF4,4);
TASK_PP(16'h4DF5,4);
TASK_PP(16'h4DF6,4);
TASK_PP(16'h4DF7,4);
TASK_PP(16'h4DF8,4);
TASK_PP(16'h4DF9,4);
TASK_PP(16'h4DFA,4);
TASK_PP(16'h4DFB,4);
TASK_PP(16'h4DFC,4);
TASK_PP(16'h4DFD,4);
TASK_PP(16'h4DFE,4);
TASK_PP(16'h4DFF,4);
TASK_PP(16'h4E00,4);
TASK_PP(16'h4E01,4);
TASK_PP(16'h4E02,4);
TASK_PP(16'h4E03,4);
TASK_PP(16'h4E04,4);
TASK_PP(16'h4E05,4);
TASK_PP(16'h4E06,4);
TASK_PP(16'h4E07,4);
TASK_PP(16'h4E08,4);
TASK_PP(16'h4E09,4);
TASK_PP(16'h4E0A,4);
TASK_PP(16'h4E0B,4);
TASK_PP(16'h4E0C,4);
TASK_PP(16'h4E0D,4);
TASK_PP(16'h4E0E,4);
TASK_PP(16'h4E0F,4);
TASK_PP(16'h4E10,4);
TASK_PP(16'h4E11,4);
TASK_PP(16'h4E12,4);
TASK_PP(16'h4E13,4);
TASK_PP(16'h4E14,4);
TASK_PP(16'h4E15,4);
TASK_PP(16'h4E16,4);
TASK_PP(16'h4E17,4);
TASK_PP(16'h4E18,4);
TASK_PP(16'h4E19,4);
TASK_PP(16'h4E1A,4);
TASK_PP(16'h4E1B,4);
TASK_PP(16'h4E1C,4);
TASK_PP(16'h4E1D,4);
TASK_PP(16'h4E1E,4);
TASK_PP(16'h4E1F,4);
TASK_PP(16'h4E20,4);
TASK_PP(16'h4E21,4);
TASK_PP(16'h4E22,4);
TASK_PP(16'h4E23,4);
TASK_PP(16'h4E24,4);
TASK_PP(16'h4E25,4);
TASK_PP(16'h4E26,4);
TASK_PP(16'h4E27,4);
TASK_PP(16'h4E28,4);
TASK_PP(16'h4E29,4);
TASK_PP(16'h4E2A,4);
TASK_PP(16'h4E2B,4);
TASK_PP(16'h4E2C,4);
TASK_PP(16'h4E2D,4);
TASK_PP(16'h4E2E,4);
TASK_PP(16'h4E2F,4);
TASK_PP(16'h4E30,4);
TASK_PP(16'h4E31,4);
TASK_PP(16'h4E32,4);
TASK_PP(16'h4E33,4);
TASK_PP(16'h4E34,4);
TASK_PP(16'h4E35,4);
TASK_PP(16'h4E36,4);
TASK_PP(16'h4E37,4);
TASK_PP(16'h4E38,4);
TASK_PP(16'h4E39,4);
TASK_PP(16'h4E3A,4);
TASK_PP(16'h4E3B,4);
TASK_PP(16'h4E3C,4);
TASK_PP(16'h4E3D,4);
TASK_PP(16'h4E3E,4);
TASK_PP(16'h4E3F,4);
TASK_PP(16'h4E40,4);
TASK_PP(16'h4E41,4);
TASK_PP(16'h4E42,4);
TASK_PP(16'h4E43,4);
TASK_PP(16'h4E44,4);
TASK_PP(16'h4E45,4);
TASK_PP(16'h4E46,4);
TASK_PP(16'h4E47,4);
TASK_PP(16'h4E48,4);
TASK_PP(16'h4E49,4);
TASK_PP(16'h4E4A,4);
TASK_PP(16'h4E4B,4);
TASK_PP(16'h4E4C,4);
TASK_PP(16'h4E4D,4);
TASK_PP(16'h4E4E,4);
TASK_PP(16'h4E4F,4);
TASK_PP(16'h4E50,4);
TASK_PP(16'h4E51,4);
TASK_PP(16'h4E52,4);
TASK_PP(16'h4E53,4);
TASK_PP(16'h4E54,4);
TASK_PP(16'h4E55,4);
TASK_PP(16'h4E56,4);
TASK_PP(16'h4E57,4);
TASK_PP(16'h4E58,4);
TASK_PP(16'h4E59,4);
TASK_PP(16'h4E5A,4);
TASK_PP(16'h4E5B,4);
TASK_PP(16'h4E5C,4);
TASK_PP(16'h4E5D,4);
TASK_PP(16'h4E5E,4);
TASK_PP(16'h4E5F,4);
TASK_PP(16'h4E60,4);
TASK_PP(16'h4E61,4);
TASK_PP(16'h4E62,4);
TASK_PP(16'h4E63,4);
TASK_PP(16'h4E64,4);
TASK_PP(16'h4E65,4);
TASK_PP(16'h4E66,4);
TASK_PP(16'h4E67,4);
TASK_PP(16'h4E68,4);
TASK_PP(16'h4E69,4);
TASK_PP(16'h4E6A,4);
TASK_PP(16'h4E6B,4);
TASK_PP(16'h4E6C,4);
TASK_PP(16'h4E6D,4);
TASK_PP(16'h4E6E,4);
TASK_PP(16'h4E6F,4);
TASK_PP(16'h4E70,4);
TASK_PP(16'h4E71,4);
TASK_PP(16'h4E72,4);
TASK_PP(16'h4E73,4);
TASK_PP(16'h4E74,4);
TASK_PP(16'h4E75,4);
TASK_PP(16'h4E76,4);
TASK_PP(16'h4E77,4);
TASK_PP(16'h4E78,4);
TASK_PP(16'h4E79,4);
TASK_PP(16'h4E7A,4);
TASK_PP(16'h4E7B,4);
TASK_PP(16'h4E7C,4);
TASK_PP(16'h4E7D,4);
TASK_PP(16'h4E7E,4);
TASK_PP(16'h4E7F,4);
TASK_PP(16'h4E80,4);
TASK_PP(16'h4E81,4);
TASK_PP(16'h4E82,4);
TASK_PP(16'h4E83,4);
TASK_PP(16'h4E84,4);
TASK_PP(16'h4E85,4);
TASK_PP(16'h4E86,4);
TASK_PP(16'h4E87,4);
TASK_PP(16'h4E88,4);
TASK_PP(16'h4E89,4);
TASK_PP(16'h4E8A,4);
TASK_PP(16'h4E8B,4);
TASK_PP(16'h4E8C,4);
TASK_PP(16'h4E8D,4);
TASK_PP(16'h4E8E,4);
TASK_PP(16'h4E8F,4);
TASK_PP(16'h4E90,4);
TASK_PP(16'h4E91,4);
TASK_PP(16'h4E92,4);
TASK_PP(16'h4E93,4);
TASK_PP(16'h4E94,4);
TASK_PP(16'h4E95,4);
TASK_PP(16'h4E96,4);
TASK_PP(16'h4E97,4);
TASK_PP(16'h4E98,4);
TASK_PP(16'h4E99,4);
TASK_PP(16'h4E9A,4);
TASK_PP(16'h4E9B,4);
TASK_PP(16'h4E9C,4);
TASK_PP(16'h4E9D,4);
TASK_PP(16'h4E9E,4);
TASK_PP(16'h4E9F,4);
TASK_PP(16'h4EA0,4);
TASK_PP(16'h4EA1,4);
TASK_PP(16'h4EA2,4);
TASK_PP(16'h4EA3,4);
TASK_PP(16'h4EA4,4);
TASK_PP(16'h4EA5,4);
TASK_PP(16'h4EA6,4);
TASK_PP(16'h4EA7,4);
TASK_PP(16'h4EA8,4);
TASK_PP(16'h4EA9,4);
TASK_PP(16'h4EAA,4);
TASK_PP(16'h4EAB,4);
TASK_PP(16'h4EAC,4);
TASK_PP(16'h4EAD,4);
TASK_PP(16'h4EAE,4);
TASK_PP(16'h4EAF,4);
TASK_PP(16'h4EB0,4);
TASK_PP(16'h4EB1,4);
TASK_PP(16'h4EB2,4);
TASK_PP(16'h4EB3,4);
TASK_PP(16'h4EB4,4);
TASK_PP(16'h4EB5,4);
TASK_PP(16'h4EB6,4);
TASK_PP(16'h4EB7,4);
TASK_PP(16'h4EB8,4);
TASK_PP(16'h4EB9,4);
TASK_PP(16'h4EBA,4);
TASK_PP(16'h4EBB,4);
TASK_PP(16'h4EBC,4);
TASK_PP(16'h4EBD,4);
TASK_PP(16'h4EBE,4);
TASK_PP(16'h4EBF,4);
TASK_PP(16'h4EC0,4);
TASK_PP(16'h4EC1,4);
TASK_PP(16'h4EC2,4);
TASK_PP(16'h4EC3,4);
TASK_PP(16'h4EC4,4);
TASK_PP(16'h4EC5,4);
TASK_PP(16'h4EC6,4);
TASK_PP(16'h4EC7,4);
TASK_PP(16'h4EC8,4);
TASK_PP(16'h4EC9,4);
TASK_PP(16'h4ECA,4);
TASK_PP(16'h4ECB,4);
TASK_PP(16'h4ECC,4);
TASK_PP(16'h4ECD,4);
TASK_PP(16'h4ECE,4);
TASK_PP(16'h4ECF,4);
TASK_PP(16'h4ED0,4);
TASK_PP(16'h4ED1,4);
TASK_PP(16'h4ED2,4);
TASK_PP(16'h4ED3,4);
TASK_PP(16'h4ED4,4);
TASK_PP(16'h4ED5,4);
TASK_PP(16'h4ED6,4);
TASK_PP(16'h4ED7,4);
TASK_PP(16'h4ED8,4);
TASK_PP(16'h4ED9,4);
TASK_PP(16'h4EDA,4);
TASK_PP(16'h4EDB,4);
TASK_PP(16'h4EDC,4);
TASK_PP(16'h4EDD,4);
TASK_PP(16'h4EDE,4);
TASK_PP(16'h4EDF,4);
TASK_PP(16'h4EE0,4);
TASK_PP(16'h4EE1,4);
TASK_PP(16'h4EE2,4);
TASK_PP(16'h4EE3,4);
TASK_PP(16'h4EE4,4);
TASK_PP(16'h4EE5,4);
TASK_PP(16'h4EE6,4);
TASK_PP(16'h4EE7,4);
TASK_PP(16'h4EE8,4);
TASK_PP(16'h4EE9,4);
TASK_PP(16'h4EEA,4);
TASK_PP(16'h4EEB,4);
TASK_PP(16'h4EEC,4);
TASK_PP(16'h4EED,4);
TASK_PP(16'h4EEE,4);
TASK_PP(16'h4EEF,4);
TASK_PP(16'h4EF0,4);
TASK_PP(16'h4EF1,4);
TASK_PP(16'h4EF2,4);
TASK_PP(16'h4EF3,4);
TASK_PP(16'h4EF4,4);
TASK_PP(16'h4EF5,4);
TASK_PP(16'h4EF6,4);
TASK_PP(16'h4EF7,4);
TASK_PP(16'h4EF8,4);
TASK_PP(16'h4EF9,4);
TASK_PP(16'h4EFA,4);
TASK_PP(16'h4EFB,4);
TASK_PP(16'h4EFC,4);
TASK_PP(16'h4EFD,4);
TASK_PP(16'h4EFE,4);
TASK_PP(16'h4EFF,4);
TASK_PP(16'h4F00,4);
TASK_PP(16'h4F01,4);
TASK_PP(16'h4F02,4);
TASK_PP(16'h4F03,4);
TASK_PP(16'h4F04,4);
TASK_PP(16'h4F05,4);
TASK_PP(16'h4F06,4);
TASK_PP(16'h4F07,4);
TASK_PP(16'h4F08,4);
TASK_PP(16'h4F09,4);
TASK_PP(16'h4F0A,4);
TASK_PP(16'h4F0B,4);
TASK_PP(16'h4F0C,4);
TASK_PP(16'h4F0D,4);
TASK_PP(16'h4F0E,4);
TASK_PP(16'h4F0F,4);
TASK_PP(16'h4F10,4);
TASK_PP(16'h4F11,4);
TASK_PP(16'h4F12,4);
TASK_PP(16'h4F13,4);
TASK_PP(16'h4F14,4);
TASK_PP(16'h4F15,4);
TASK_PP(16'h4F16,4);
TASK_PP(16'h4F17,4);
TASK_PP(16'h4F18,4);
TASK_PP(16'h4F19,4);
TASK_PP(16'h4F1A,4);
TASK_PP(16'h4F1B,4);
TASK_PP(16'h4F1C,4);
TASK_PP(16'h4F1D,4);
TASK_PP(16'h4F1E,4);
TASK_PP(16'h4F1F,4);
TASK_PP(16'h4F20,4);
TASK_PP(16'h4F21,4);
TASK_PP(16'h4F22,4);
TASK_PP(16'h4F23,4);
TASK_PP(16'h4F24,4);
TASK_PP(16'h4F25,4);
TASK_PP(16'h4F26,4);
TASK_PP(16'h4F27,4);
TASK_PP(16'h4F28,4);
TASK_PP(16'h4F29,4);
TASK_PP(16'h4F2A,4);
TASK_PP(16'h4F2B,4);
TASK_PP(16'h4F2C,4);
TASK_PP(16'h4F2D,4);
TASK_PP(16'h4F2E,4);
TASK_PP(16'h4F2F,4);
TASK_PP(16'h4F30,4);
TASK_PP(16'h4F31,4);
TASK_PP(16'h4F32,4);
TASK_PP(16'h4F33,4);
TASK_PP(16'h4F34,4);
TASK_PP(16'h4F35,4);
TASK_PP(16'h4F36,4);
TASK_PP(16'h4F37,4);
TASK_PP(16'h4F38,4);
TASK_PP(16'h4F39,4);
TASK_PP(16'h4F3A,4);
TASK_PP(16'h4F3B,4);
TASK_PP(16'h4F3C,4);
TASK_PP(16'h4F3D,4);
TASK_PP(16'h4F3E,4);
TASK_PP(16'h4F3F,4);
TASK_PP(16'h4F40,4);
TASK_PP(16'h4F41,4);
TASK_PP(16'h4F42,4);
TASK_PP(16'h4F43,4);
TASK_PP(16'h4F44,4);
TASK_PP(16'h4F45,4);
TASK_PP(16'h4F46,4);
TASK_PP(16'h4F47,4);
TASK_PP(16'h4F48,4);
TASK_PP(16'h4F49,4);
TASK_PP(16'h4F4A,4);
TASK_PP(16'h4F4B,4);
TASK_PP(16'h4F4C,4);
TASK_PP(16'h4F4D,4);
TASK_PP(16'h4F4E,4);
TASK_PP(16'h4F4F,4);
TASK_PP(16'h4F50,4);
TASK_PP(16'h4F51,4);
TASK_PP(16'h4F52,4);
TASK_PP(16'h4F53,4);
TASK_PP(16'h4F54,4);
TASK_PP(16'h4F55,4);
TASK_PP(16'h4F56,4);
TASK_PP(16'h4F57,4);
TASK_PP(16'h4F58,4);
TASK_PP(16'h4F59,4);
TASK_PP(16'h4F5A,4);
TASK_PP(16'h4F5B,4);
TASK_PP(16'h4F5C,4);
TASK_PP(16'h4F5D,4);
TASK_PP(16'h4F5E,4);
TASK_PP(16'h4F5F,4);
TASK_PP(16'h4F60,4);
TASK_PP(16'h4F61,4);
TASK_PP(16'h4F62,4);
TASK_PP(16'h4F63,4);
TASK_PP(16'h4F64,4);
TASK_PP(16'h4F65,4);
TASK_PP(16'h4F66,4);
TASK_PP(16'h4F67,4);
TASK_PP(16'h4F68,4);
TASK_PP(16'h4F69,4);
TASK_PP(16'h4F6A,4);
TASK_PP(16'h4F6B,4);
TASK_PP(16'h4F6C,4);
TASK_PP(16'h4F6D,4);
TASK_PP(16'h4F6E,4);
TASK_PP(16'h4F6F,4);
TASK_PP(16'h4F70,4);
TASK_PP(16'h4F71,4);
TASK_PP(16'h4F72,4);
TASK_PP(16'h4F73,4);
TASK_PP(16'h4F74,4);
TASK_PP(16'h4F75,4);
TASK_PP(16'h4F76,4);
TASK_PP(16'h4F77,4);
TASK_PP(16'h4F78,4);
TASK_PP(16'h4F79,4);
TASK_PP(16'h4F7A,4);
TASK_PP(16'h4F7B,4);
TASK_PP(16'h4F7C,4);
TASK_PP(16'h4F7D,4);
TASK_PP(16'h4F7E,4);
TASK_PP(16'h4F7F,4);
TASK_PP(16'h4F80,4);
TASK_PP(16'h4F81,4);
TASK_PP(16'h4F82,4);
TASK_PP(16'h4F83,4);
TASK_PP(16'h4F84,4);
TASK_PP(16'h4F85,4);
TASK_PP(16'h4F86,4);
TASK_PP(16'h4F87,4);
TASK_PP(16'h4F88,4);
TASK_PP(16'h4F89,4);
TASK_PP(16'h4F8A,4);
TASK_PP(16'h4F8B,4);
TASK_PP(16'h4F8C,4);
TASK_PP(16'h4F8D,4);
TASK_PP(16'h4F8E,4);
TASK_PP(16'h4F8F,4);
TASK_PP(16'h4F90,4);
TASK_PP(16'h4F91,4);
TASK_PP(16'h4F92,4);
TASK_PP(16'h4F93,4);
TASK_PP(16'h4F94,4);
TASK_PP(16'h4F95,4);
TASK_PP(16'h4F96,4);
TASK_PP(16'h4F97,4);
TASK_PP(16'h4F98,4);
TASK_PP(16'h4F99,4);
TASK_PP(16'h4F9A,4);
TASK_PP(16'h4F9B,4);
TASK_PP(16'h4F9C,4);
TASK_PP(16'h4F9D,4);
TASK_PP(16'h4F9E,4);
TASK_PP(16'h4F9F,4);
TASK_PP(16'h4FA0,4);
TASK_PP(16'h4FA1,4);
TASK_PP(16'h4FA2,4);
TASK_PP(16'h4FA3,4);
TASK_PP(16'h4FA4,4);
TASK_PP(16'h4FA5,4);
TASK_PP(16'h4FA6,4);
TASK_PP(16'h4FA7,4);
TASK_PP(16'h4FA8,4);
TASK_PP(16'h4FA9,4);
TASK_PP(16'h4FAA,4);
TASK_PP(16'h4FAB,4);
TASK_PP(16'h4FAC,4);
TASK_PP(16'h4FAD,4);
TASK_PP(16'h4FAE,4);
TASK_PP(16'h4FAF,4);
TASK_PP(16'h4FB0,4);
TASK_PP(16'h4FB1,4);
TASK_PP(16'h4FB2,4);
TASK_PP(16'h4FB3,4);
TASK_PP(16'h4FB4,4);
TASK_PP(16'h4FB5,4);
TASK_PP(16'h4FB6,4);
TASK_PP(16'h4FB7,4);
TASK_PP(16'h4FB8,4);
TASK_PP(16'h4FB9,4);
TASK_PP(16'h4FBA,4);
TASK_PP(16'h4FBB,4);
TASK_PP(16'h4FBC,4);
TASK_PP(16'h4FBD,4);
TASK_PP(16'h4FBE,4);
TASK_PP(16'h4FBF,4);
TASK_PP(16'h4FC0,4);
TASK_PP(16'h4FC1,4);
TASK_PP(16'h4FC2,4);
TASK_PP(16'h4FC3,4);
TASK_PP(16'h4FC4,4);
TASK_PP(16'h4FC5,4);
TASK_PP(16'h4FC6,4);
TASK_PP(16'h4FC7,4);
TASK_PP(16'h4FC8,4);
TASK_PP(16'h4FC9,4);
TASK_PP(16'h4FCA,4);
TASK_PP(16'h4FCB,4);
TASK_PP(16'h4FCC,4);
TASK_PP(16'h4FCD,4);
TASK_PP(16'h4FCE,4);
TASK_PP(16'h4FCF,4);
TASK_PP(16'h4FD0,4);
TASK_PP(16'h4FD1,4);
TASK_PP(16'h4FD2,4);
TASK_PP(16'h4FD3,4);
TASK_PP(16'h4FD4,4);
TASK_PP(16'h4FD5,4);
TASK_PP(16'h4FD6,4);
TASK_PP(16'h4FD7,4);
TASK_PP(16'h4FD8,4);
TASK_PP(16'h4FD9,4);
TASK_PP(16'h4FDA,4);
TASK_PP(16'h4FDB,4);
TASK_PP(16'h4FDC,4);
TASK_PP(16'h4FDD,4);
TASK_PP(16'h4FDE,4);
TASK_PP(16'h4FDF,4);
TASK_PP(16'h4FE0,4);
TASK_PP(16'h4FE1,4);
TASK_PP(16'h4FE2,4);
TASK_PP(16'h4FE3,4);
TASK_PP(16'h4FE4,4);
TASK_PP(16'h4FE5,4);
TASK_PP(16'h4FE6,4);
TASK_PP(16'h4FE7,4);
TASK_PP(16'h4FE8,4);
TASK_PP(16'h4FE9,4);
TASK_PP(16'h4FEA,4);
TASK_PP(16'h4FEB,4);
TASK_PP(16'h4FEC,4);
TASK_PP(16'h4FED,4);
TASK_PP(16'h4FEE,4);
TASK_PP(16'h4FEF,4);
TASK_PP(16'h4FF0,4);
TASK_PP(16'h4FF1,4);
TASK_PP(16'h4FF2,4);
TASK_PP(16'h4FF3,4);
TASK_PP(16'h4FF4,4);
TASK_PP(16'h4FF5,4);
TASK_PP(16'h4FF6,4);
TASK_PP(16'h4FF7,4);
TASK_PP(16'h4FF8,4);
TASK_PP(16'h4FF9,4);
TASK_PP(16'h4FFA,4);
TASK_PP(16'h4FFB,4);
TASK_PP(16'h4FFC,4);
TASK_PP(16'h4FFD,4);
TASK_PP(16'h4FFE,4);
TASK_PP(16'h4FFF,4);
TASK_PP(16'h5000,4);
TASK_PP(16'h5001,4);
TASK_PP(16'h5002,4);
TASK_PP(16'h5003,4);
TASK_PP(16'h5004,4);
TASK_PP(16'h5005,4);
TASK_PP(16'h5006,4);
TASK_PP(16'h5007,4);
TASK_PP(16'h5008,4);
TASK_PP(16'h5009,4);
TASK_PP(16'h500A,4);
TASK_PP(16'h500B,4);
TASK_PP(16'h500C,4);
TASK_PP(16'h500D,4);
TASK_PP(16'h500E,4);
TASK_PP(16'h500F,4);
TASK_PP(16'h5010,4);
TASK_PP(16'h5011,4);
TASK_PP(16'h5012,4);
TASK_PP(16'h5013,4);
TASK_PP(16'h5014,4);
TASK_PP(16'h5015,4);
TASK_PP(16'h5016,4);
TASK_PP(16'h5017,4);
TASK_PP(16'h5018,4);
TASK_PP(16'h5019,4);
TASK_PP(16'h501A,4);
TASK_PP(16'h501B,4);
TASK_PP(16'h501C,4);
TASK_PP(16'h501D,4);
TASK_PP(16'h501E,4);
TASK_PP(16'h501F,4);
TASK_PP(16'h5020,4);
TASK_PP(16'h5021,4);
TASK_PP(16'h5022,4);
TASK_PP(16'h5023,4);
TASK_PP(16'h5024,4);
TASK_PP(16'h5025,4);
TASK_PP(16'h5026,4);
TASK_PP(16'h5027,4);
TASK_PP(16'h5028,4);
TASK_PP(16'h5029,4);
TASK_PP(16'h502A,4);
TASK_PP(16'h502B,4);
TASK_PP(16'h502C,4);
TASK_PP(16'h502D,4);
TASK_PP(16'h502E,4);
TASK_PP(16'h502F,4);
TASK_PP(16'h5030,4);
TASK_PP(16'h5031,4);
TASK_PP(16'h5032,4);
TASK_PP(16'h5033,4);
TASK_PP(16'h5034,4);
TASK_PP(16'h5035,4);
TASK_PP(16'h5036,4);
TASK_PP(16'h5037,4);
TASK_PP(16'h5038,4);
TASK_PP(16'h5039,4);
TASK_PP(16'h503A,4);
TASK_PP(16'h503B,4);
TASK_PP(16'h503C,4);
TASK_PP(16'h503D,4);
TASK_PP(16'h503E,4);
TASK_PP(16'h503F,4);
TASK_PP(16'h5040,4);
TASK_PP(16'h5041,4);
TASK_PP(16'h5042,4);
TASK_PP(16'h5043,4);
TASK_PP(16'h5044,4);
TASK_PP(16'h5045,4);
TASK_PP(16'h5046,4);
TASK_PP(16'h5047,4);
TASK_PP(16'h5048,4);
TASK_PP(16'h5049,4);
TASK_PP(16'h504A,4);
TASK_PP(16'h504B,4);
TASK_PP(16'h504C,4);
TASK_PP(16'h504D,4);
TASK_PP(16'h504E,4);
TASK_PP(16'h504F,4);
TASK_PP(16'h5050,4);
TASK_PP(16'h5051,4);
TASK_PP(16'h5052,4);
TASK_PP(16'h5053,4);
TASK_PP(16'h5054,4);
TASK_PP(16'h5055,4);
TASK_PP(16'h5056,4);
TASK_PP(16'h5057,4);
TASK_PP(16'h5058,4);
TASK_PP(16'h5059,4);
TASK_PP(16'h505A,4);
TASK_PP(16'h505B,4);
TASK_PP(16'h505C,4);
TASK_PP(16'h505D,4);
TASK_PP(16'h505E,4);
TASK_PP(16'h505F,4);
TASK_PP(16'h5060,4);
TASK_PP(16'h5061,4);
TASK_PP(16'h5062,4);
TASK_PP(16'h5063,4);
TASK_PP(16'h5064,4);
TASK_PP(16'h5065,4);
TASK_PP(16'h5066,4);
TASK_PP(16'h5067,4);
TASK_PP(16'h5068,4);
TASK_PP(16'h5069,4);
TASK_PP(16'h506A,4);
TASK_PP(16'h506B,4);
TASK_PP(16'h506C,4);
TASK_PP(16'h506D,4);
TASK_PP(16'h506E,4);
TASK_PP(16'h506F,4);
TASK_PP(16'h5070,4);
TASK_PP(16'h5071,4);
TASK_PP(16'h5072,4);
TASK_PP(16'h5073,4);
TASK_PP(16'h5074,4);
TASK_PP(16'h5075,4);
TASK_PP(16'h5076,4);
TASK_PP(16'h5077,4);
TASK_PP(16'h5078,4);
TASK_PP(16'h5079,4);
TASK_PP(16'h507A,4);
TASK_PP(16'h507B,4);
TASK_PP(16'h507C,4);
TASK_PP(16'h507D,4);
TASK_PP(16'h507E,4);
TASK_PP(16'h507F,4);
TASK_PP(16'h5080,4);
TASK_PP(16'h5081,4);
TASK_PP(16'h5082,4);
TASK_PP(16'h5083,4);
TASK_PP(16'h5084,4);
TASK_PP(16'h5085,4);
TASK_PP(16'h5086,4);
TASK_PP(16'h5087,4);
TASK_PP(16'h5088,4);
TASK_PP(16'h5089,4);
TASK_PP(16'h508A,4);
TASK_PP(16'h508B,4);
TASK_PP(16'h508C,4);
TASK_PP(16'h508D,4);
TASK_PP(16'h508E,4);
TASK_PP(16'h508F,4);
TASK_PP(16'h5090,4);
TASK_PP(16'h5091,4);
TASK_PP(16'h5092,4);
TASK_PP(16'h5093,4);
TASK_PP(16'h5094,4);
TASK_PP(16'h5095,4);
TASK_PP(16'h5096,4);
TASK_PP(16'h5097,4);
TASK_PP(16'h5098,4);
TASK_PP(16'h5099,4);
TASK_PP(16'h509A,4);
TASK_PP(16'h509B,4);
TASK_PP(16'h509C,4);
TASK_PP(16'h509D,4);
TASK_PP(16'h509E,4);
TASK_PP(16'h509F,4);
TASK_PP(16'h50A0,4);
TASK_PP(16'h50A1,4);
TASK_PP(16'h50A2,4);
TASK_PP(16'h50A3,4);
TASK_PP(16'h50A4,4);
TASK_PP(16'h50A5,4);
TASK_PP(16'h50A6,4);
TASK_PP(16'h50A7,4);
TASK_PP(16'h50A8,4);
TASK_PP(16'h50A9,4);
TASK_PP(16'h50AA,4);
TASK_PP(16'h50AB,4);
TASK_PP(16'h50AC,4);
TASK_PP(16'h50AD,4);
TASK_PP(16'h50AE,4);
TASK_PP(16'h50AF,4);
TASK_PP(16'h50B0,4);
TASK_PP(16'h50B1,4);
TASK_PP(16'h50B2,4);
TASK_PP(16'h50B3,4);
TASK_PP(16'h50B4,4);
TASK_PP(16'h50B5,4);
TASK_PP(16'h50B6,4);
TASK_PP(16'h50B7,4);
TASK_PP(16'h50B8,4);
TASK_PP(16'h50B9,4);
TASK_PP(16'h50BA,4);
TASK_PP(16'h50BB,4);
TASK_PP(16'h50BC,4);
TASK_PP(16'h50BD,4);
TASK_PP(16'h50BE,4);
TASK_PP(16'h50BF,4);
TASK_PP(16'h50C0,4);
TASK_PP(16'h50C1,4);
TASK_PP(16'h50C2,4);
TASK_PP(16'h50C3,4);
TASK_PP(16'h50C4,4);
TASK_PP(16'h50C5,4);
TASK_PP(16'h50C6,4);
TASK_PP(16'h50C7,4);
TASK_PP(16'h50C8,4);
TASK_PP(16'h50C9,4);
TASK_PP(16'h50CA,4);
TASK_PP(16'h50CB,4);
TASK_PP(16'h50CC,4);
TASK_PP(16'h50CD,4);
TASK_PP(16'h50CE,4);
TASK_PP(16'h50CF,4);
TASK_PP(16'h50D0,4);
TASK_PP(16'h50D1,4);
TASK_PP(16'h50D2,4);
TASK_PP(16'h50D3,4);
TASK_PP(16'h50D4,4);
TASK_PP(16'h50D5,4);
TASK_PP(16'h50D6,4);
TASK_PP(16'h50D7,4);
TASK_PP(16'h50D8,4);
TASK_PP(16'h50D9,4);
TASK_PP(16'h50DA,4);
TASK_PP(16'h50DB,4);
TASK_PP(16'h50DC,4);
TASK_PP(16'h50DD,4);
TASK_PP(16'h50DE,4);
TASK_PP(16'h50DF,4);
TASK_PP(16'h50E0,4);
TASK_PP(16'h50E1,4);
TASK_PP(16'h50E2,4);
TASK_PP(16'h50E3,4);
TASK_PP(16'h50E4,4);
TASK_PP(16'h50E5,4);
TASK_PP(16'h50E6,4);
TASK_PP(16'h50E7,4);
TASK_PP(16'h50E8,4);
TASK_PP(16'h50E9,4);
TASK_PP(16'h50EA,4);
TASK_PP(16'h50EB,4);
TASK_PP(16'h50EC,4);
TASK_PP(16'h50ED,4);
TASK_PP(16'h50EE,4);
TASK_PP(16'h50EF,4);
TASK_PP(16'h50F0,4);
TASK_PP(16'h50F1,4);
TASK_PP(16'h50F2,4);
TASK_PP(16'h50F3,4);
TASK_PP(16'h50F4,4);
TASK_PP(16'h50F5,4);
TASK_PP(16'h50F6,4);
TASK_PP(16'h50F7,4);
TASK_PP(16'h50F8,4);
TASK_PP(16'h50F9,4);
TASK_PP(16'h50FA,4);
TASK_PP(16'h50FB,4);
TASK_PP(16'h50FC,4);
TASK_PP(16'h50FD,4);
TASK_PP(16'h50FE,4);
TASK_PP(16'h50FF,4);
TASK_PP(16'h5100,4);
TASK_PP(16'h5101,4);
TASK_PP(16'h5102,4);
TASK_PP(16'h5103,4);
TASK_PP(16'h5104,4);
TASK_PP(16'h5105,4);
TASK_PP(16'h5106,4);
TASK_PP(16'h5107,4);
TASK_PP(16'h5108,4);
TASK_PP(16'h5109,4);
TASK_PP(16'h510A,4);
TASK_PP(16'h510B,4);
TASK_PP(16'h510C,4);
TASK_PP(16'h510D,4);
TASK_PP(16'h510E,4);
TASK_PP(16'h510F,4);
TASK_PP(16'h5110,4);
TASK_PP(16'h5111,4);
TASK_PP(16'h5112,4);
TASK_PP(16'h5113,4);
TASK_PP(16'h5114,4);
TASK_PP(16'h5115,4);
TASK_PP(16'h5116,4);
TASK_PP(16'h5117,4);
TASK_PP(16'h5118,4);
TASK_PP(16'h5119,4);
TASK_PP(16'h511A,4);
TASK_PP(16'h511B,4);
TASK_PP(16'h511C,4);
TASK_PP(16'h511D,4);
TASK_PP(16'h511E,4);
TASK_PP(16'h511F,4);
TASK_PP(16'h5120,4);
TASK_PP(16'h5121,4);
TASK_PP(16'h5122,4);
TASK_PP(16'h5123,4);
TASK_PP(16'h5124,4);
TASK_PP(16'h5125,4);
TASK_PP(16'h5126,4);
TASK_PP(16'h5127,4);
TASK_PP(16'h5128,4);
TASK_PP(16'h5129,4);
TASK_PP(16'h512A,4);
TASK_PP(16'h512B,4);
TASK_PP(16'h512C,4);
TASK_PP(16'h512D,4);
TASK_PP(16'h512E,4);
TASK_PP(16'h512F,4);
TASK_PP(16'h5130,4);
TASK_PP(16'h5131,4);
TASK_PP(16'h5132,4);
TASK_PP(16'h5133,4);
TASK_PP(16'h5134,4);
TASK_PP(16'h5135,4);
TASK_PP(16'h5136,4);
TASK_PP(16'h5137,4);
TASK_PP(16'h5138,4);
TASK_PP(16'h5139,4);
TASK_PP(16'h513A,4);
TASK_PP(16'h513B,4);
TASK_PP(16'h513C,4);
TASK_PP(16'h513D,4);
TASK_PP(16'h513E,4);
TASK_PP(16'h513F,4);
TASK_PP(16'h5140,4);
TASK_PP(16'h5141,4);
TASK_PP(16'h5142,4);
TASK_PP(16'h5143,4);
TASK_PP(16'h5144,4);
TASK_PP(16'h5145,4);
TASK_PP(16'h5146,4);
TASK_PP(16'h5147,4);
TASK_PP(16'h5148,4);
TASK_PP(16'h5149,4);
TASK_PP(16'h514A,4);
TASK_PP(16'h514B,4);
TASK_PP(16'h514C,4);
TASK_PP(16'h514D,4);
TASK_PP(16'h514E,4);
TASK_PP(16'h514F,4);
TASK_PP(16'h5150,4);
TASK_PP(16'h5151,4);
TASK_PP(16'h5152,4);
TASK_PP(16'h5153,4);
TASK_PP(16'h5154,4);
TASK_PP(16'h5155,4);
TASK_PP(16'h5156,4);
TASK_PP(16'h5157,4);
TASK_PP(16'h5158,4);
TASK_PP(16'h5159,4);
TASK_PP(16'h515A,4);
TASK_PP(16'h515B,4);
TASK_PP(16'h515C,4);
TASK_PP(16'h515D,4);
TASK_PP(16'h515E,4);
TASK_PP(16'h515F,4);
TASK_PP(16'h5160,4);
TASK_PP(16'h5161,4);
TASK_PP(16'h5162,4);
TASK_PP(16'h5163,4);
TASK_PP(16'h5164,4);
TASK_PP(16'h5165,4);
TASK_PP(16'h5166,4);
TASK_PP(16'h5167,4);
TASK_PP(16'h5168,4);
TASK_PP(16'h5169,4);
TASK_PP(16'h516A,4);
TASK_PP(16'h516B,4);
TASK_PP(16'h516C,4);
TASK_PP(16'h516D,4);
TASK_PP(16'h516E,4);
TASK_PP(16'h516F,4);
TASK_PP(16'h5170,4);
TASK_PP(16'h5171,4);
TASK_PP(16'h5172,4);
TASK_PP(16'h5173,4);
TASK_PP(16'h5174,4);
TASK_PP(16'h5175,4);
TASK_PP(16'h5176,4);
TASK_PP(16'h5177,4);
TASK_PP(16'h5178,4);
TASK_PP(16'h5179,4);
TASK_PP(16'h517A,4);
TASK_PP(16'h517B,4);
TASK_PP(16'h517C,4);
TASK_PP(16'h517D,4);
TASK_PP(16'h517E,4);
TASK_PP(16'h517F,4);
TASK_PP(16'h5180,4);
TASK_PP(16'h5181,4);
TASK_PP(16'h5182,4);
TASK_PP(16'h5183,4);
TASK_PP(16'h5184,4);
TASK_PP(16'h5185,4);
TASK_PP(16'h5186,4);
TASK_PP(16'h5187,4);
TASK_PP(16'h5188,4);
TASK_PP(16'h5189,4);
TASK_PP(16'h518A,4);
TASK_PP(16'h518B,4);
TASK_PP(16'h518C,4);
TASK_PP(16'h518D,4);
TASK_PP(16'h518E,4);
TASK_PP(16'h518F,4);
TASK_PP(16'h5190,4);
TASK_PP(16'h5191,4);
TASK_PP(16'h5192,4);
TASK_PP(16'h5193,4);
TASK_PP(16'h5194,4);
TASK_PP(16'h5195,4);
TASK_PP(16'h5196,4);
TASK_PP(16'h5197,4);
TASK_PP(16'h5198,4);
TASK_PP(16'h5199,4);
TASK_PP(16'h519A,4);
TASK_PP(16'h519B,4);
TASK_PP(16'h519C,4);
TASK_PP(16'h519D,4);
TASK_PP(16'h519E,4);
TASK_PP(16'h519F,4);
TASK_PP(16'h51A0,4);
TASK_PP(16'h51A1,4);
TASK_PP(16'h51A2,4);
TASK_PP(16'h51A3,4);
TASK_PP(16'h51A4,4);
TASK_PP(16'h51A5,4);
TASK_PP(16'h51A6,4);
TASK_PP(16'h51A7,4);
TASK_PP(16'h51A8,4);
TASK_PP(16'h51A9,4);
TASK_PP(16'h51AA,4);
TASK_PP(16'h51AB,4);
TASK_PP(16'h51AC,4);
TASK_PP(16'h51AD,4);
TASK_PP(16'h51AE,4);
TASK_PP(16'h51AF,4);
TASK_PP(16'h51B0,4);
TASK_PP(16'h51B1,4);
TASK_PP(16'h51B2,4);
TASK_PP(16'h51B3,4);
TASK_PP(16'h51B4,4);
TASK_PP(16'h51B5,4);
TASK_PP(16'h51B6,4);
TASK_PP(16'h51B7,4);
TASK_PP(16'h51B8,4);
TASK_PP(16'h51B9,4);
TASK_PP(16'h51BA,4);
TASK_PP(16'h51BB,4);
TASK_PP(16'h51BC,4);
TASK_PP(16'h51BD,4);
TASK_PP(16'h51BE,4);
TASK_PP(16'h51BF,4);
TASK_PP(16'h51C0,4);
TASK_PP(16'h51C1,4);
TASK_PP(16'h51C2,4);
TASK_PP(16'h51C3,4);
TASK_PP(16'h51C4,4);
TASK_PP(16'h51C5,4);
TASK_PP(16'h51C6,4);
TASK_PP(16'h51C7,4);
TASK_PP(16'h51C8,4);
TASK_PP(16'h51C9,4);
TASK_PP(16'h51CA,4);
TASK_PP(16'h51CB,4);
TASK_PP(16'h51CC,4);
TASK_PP(16'h51CD,4);
TASK_PP(16'h51CE,4);
TASK_PP(16'h51CF,4);
TASK_PP(16'h51D0,4);
TASK_PP(16'h51D1,4);
TASK_PP(16'h51D2,4);
TASK_PP(16'h51D3,4);
TASK_PP(16'h51D4,4);
TASK_PP(16'h51D5,4);
TASK_PP(16'h51D6,4);
TASK_PP(16'h51D7,4);
TASK_PP(16'h51D8,4);
TASK_PP(16'h51D9,4);
TASK_PP(16'h51DA,4);
TASK_PP(16'h51DB,4);
TASK_PP(16'h51DC,4);
TASK_PP(16'h51DD,4);
TASK_PP(16'h51DE,4);
TASK_PP(16'h51DF,4);
TASK_PP(16'h51E0,4);
TASK_PP(16'h51E1,4);
TASK_PP(16'h51E2,4);
TASK_PP(16'h51E3,4);
TASK_PP(16'h51E4,4);
TASK_PP(16'h51E5,4);
TASK_PP(16'h51E6,4);
TASK_PP(16'h51E7,4);
TASK_PP(16'h51E8,4);
TASK_PP(16'h51E9,4);
TASK_PP(16'h51EA,4);
TASK_PP(16'h51EB,4);
TASK_PP(16'h51EC,4);
TASK_PP(16'h51ED,4);
TASK_PP(16'h51EE,4);
TASK_PP(16'h51EF,4);
TASK_PP(16'h51F0,4);
TASK_PP(16'h51F1,4);
TASK_PP(16'h51F2,4);
TASK_PP(16'h51F3,4);
TASK_PP(16'h51F4,4);
TASK_PP(16'h51F5,4);
TASK_PP(16'h51F6,4);
TASK_PP(16'h51F7,4);
TASK_PP(16'h51F8,4);
TASK_PP(16'h51F9,4);
TASK_PP(16'h51FA,4);
TASK_PP(16'h51FB,4);
TASK_PP(16'h51FC,4);
TASK_PP(16'h51FD,4);
TASK_PP(16'h51FE,4);
TASK_PP(16'h51FF,4);
TASK_PP(16'h5200,4);
TASK_PP(16'h5201,4);
TASK_PP(16'h5202,4);
TASK_PP(16'h5203,4);
TASK_PP(16'h5204,4);
TASK_PP(16'h5205,4);
TASK_PP(16'h5206,4);
TASK_PP(16'h5207,4);
TASK_PP(16'h5208,4);
TASK_PP(16'h5209,4);
TASK_PP(16'h520A,4);
TASK_PP(16'h520B,4);
TASK_PP(16'h520C,4);
TASK_PP(16'h520D,4);
TASK_PP(16'h520E,4);
TASK_PP(16'h520F,4);
TASK_PP(16'h5210,4);
TASK_PP(16'h5211,4);
TASK_PP(16'h5212,4);
TASK_PP(16'h5213,4);
TASK_PP(16'h5214,4);
TASK_PP(16'h5215,4);
TASK_PP(16'h5216,4);
TASK_PP(16'h5217,4);
TASK_PP(16'h5218,4);
TASK_PP(16'h5219,4);
TASK_PP(16'h521A,4);
TASK_PP(16'h521B,4);
TASK_PP(16'h521C,4);
TASK_PP(16'h521D,4);
TASK_PP(16'h521E,4);
TASK_PP(16'h521F,4);
TASK_PP(16'h5220,4);
TASK_PP(16'h5221,4);
TASK_PP(16'h5222,4);
TASK_PP(16'h5223,4);
TASK_PP(16'h5224,4);
TASK_PP(16'h5225,4);
TASK_PP(16'h5226,4);
TASK_PP(16'h5227,4);
TASK_PP(16'h5228,4);
TASK_PP(16'h5229,4);
TASK_PP(16'h522A,4);
TASK_PP(16'h522B,4);
TASK_PP(16'h522C,4);
TASK_PP(16'h522D,4);
TASK_PP(16'h522E,4);
TASK_PP(16'h522F,4);
TASK_PP(16'h5230,4);
TASK_PP(16'h5231,4);
TASK_PP(16'h5232,4);
TASK_PP(16'h5233,4);
TASK_PP(16'h5234,4);
TASK_PP(16'h5235,4);
TASK_PP(16'h5236,4);
TASK_PP(16'h5237,4);
TASK_PP(16'h5238,4);
TASK_PP(16'h5239,4);
TASK_PP(16'h523A,4);
TASK_PP(16'h523B,4);
TASK_PP(16'h523C,4);
TASK_PP(16'h523D,4);
TASK_PP(16'h523E,4);
TASK_PP(16'h523F,4);
TASK_PP(16'h5240,4);
TASK_PP(16'h5241,4);
TASK_PP(16'h5242,4);
TASK_PP(16'h5243,4);
TASK_PP(16'h5244,4);
TASK_PP(16'h5245,4);
TASK_PP(16'h5246,4);
TASK_PP(16'h5247,4);
TASK_PP(16'h5248,4);
TASK_PP(16'h5249,4);
TASK_PP(16'h524A,4);
TASK_PP(16'h524B,4);
TASK_PP(16'h524C,4);
TASK_PP(16'h524D,4);
TASK_PP(16'h524E,4);
TASK_PP(16'h524F,4);
TASK_PP(16'h5250,4);
TASK_PP(16'h5251,4);
TASK_PP(16'h5252,4);
TASK_PP(16'h5253,4);
TASK_PP(16'h5254,4);
TASK_PP(16'h5255,4);
TASK_PP(16'h5256,4);
TASK_PP(16'h5257,4);
TASK_PP(16'h5258,4);
TASK_PP(16'h5259,4);
TASK_PP(16'h525A,4);
TASK_PP(16'h525B,4);
TASK_PP(16'h525C,4);
TASK_PP(16'h525D,4);
TASK_PP(16'h525E,4);
TASK_PP(16'h525F,4);
TASK_PP(16'h5260,4);
TASK_PP(16'h5261,4);
TASK_PP(16'h5262,4);
TASK_PP(16'h5263,4);
TASK_PP(16'h5264,4);
TASK_PP(16'h5265,4);
TASK_PP(16'h5266,4);
TASK_PP(16'h5267,4);
TASK_PP(16'h5268,4);
TASK_PP(16'h5269,4);
TASK_PP(16'h526A,4);
TASK_PP(16'h526B,4);
TASK_PP(16'h526C,4);
TASK_PP(16'h526D,4);
TASK_PP(16'h526E,4);
TASK_PP(16'h526F,4);
TASK_PP(16'h5270,4);
TASK_PP(16'h5271,4);
TASK_PP(16'h5272,4);
TASK_PP(16'h5273,4);
TASK_PP(16'h5274,4);
TASK_PP(16'h5275,4);
TASK_PP(16'h5276,4);
TASK_PP(16'h5277,4);
TASK_PP(16'h5278,4);
TASK_PP(16'h5279,4);
TASK_PP(16'h527A,4);
TASK_PP(16'h527B,4);
TASK_PP(16'h527C,4);
TASK_PP(16'h527D,4);
TASK_PP(16'h527E,4);
TASK_PP(16'h527F,4);
TASK_PP(16'h5280,4);
TASK_PP(16'h5281,4);
TASK_PP(16'h5282,4);
TASK_PP(16'h5283,4);
TASK_PP(16'h5284,4);
TASK_PP(16'h5285,4);
TASK_PP(16'h5286,4);
TASK_PP(16'h5287,4);
TASK_PP(16'h5288,4);
TASK_PP(16'h5289,4);
TASK_PP(16'h528A,4);
TASK_PP(16'h528B,4);
TASK_PP(16'h528C,4);
TASK_PP(16'h528D,4);
TASK_PP(16'h528E,4);
TASK_PP(16'h528F,4);
TASK_PP(16'h5290,4);
TASK_PP(16'h5291,4);
TASK_PP(16'h5292,4);
TASK_PP(16'h5293,4);
TASK_PP(16'h5294,4);
TASK_PP(16'h5295,4);
TASK_PP(16'h5296,4);
TASK_PP(16'h5297,4);
TASK_PP(16'h5298,4);
TASK_PP(16'h5299,4);
TASK_PP(16'h529A,4);
TASK_PP(16'h529B,4);
TASK_PP(16'h529C,4);
TASK_PP(16'h529D,4);
TASK_PP(16'h529E,4);
TASK_PP(16'h529F,4);
TASK_PP(16'h52A0,4);
TASK_PP(16'h52A1,4);
TASK_PP(16'h52A2,4);
TASK_PP(16'h52A3,4);
TASK_PP(16'h52A4,4);
TASK_PP(16'h52A5,4);
TASK_PP(16'h52A6,4);
TASK_PP(16'h52A7,4);
TASK_PP(16'h52A8,4);
TASK_PP(16'h52A9,4);
TASK_PP(16'h52AA,4);
TASK_PP(16'h52AB,4);
TASK_PP(16'h52AC,4);
TASK_PP(16'h52AD,4);
TASK_PP(16'h52AE,4);
TASK_PP(16'h52AF,4);
TASK_PP(16'h52B0,4);
TASK_PP(16'h52B1,4);
TASK_PP(16'h52B2,4);
TASK_PP(16'h52B3,4);
TASK_PP(16'h52B4,4);
TASK_PP(16'h52B5,4);
TASK_PP(16'h52B6,4);
TASK_PP(16'h52B7,4);
TASK_PP(16'h52B8,4);
TASK_PP(16'h52B9,4);
TASK_PP(16'h52BA,4);
TASK_PP(16'h52BB,4);
TASK_PP(16'h52BC,4);
TASK_PP(16'h52BD,4);
TASK_PP(16'h52BE,4);
TASK_PP(16'h52BF,4);
TASK_PP(16'h52C0,4);
TASK_PP(16'h52C1,4);
TASK_PP(16'h52C2,4);
TASK_PP(16'h52C3,4);
TASK_PP(16'h52C4,4);
TASK_PP(16'h52C5,4);
TASK_PP(16'h52C6,4);
TASK_PP(16'h52C7,4);
TASK_PP(16'h52C8,4);
TASK_PP(16'h52C9,4);
TASK_PP(16'h52CA,4);
TASK_PP(16'h52CB,4);
TASK_PP(16'h52CC,4);
TASK_PP(16'h52CD,4);
TASK_PP(16'h52CE,4);
TASK_PP(16'h52CF,4);
TASK_PP(16'h52D0,4);
TASK_PP(16'h52D1,4);
TASK_PP(16'h52D2,4);
TASK_PP(16'h52D3,4);
TASK_PP(16'h52D4,4);
TASK_PP(16'h52D5,4);
TASK_PP(16'h52D6,4);
TASK_PP(16'h52D7,4);
TASK_PP(16'h52D8,4);
TASK_PP(16'h52D9,4);
TASK_PP(16'h52DA,4);
TASK_PP(16'h52DB,4);
TASK_PP(16'h52DC,4);
TASK_PP(16'h52DD,4);
TASK_PP(16'h52DE,4);
TASK_PP(16'h52DF,4);
TASK_PP(16'h52E0,4);
TASK_PP(16'h52E1,4);
TASK_PP(16'h52E2,4);
TASK_PP(16'h52E3,4);
TASK_PP(16'h52E4,4);
TASK_PP(16'h52E5,4);
TASK_PP(16'h52E6,4);
TASK_PP(16'h52E7,4);
TASK_PP(16'h52E8,4);
TASK_PP(16'h52E9,4);
TASK_PP(16'h52EA,4);
TASK_PP(16'h52EB,4);
TASK_PP(16'h52EC,4);
TASK_PP(16'h52ED,4);
TASK_PP(16'h52EE,4);
TASK_PP(16'h52EF,4);
TASK_PP(16'h52F0,4);
TASK_PP(16'h52F1,4);
TASK_PP(16'h52F2,4);
TASK_PP(16'h52F3,4);
TASK_PP(16'h52F4,4);
TASK_PP(16'h52F5,4);
TASK_PP(16'h52F6,4);
TASK_PP(16'h52F7,4);
TASK_PP(16'h52F8,4);
TASK_PP(16'h52F9,4);
TASK_PP(16'h52FA,4);
TASK_PP(16'h52FB,4);
TASK_PP(16'h52FC,4);
TASK_PP(16'h52FD,4);
TASK_PP(16'h52FE,4);
TASK_PP(16'h52FF,4);
TASK_PP(16'h5300,4);
TASK_PP(16'h5301,4);
TASK_PP(16'h5302,4);
TASK_PP(16'h5303,4);
TASK_PP(16'h5304,4);
TASK_PP(16'h5305,4);
TASK_PP(16'h5306,4);
TASK_PP(16'h5307,4);
TASK_PP(16'h5308,4);
TASK_PP(16'h5309,4);
TASK_PP(16'h530A,4);
TASK_PP(16'h530B,4);
TASK_PP(16'h530C,4);
TASK_PP(16'h530D,4);
TASK_PP(16'h530E,4);
TASK_PP(16'h530F,4);
TASK_PP(16'h5310,4);
TASK_PP(16'h5311,4);
TASK_PP(16'h5312,4);
TASK_PP(16'h5313,4);
TASK_PP(16'h5314,4);
TASK_PP(16'h5315,4);
TASK_PP(16'h5316,4);
TASK_PP(16'h5317,4);
TASK_PP(16'h5318,4);
TASK_PP(16'h5319,4);
TASK_PP(16'h531A,4);
TASK_PP(16'h531B,4);
TASK_PP(16'h531C,4);
TASK_PP(16'h531D,4);
TASK_PP(16'h531E,4);
TASK_PP(16'h531F,4);
TASK_PP(16'h5320,4);
TASK_PP(16'h5321,4);
TASK_PP(16'h5322,4);
TASK_PP(16'h5323,4);
TASK_PP(16'h5324,4);
TASK_PP(16'h5325,4);
TASK_PP(16'h5326,4);
TASK_PP(16'h5327,4);
TASK_PP(16'h5328,4);
TASK_PP(16'h5329,4);
TASK_PP(16'h532A,4);
TASK_PP(16'h532B,4);
TASK_PP(16'h532C,4);
TASK_PP(16'h532D,4);
TASK_PP(16'h532E,4);
TASK_PP(16'h532F,4);
TASK_PP(16'h5330,4);
TASK_PP(16'h5331,4);
TASK_PP(16'h5332,4);
TASK_PP(16'h5333,4);
TASK_PP(16'h5334,4);
TASK_PP(16'h5335,4);
TASK_PP(16'h5336,4);
TASK_PP(16'h5337,4);
TASK_PP(16'h5338,4);
TASK_PP(16'h5339,4);
TASK_PP(16'h533A,4);
TASK_PP(16'h533B,4);
TASK_PP(16'h533C,4);
TASK_PP(16'h533D,4);
TASK_PP(16'h533E,4);
TASK_PP(16'h533F,4);
TASK_PP(16'h5340,4);
TASK_PP(16'h5341,4);
TASK_PP(16'h5342,4);
TASK_PP(16'h5343,4);
TASK_PP(16'h5344,4);
TASK_PP(16'h5345,4);
TASK_PP(16'h5346,4);
TASK_PP(16'h5347,4);
TASK_PP(16'h5348,4);
TASK_PP(16'h5349,4);
TASK_PP(16'h534A,4);
TASK_PP(16'h534B,4);
TASK_PP(16'h534C,4);
TASK_PP(16'h534D,4);
TASK_PP(16'h534E,4);
TASK_PP(16'h534F,4);
TASK_PP(16'h5350,4);
TASK_PP(16'h5351,4);
TASK_PP(16'h5352,4);
TASK_PP(16'h5353,4);
TASK_PP(16'h5354,4);
TASK_PP(16'h5355,4);
TASK_PP(16'h5356,4);
TASK_PP(16'h5357,4);
TASK_PP(16'h5358,4);
TASK_PP(16'h5359,4);
TASK_PP(16'h535A,4);
TASK_PP(16'h535B,4);
TASK_PP(16'h535C,4);
TASK_PP(16'h535D,4);
TASK_PP(16'h535E,4);
TASK_PP(16'h535F,4);
TASK_PP(16'h5360,4);
TASK_PP(16'h5361,4);
TASK_PP(16'h5362,4);
TASK_PP(16'h5363,4);
TASK_PP(16'h5364,4);
TASK_PP(16'h5365,4);
TASK_PP(16'h5366,4);
TASK_PP(16'h5367,4);
TASK_PP(16'h5368,4);
TASK_PP(16'h5369,4);
TASK_PP(16'h536A,4);
TASK_PP(16'h536B,4);
TASK_PP(16'h536C,4);
TASK_PP(16'h536D,4);
TASK_PP(16'h536E,4);
TASK_PP(16'h536F,4);
TASK_PP(16'h5370,4);
TASK_PP(16'h5371,4);
TASK_PP(16'h5372,4);
TASK_PP(16'h5373,4);
TASK_PP(16'h5374,4);
TASK_PP(16'h5375,4);
TASK_PP(16'h5376,4);
TASK_PP(16'h5377,4);
TASK_PP(16'h5378,4);
TASK_PP(16'h5379,4);
TASK_PP(16'h537A,4);
TASK_PP(16'h537B,4);
TASK_PP(16'h537C,4);
TASK_PP(16'h537D,4);
TASK_PP(16'h537E,4);
TASK_PP(16'h537F,4);
TASK_PP(16'h5380,4);
TASK_PP(16'h5381,4);
TASK_PP(16'h5382,4);
TASK_PP(16'h5383,4);
TASK_PP(16'h5384,4);
TASK_PP(16'h5385,4);
TASK_PP(16'h5386,4);
TASK_PP(16'h5387,4);
TASK_PP(16'h5388,4);
TASK_PP(16'h5389,4);
TASK_PP(16'h538A,4);
TASK_PP(16'h538B,4);
TASK_PP(16'h538C,4);
TASK_PP(16'h538D,4);
TASK_PP(16'h538E,4);
TASK_PP(16'h538F,4);
TASK_PP(16'h5390,4);
TASK_PP(16'h5391,4);
TASK_PP(16'h5392,4);
TASK_PP(16'h5393,4);
TASK_PP(16'h5394,4);
TASK_PP(16'h5395,4);
TASK_PP(16'h5396,4);
TASK_PP(16'h5397,4);
TASK_PP(16'h5398,4);
TASK_PP(16'h5399,4);
TASK_PP(16'h539A,4);
TASK_PP(16'h539B,4);
TASK_PP(16'h539C,4);
TASK_PP(16'h539D,4);
TASK_PP(16'h539E,4);
TASK_PP(16'h539F,4);
TASK_PP(16'h53A0,4);
TASK_PP(16'h53A1,4);
TASK_PP(16'h53A2,4);
TASK_PP(16'h53A3,4);
TASK_PP(16'h53A4,4);
TASK_PP(16'h53A5,4);
TASK_PP(16'h53A6,4);
TASK_PP(16'h53A7,4);
TASK_PP(16'h53A8,4);
TASK_PP(16'h53A9,4);
TASK_PP(16'h53AA,4);
TASK_PP(16'h53AB,4);
TASK_PP(16'h53AC,4);
TASK_PP(16'h53AD,4);
TASK_PP(16'h53AE,4);
TASK_PP(16'h53AF,4);
TASK_PP(16'h53B0,4);
TASK_PP(16'h53B1,4);
TASK_PP(16'h53B2,4);
TASK_PP(16'h53B3,4);
TASK_PP(16'h53B4,4);
TASK_PP(16'h53B5,4);
TASK_PP(16'h53B6,4);
TASK_PP(16'h53B7,4);
TASK_PP(16'h53B8,4);
TASK_PP(16'h53B9,4);
TASK_PP(16'h53BA,4);
TASK_PP(16'h53BB,4);
TASK_PP(16'h53BC,4);
TASK_PP(16'h53BD,4);
TASK_PP(16'h53BE,4);
TASK_PP(16'h53BF,4);
TASK_PP(16'h53C0,4);
TASK_PP(16'h53C1,4);
TASK_PP(16'h53C2,4);
TASK_PP(16'h53C3,4);
TASK_PP(16'h53C4,4);
TASK_PP(16'h53C5,4);
TASK_PP(16'h53C6,4);
TASK_PP(16'h53C7,4);
TASK_PP(16'h53C8,4);
TASK_PP(16'h53C9,4);
TASK_PP(16'h53CA,4);
TASK_PP(16'h53CB,4);
TASK_PP(16'h53CC,4);
TASK_PP(16'h53CD,4);
TASK_PP(16'h53CE,4);
TASK_PP(16'h53CF,4);
TASK_PP(16'h53D0,4);
TASK_PP(16'h53D1,4);
TASK_PP(16'h53D2,4);
TASK_PP(16'h53D3,4);
TASK_PP(16'h53D4,4);
TASK_PP(16'h53D5,4);
TASK_PP(16'h53D6,4);
TASK_PP(16'h53D7,4);
TASK_PP(16'h53D8,4);
TASK_PP(16'h53D9,4);
TASK_PP(16'h53DA,4);
TASK_PP(16'h53DB,4);
TASK_PP(16'h53DC,4);
TASK_PP(16'h53DD,4);
TASK_PP(16'h53DE,4);
TASK_PP(16'h53DF,4);
TASK_PP(16'h53E0,4);
TASK_PP(16'h53E1,4);
TASK_PP(16'h53E2,4);
TASK_PP(16'h53E3,4);
TASK_PP(16'h53E4,4);
TASK_PP(16'h53E5,4);
TASK_PP(16'h53E6,4);
TASK_PP(16'h53E7,4);
TASK_PP(16'h53E8,4);
TASK_PP(16'h53E9,4);
TASK_PP(16'h53EA,4);
TASK_PP(16'h53EB,4);
TASK_PP(16'h53EC,4);
TASK_PP(16'h53ED,4);
TASK_PP(16'h53EE,4);
TASK_PP(16'h53EF,4);
TASK_PP(16'h53F0,4);
TASK_PP(16'h53F1,4);
TASK_PP(16'h53F2,4);
TASK_PP(16'h53F3,4);
TASK_PP(16'h53F4,4);
TASK_PP(16'h53F5,4);
TASK_PP(16'h53F6,4);
TASK_PP(16'h53F7,4);
TASK_PP(16'h53F8,4);
TASK_PP(16'h53F9,4);
TASK_PP(16'h53FA,4);
TASK_PP(16'h53FB,4);
TASK_PP(16'h53FC,4);
TASK_PP(16'h53FD,4);
TASK_PP(16'h53FE,4);
TASK_PP(16'h53FF,4);
TASK_PP(16'h5400,4);
TASK_PP(16'h5401,4);
TASK_PP(16'h5402,4);
TASK_PP(16'h5403,4);
TASK_PP(16'h5404,4);
TASK_PP(16'h5405,4);
TASK_PP(16'h5406,4);
TASK_PP(16'h5407,4);
TASK_PP(16'h5408,4);
TASK_PP(16'h5409,4);
TASK_PP(16'h540A,4);
TASK_PP(16'h540B,4);
TASK_PP(16'h540C,4);
TASK_PP(16'h540D,4);
TASK_PP(16'h540E,4);
TASK_PP(16'h540F,4);
TASK_PP(16'h5410,4);
TASK_PP(16'h5411,4);
TASK_PP(16'h5412,4);
TASK_PP(16'h5413,4);
TASK_PP(16'h5414,4);
TASK_PP(16'h5415,4);
TASK_PP(16'h5416,4);
TASK_PP(16'h5417,4);
TASK_PP(16'h5418,4);
TASK_PP(16'h5419,4);
TASK_PP(16'h541A,4);
TASK_PP(16'h541B,4);
TASK_PP(16'h541C,4);
TASK_PP(16'h541D,4);
TASK_PP(16'h541E,4);
TASK_PP(16'h541F,4);
TASK_PP(16'h5420,4);
TASK_PP(16'h5421,4);
TASK_PP(16'h5422,4);
TASK_PP(16'h5423,4);
TASK_PP(16'h5424,4);
TASK_PP(16'h5425,4);
TASK_PP(16'h5426,4);
TASK_PP(16'h5427,4);
TASK_PP(16'h5428,4);
TASK_PP(16'h5429,4);
TASK_PP(16'h542A,4);
TASK_PP(16'h542B,4);
TASK_PP(16'h542C,4);
TASK_PP(16'h542D,4);
TASK_PP(16'h542E,4);
TASK_PP(16'h542F,4);
TASK_PP(16'h5430,4);
TASK_PP(16'h5431,4);
TASK_PP(16'h5432,4);
TASK_PP(16'h5433,4);
TASK_PP(16'h5434,4);
TASK_PP(16'h5435,4);
TASK_PP(16'h5436,4);
TASK_PP(16'h5437,4);
TASK_PP(16'h5438,4);
TASK_PP(16'h5439,4);
TASK_PP(16'h543A,4);
TASK_PP(16'h543B,4);
TASK_PP(16'h543C,4);
TASK_PP(16'h543D,4);
TASK_PP(16'h543E,4);
TASK_PP(16'h543F,4);
TASK_PP(16'h5440,4);
TASK_PP(16'h5441,4);
TASK_PP(16'h5442,4);
TASK_PP(16'h5443,4);
TASK_PP(16'h5444,4);
TASK_PP(16'h5445,4);
TASK_PP(16'h5446,4);
TASK_PP(16'h5447,4);
TASK_PP(16'h5448,4);
TASK_PP(16'h5449,4);
TASK_PP(16'h544A,4);
TASK_PP(16'h544B,4);
TASK_PP(16'h544C,4);
TASK_PP(16'h544D,4);
TASK_PP(16'h544E,4);
TASK_PP(16'h544F,4);
TASK_PP(16'h5450,4);
TASK_PP(16'h5451,4);
TASK_PP(16'h5452,4);
TASK_PP(16'h5453,4);
TASK_PP(16'h5454,4);
TASK_PP(16'h5455,4);
TASK_PP(16'h5456,4);
TASK_PP(16'h5457,4);
TASK_PP(16'h5458,4);
TASK_PP(16'h5459,4);
TASK_PP(16'h545A,4);
TASK_PP(16'h545B,4);
TASK_PP(16'h545C,4);
TASK_PP(16'h545D,4);
TASK_PP(16'h545E,4);
TASK_PP(16'h545F,4);
TASK_PP(16'h5460,4);
TASK_PP(16'h5461,4);
TASK_PP(16'h5462,4);
TASK_PP(16'h5463,4);
TASK_PP(16'h5464,4);
TASK_PP(16'h5465,4);
TASK_PP(16'h5466,4);
TASK_PP(16'h5467,4);
TASK_PP(16'h5468,4);
TASK_PP(16'h5469,4);
TASK_PP(16'h546A,4);
TASK_PP(16'h546B,4);
TASK_PP(16'h546C,4);
TASK_PP(16'h546D,4);
TASK_PP(16'h546E,4);
TASK_PP(16'h546F,4);
TASK_PP(16'h5470,4);
TASK_PP(16'h5471,4);
TASK_PP(16'h5472,4);
TASK_PP(16'h5473,4);
TASK_PP(16'h5474,4);
TASK_PP(16'h5475,4);
TASK_PP(16'h5476,4);
TASK_PP(16'h5477,4);
TASK_PP(16'h5478,4);
TASK_PP(16'h5479,4);
TASK_PP(16'h547A,4);
TASK_PP(16'h547B,4);
TASK_PP(16'h547C,4);
TASK_PP(16'h547D,4);
TASK_PP(16'h547E,4);
TASK_PP(16'h547F,4);
TASK_PP(16'h5480,4);
TASK_PP(16'h5481,4);
TASK_PP(16'h5482,4);
TASK_PP(16'h5483,4);
TASK_PP(16'h5484,4);
TASK_PP(16'h5485,4);
TASK_PP(16'h5486,4);
TASK_PP(16'h5487,4);
TASK_PP(16'h5488,4);
TASK_PP(16'h5489,4);
TASK_PP(16'h548A,4);
TASK_PP(16'h548B,4);
TASK_PP(16'h548C,4);
TASK_PP(16'h548D,4);
TASK_PP(16'h548E,4);
TASK_PP(16'h548F,4);
TASK_PP(16'h5490,4);
TASK_PP(16'h5491,4);
TASK_PP(16'h5492,4);
TASK_PP(16'h5493,4);
TASK_PP(16'h5494,4);
TASK_PP(16'h5495,4);
TASK_PP(16'h5496,4);
TASK_PP(16'h5497,4);
TASK_PP(16'h5498,4);
TASK_PP(16'h5499,4);
TASK_PP(16'h549A,4);
TASK_PP(16'h549B,4);
TASK_PP(16'h549C,4);
TASK_PP(16'h549D,4);
TASK_PP(16'h549E,4);
TASK_PP(16'h549F,4);
TASK_PP(16'h54A0,4);
TASK_PP(16'h54A1,4);
TASK_PP(16'h54A2,4);
TASK_PP(16'h54A3,4);
TASK_PP(16'h54A4,4);
TASK_PP(16'h54A5,4);
TASK_PP(16'h54A6,4);
TASK_PP(16'h54A7,4);
TASK_PP(16'h54A8,4);
TASK_PP(16'h54A9,4);
TASK_PP(16'h54AA,4);
TASK_PP(16'h54AB,4);
TASK_PP(16'h54AC,4);
TASK_PP(16'h54AD,4);
TASK_PP(16'h54AE,4);
TASK_PP(16'h54AF,4);
TASK_PP(16'h54B0,4);
TASK_PP(16'h54B1,4);
TASK_PP(16'h54B2,4);
TASK_PP(16'h54B3,4);
TASK_PP(16'h54B4,4);
TASK_PP(16'h54B5,4);
TASK_PP(16'h54B6,4);
TASK_PP(16'h54B7,4);
TASK_PP(16'h54B8,4);
TASK_PP(16'h54B9,4);
TASK_PP(16'h54BA,4);
TASK_PP(16'h54BB,4);
TASK_PP(16'h54BC,4);
TASK_PP(16'h54BD,4);
TASK_PP(16'h54BE,4);
TASK_PP(16'h54BF,4);
TASK_PP(16'h54C0,4);
TASK_PP(16'h54C1,4);
TASK_PP(16'h54C2,4);
TASK_PP(16'h54C3,4);
TASK_PP(16'h54C4,4);
TASK_PP(16'h54C5,4);
TASK_PP(16'h54C6,4);
TASK_PP(16'h54C7,4);
TASK_PP(16'h54C8,4);
TASK_PP(16'h54C9,4);
TASK_PP(16'h54CA,4);
TASK_PP(16'h54CB,4);
TASK_PP(16'h54CC,4);
TASK_PP(16'h54CD,4);
TASK_PP(16'h54CE,4);
TASK_PP(16'h54CF,4);
TASK_PP(16'h54D0,4);
TASK_PP(16'h54D1,4);
TASK_PP(16'h54D2,4);
TASK_PP(16'h54D3,4);
TASK_PP(16'h54D4,4);
TASK_PP(16'h54D5,4);
TASK_PP(16'h54D6,4);
TASK_PP(16'h54D7,4);
TASK_PP(16'h54D8,4);
TASK_PP(16'h54D9,4);
TASK_PP(16'h54DA,4);
TASK_PP(16'h54DB,4);
TASK_PP(16'h54DC,4);
TASK_PP(16'h54DD,4);
TASK_PP(16'h54DE,4);
TASK_PP(16'h54DF,4);
TASK_PP(16'h54E0,4);
TASK_PP(16'h54E1,4);
TASK_PP(16'h54E2,4);
TASK_PP(16'h54E3,4);
TASK_PP(16'h54E4,4);
TASK_PP(16'h54E5,4);
TASK_PP(16'h54E6,4);
TASK_PP(16'h54E7,4);
TASK_PP(16'h54E8,4);
TASK_PP(16'h54E9,4);
TASK_PP(16'h54EA,4);
TASK_PP(16'h54EB,4);
TASK_PP(16'h54EC,4);
TASK_PP(16'h54ED,4);
TASK_PP(16'h54EE,4);
TASK_PP(16'h54EF,4);
TASK_PP(16'h54F0,4);
TASK_PP(16'h54F1,4);
TASK_PP(16'h54F2,4);
TASK_PP(16'h54F3,4);
TASK_PP(16'h54F4,4);
TASK_PP(16'h54F5,4);
TASK_PP(16'h54F6,4);
TASK_PP(16'h54F7,4);
TASK_PP(16'h54F8,4);
TASK_PP(16'h54F9,4);
TASK_PP(16'h54FA,4);
TASK_PP(16'h54FB,4);
TASK_PP(16'h54FC,4);
TASK_PP(16'h54FD,4);
TASK_PP(16'h54FE,4);
TASK_PP(16'h54FF,4);
TASK_PP(16'h5500,4);
TASK_PP(16'h5501,4);
TASK_PP(16'h5502,4);
TASK_PP(16'h5503,4);
TASK_PP(16'h5504,4);
TASK_PP(16'h5505,4);
TASK_PP(16'h5506,4);
TASK_PP(16'h5507,4);
TASK_PP(16'h5508,4);
TASK_PP(16'h5509,4);
TASK_PP(16'h550A,4);
TASK_PP(16'h550B,4);
TASK_PP(16'h550C,4);
TASK_PP(16'h550D,4);
TASK_PP(16'h550E,4);
TASK_PP(16'h550F,4);
TASK_PP(16'h5510,4);
TASK_PP(16'h5511,4);
TASK_PP(16'h5512,4);
TASK_PP(16'h5513,4);
TASK_PP(16'h5514,4);
TASK_PP(16'h5515,4);
TASK_PP(16'h5516,4);
TASK_PP(16'h5517,4);
TASK_PP(16'h5518,4);
TASK_PP(16'h5519,4);
TASK_PP(16'h551A,4);
TASK_PP(16'h551B,4);
TASK_PP(16'h551C,4);
TASK_PP(16'h551D,4);
TASK_PP(16'h551E,4);
TASK_PP(16'h551F,4);
TASK_PP(16'h5520,4);
TASK_PP(16'h5521,4);
TASK_PP(16'h5522,4);
TASK_PP(16'h5523,4);
TASK_PP(16'h5524,4);
TASK_PP(16'h5525,4);
TASK_PP(16'h5526,4);
TASK_PP(16'h5527,4);
TASK_PP(16'h5528,4);
TASK_PP(16'h5529,4);
TASK_PP(16'h552A,4);
TASK_PP(16'h552B,4);
TASK_PP(16'h552C,4);
TASK_PP(16'h552D,4);
TASK_PP(16'h552E,4);
TASK_PP(16'h552F,4);
TASK_PP(16'h5530,4);
TASK_PP(16'h5531,4);
TASK_PP(16'h5532,4);
TASK_PP(16'h5533,4);
TASK_PP(16'h5534,4);
TASK_PP(16'h5535,4);
TASK_PP(16'h5536,4);
TASK_PP(16'h5537,4);
TASK_PP(16'h5538,4);
TASK_PP(16'h5539,4);
TASK_PP(16'h553A,4);
TASK_PP(16'h553B,4);
TASK_PP(16'h553C,4);
TASK_PP(16'h553D,4);
TASK_PP(16'h553E,4);
TASK_PP(16'h553F,4);
TASK_PP(16'h5540,4);
TASK_PP(16'h5541,4);
TASK_PP(16'h5542,4);
TASK_PP(16'h5543,4);
TASK_PP(16'h5544,4);
TASK_PP(16'h5545,4);
TASK_PP(16'h5546,4);
TASK_PP(16'h5547,4);
TASK_PP(16'h5548,4);
TASK_PP(16'h5549,4);
TASK_PP(16'h554A,4);
TASK_PP(16'h554B,4);
TASK_PP(16'h554C,4);
TASK_PP(16'h554D,4);
TASK_PP(16'h554E,4);
TASK_PP(16'h554F,4);
TASK_PP(16'h5550,4);
TASK_PP(16'h5551,4);
TASK_PP(16'h5552,4);
TASK_PP(16'h5553,4);
TASK_PP(16'h5554,4);
TASK_PP(16'h5555,4);
TASK_PP(16'h5556,4);
TASK_PP(16'h5557,4);
TASK_PP(16'h5558,4);
TASK_PP(16'h5559,4);
TASK_PP(16'h555A,4);
TASK_PP(16'h555B,4);
TASK_PP(16'h555C,4);
TASK_PP(16'h555D,4);
TASK_PP(16'h555E,4);
TASK_PP(16'h555F,4);
TASK_PP(16'h5560,4);
TASK_PP(16'h5561,4);
TASK_PP(16'h5562,4);
TASK_PP(16'h5563,4);
TASK_PP(16'h5564,4);
TASK_PP(16'h5565,4);
TASK_PP(16'h5566,4);
TASK_PP(16'h5567,4);
TASK_PP(16'h5568,4);
TASK_PP(16'h5569,4);
TASK_PP(16'h556A,4);
TASK_PP(16'h556B,4);
TASK_PP(16'h556C,4);
TASK_PP(16'h556D,4);
TASK_PP(16'h556E,4);
TASK_PP(16'h556F,4);
TASK_PP(16'h5570,4);
TASK_PP(16'h5571,4);
TASK_PP(16'h5572,4);
TASK_PP(16'h5573,4);
TASK_PP(16'h5574,4);
TASK_PP(16'h5575,4);
TASK_PP(16'h5576,4);
TASK_PP(16'h5577,4);
TASK_PP(16'h5578,4);
TASK_PP(16'h5579,4);
TASK_PP(16'h557A,4);
TASK_PP(16'h557B,4);
TASK_PP(16'h557C,4);
TASK_PP(16'h557D,4);
TASK_PP(16'h557E,4);
TASK_PP(16'h557F,4);
TASK_PP(16'h5580,4);
TASK_PP(16'h5581,4);
TASK_PP(16'h5582,4);
TASK_PP(16'h5583,4);
TASK_PP(16'h5584,4);
TASK_PP(16'h5585,4);
TASK_PP(16'h5586,4);
TASK_PP(16'h5587,4);
TASK_PP(16'h5588,4);
TASK_PP(16'h5589,4);
TASK_PP(16'h558A,4);
TASK_PP(16'h558B,4);
TASK_PP(16'h558C,4);
TASK_PP(16'h558D,4);
TASK_PP(16'h558E,4);
TASK_PP(16'h558F,4);
TASK_PP(16'h5590,4);
TASK_PP(16'h5591,4);
TASK_PP(16'h5592,4);
TASK_PP(16'h5593,4);
TASK_PP(16'h5594,4);
TASK_PP(16'h5595,4);
TASK_PP(16'h5596,4);
TASK_PP(16'h5597,4);
TASK_PP(16'h5598,4);
TASK_PP(16'h5599,4);
TASK_PP(16'h559A,4);
TASK_PP(16'h559B,4);
TASK_PP(16'h559C,4);
TASK_PP(16'h559D,4);
TASK_PP(16'h559E,4);
TASK_PP(16'h559F,4);
TASK_PP(16'h55A0,4);
TASK_PP(16'h55A1,4);
TASK_PP(16'h55A2,4);
TASK_PP(16'h55A3,4);
TASK_PP(16'h55A4,4);
TASK_PP(16'h55A5,4);
TASK_PP(16'h55A6,4);
TASK_PP(16'h55A7,4);
TASK_PP(16'h55A8,4);
TASK_PP(16'h55A9,4);
TASK_PP(16'h55AA,4);
TASK_PP(16'h55AB,4);
TASK_PP(16'h55AC,4);
TASK_PP(16'h55AD,4);
TASK_PP(16'h55AE,4);
TASK_PP(16'h55AF,4);
TASK_PP(16'h55B0,4);
TASK_PP(16'h55B1,4);
TASK_PP(16'h55B2,4);
TASK_PP(16'h55B3,4);
TASK_PP(16'h55B4,4);
TASK_PP(16'h55B5,4);
TASK_PP(16'h55B6,4);
TASK_PP(16'h55B7,4);
TASK_PP(16'h55B8,4);
TASK_PP(16'h55B9,4);
TASK_PP(16'h55BA,4);
TASK_PP(16'h55BB,4);
TASK_PP(16'h55BC,4);
TASK_PP(16'h55BD,4);
TASK_PP(16'h55BE,4);
TASK_PP(16'h55BF,4);
TASK_PP(16'h55C0,4);
TASK_PP(16'h55C1,4);
TASK_PP(16'h55C2,4);
TASK_PP(16'h55C3,4);
TASK_PP(16'h55C4,4);
TASK_PP(16'h55C5,4);
TASK_PP(16'h55C6,4);
TASK_PP(16'h55C7,4);
TASK_PP(16'h55C8,4);
TASK_PP(16'h55C9,4);
TASK_PP(16'h55CA,4);
TASK_PP(16'h55CB,4);
TASK_PP(16'h55CC,4);
TASK_PP(16'h55CD,4);
TASK_PP(16'h55CE,4);
TASK_PP(16'h55CF,4);
TASK_PP(16'h55D0,4);
TASK_PP(16'h55D1,4);
TASK_PP(16'h55D2,4);
TASK_PP(16'h55D3,4);
TASK_PP(16'h55D4,4);
TASK_PP(16'h55D5,4);
TASK_PP(16'h55D6,4);
TASK_PP(16'h55D7,4);
TASK_PP(16'h55D8,4);
TASK_PP(16'h55D9,4);
TASK_PP(16'h55DA,4);
TASK_PP(16'h55DB,4);
TASK_PP(16'h55DC,4);
TASK_PP(16'h55DD,4);
TASK_PP(16'h55DE,4);
TASK_PP(16'h55DF,4);
TASK_PP(16'h55E0,4);
TASK_PP(16'h55E1,4);
TASK_PP(16'h55E2,4);
TASK_PP(16'h55E3,4);
TASK_PP(16'h55E4,4);
TASK_PP(16'h55E5,4);
TASK_PP(16'h55E6,4);
TASK_PP(16'h55E7,4);
TASK_PP(16'h55E8,4);
TASK_PP(16'h55E9,4);
TASK_PP(16'h55EA,4);
TASK_PP(16'h55EB,4);
TASK_PP(16'h55EC,4);
TASK_PP(16'h55ED,4);
TASK_PP(16'h55EE,4);
TASK_PP(16'h55EF,4);
TASK_PP(16'h55F0,4);
TASK_PP(16'h55F1,4);
TASK_PP(16'h55F2,4);
TASK_PP(16'h55F3,4);
TASK_PP(16'h55F4,4);
TASK_PP(16'h55F5,4);
TASK_PP(16'h55F6,4);
TASK_PP(16'h55F7,4);
TASK_PP(16'h55F8,4);
TASK_PP(16'h55F9,4);
TASK_PP(16'h55FA,4);
TASK_PP(16'h55FB,4);
TASK_PP(16'h55FC,4);
TASK_PP(16'h55FD,4);
TASK_PP(16'h55FE,4);
TASK_PP(16'h55FF,4);
TASK_PP(16'h5600,4);
TASK_PP(16'h5601,4);
TASK_PP(16'h5602,4);
TASK_PP(16'h5603,4);
TASK_PP(16'h5604,4);
TASK_PP(16'h5605,4);
TASK_PP(16'h5606,4);
TASK_PP(16'h5607,4);
TASK_PP(16'h5608,4);
TASK_PP(16'h5609,4);
TASK_PP(16'h560A,4);
TASK_PP(16'h560B,4);
TASK_PP(16'h560C,4);
TASK_PP(16'h560D,4);
TASK_PP(16'h560E,4);
TASK_PP(16'h560F,4);
TASK_PP(16'h5610,4);
TASK_PP(16'h5611,4);
TASK_PP(16'h5612,4);
TASK_PP(16'h5613,4);
TASK_PP(16'h5614,4);
TASK_PP(16'h5615,4);
TASK_PP(16'h5616,4);
TASK_PP(16'h5617,4);
TASK_PP(16'h5618,4);
TASK_PP(16'h5619,4);
TASK_PP(16'h561A,4);
TASK_PP(16'h561B,4);
TASK_PP(16'h561C,4);
TASK_PP(16'h561D,4);
TASK_PP(16'h561E,4);
TASK_PP(16'h561F,4);
TASK_PP(16'h5620,4);
TASK_PP(16'h5621,4);
TASK_PP(16'h5622,4);
TASK_PP(16'h5623,4);
TASK_PP(16'h5624,4);
TASK_PP(16'h5625,4);
TASK_PP(16'h5626,4);
TASK_PP(16'h5627,4);
TASK_PP(16'h5628,4);
TASK_PP(16'h5629,4);
TASK_PP(16'h562A,4);
TASK_PP(16'h562B,4);
TASK_PP(16'h562C,4);
TASK_PP(16'h562D,4);
TASK_PP(16'h562E,4);
TASK_PP(16'h562F,4);
TASK_PP(16'h5630,4);
TASK_PP(16'h5631,4);
TASK_PP(16'h5632,4);
TASK_PP(16'h5633,4);
TASK_PP(16'h5634,4);
TASK_PP(16'h5635,4);
TASK_PP(16'h5636,4);
TASK_PP(16'h5637,4);
TASK_PP(16'h5638,4);
TASK_PP(16'h5639,4);
TASK_PP(16'h563A,4);
TASK_PP(16'h563B,4);
TASK_PP(16'h563C,4);
TASK_PP(16'h563D,4);
TASK_PP(16'h563E,4);
TASK_PP(16'h563F,4);
TASK_PP(16'h5640,4);
TASK_PP(16'h5641,4);
TASK_PP(16'h5642,4);
TASK_PP(16'h5643,4);
TASK_PP(16'h5644,4);
TASK_PP(16'h5645,4);
TASK_PP(16'h5646,4);
TASK_PP(16'h5647,4);
TASK_PP(16'h5648,4);
TASK_PP(16'h5649,4);
TASK_PP(16'h564A,4);
TASK_PP(16'h564B,4);
TASK_PP(16'h564C,4);
TASK_PP(16'h564D,4);
TASK_PP(16'h564E,4);
TASK_PP(16'h564F,4);
TASK_PP(16'h5650,4);
TASK_PP(16'h5651,4);
TASK_PP(16'h5652,4);
TASK_PP(16'h5653,4);
TASK_PP(16'h5654,4);
TASK_PP(16'h5655,4);
TASK_PP(16'h5656,4);
TASK_PP(16'h5657,4);
TASK_PP(16'h5658,4);
TASK_PP(16'h5659,4);
TASK_PP(16'h565A,4);
TASK_PP(16'h565B,4);
TASK_PP(16'h565C,4);
TASK_PP(16'h565D,4);
TASK_PP(16'h565E,4);
TASK_PP(16'h565F,4);
TASK_PP(16'h5660,4);
TASK_PP(16'h5661,4);
TASK_PP(16'h5662,4);
TASK_PP(16'h5663,4);
TASK_PP(16'h5664,4);
TASK_PP(16'h5665,4);
TASK_PP(16'h5666,4);
TASK_PP(16'h5667,4);
TASK_PP(16'h5668,4);
TASK_PP(16'h5669,4);
TASK_PP(16'h566A,4);
TASK_PP(16'h566B,4);
TASK_PP(16'h566C,4);
TASK_PP(16'h566D,4);
TASK_PP(16'h566E,4);
TASK_PP(16'h566F,4);
TASK_PP(16'h5670,4);
TASK_PP(16'h5671,4);
TASK_PP(16'h5672,4);
TASK_PP(16'h5673,4);
TASK_PP(16'h5674,4);
TASK_PP(16'h5675,4);
TASK_PP(16'h5676,4);
TASK_PP(16'h5677,4);
TASK_PP(16'h5678,4);
TASK_PP(16'h5679,4);
TASK_PP(16'h567A,4);
TASK_PP(16'h567B,4);
TASK_PP(16'h567C,4);
TASK_PP(16'h567D,4);
TASK_PP(16'h567E,4);
TASK_PP(16'h567F,4);
TASK_PP(16'h5680,4);
TASK_PP(16'h5681,4);
TASK_PP(16'h5682,4);
TASK_PP(16'h5683,4);
TASK_PP(16'h5684,4);
TASK_PP(16'h5685,4);
TASK_PP(16'h5686,4);
TASK_PP(16'h5687,4);
TASK_PP(16'h5688,4);
TASK_PP(16'h5689,4);
TASK_PP(16'h568A,4);
TASK_PP(16'h568B,4);
TASK_PP(16'h568C,4);
TASK_PP(16'h568D,4);
TASK_PP(16'h568E,4);
TASK_PP(16'h568F,4);
TASK_PP(16'h5690,4);
TASK_PP(16'h5691,4);
TASK_PP(16'h5692,4);
TASK_PP(16'h5693,4);
TASK_PP(16'h5694,4);
TASK_PP(16'h5695,4);
TASK_PP(16'h5696,4);
TASK_PP(16'h5697,4);
TASK_PP(16'h5698,4);
TASK_PP(16'h5699,4);
TASK_PP(16'h569A,4);
TASK_PP(16'h569B,4);
TASK_PP(16'h569C,4);
TASK_PP(16'h569D,4);
TASK_PP(16'h569E,4);
TASK_PP(16'h569F,4);
TASK_PP(16'h56A0,4);
TASK_PP(16'h56A1,4);
TASK_PP(16'h56A2,4);
TASK_PP(16'h56A3,4);
TASK_PP(16'h56A4,4);
TASK_PP(16'h56A5,4);
TASK_PP(16'h56A6,4);
TASK_PP(16'h56A7,4);
TASK_PP(16'h56A8,4);
TASK_PP(16'h56A9,4);
TASK_PP(16'h56AA,4);
TASK_PP(16'h56AB,4);
TASK_PP(16'h56AC,4);
TASK_PP(16'h56AD,4);
TASK_PP(16'h56AE,4);
TASK_PP(16'h56AF,4);
TASK_PP(16'h56B0,4);
TASK_PP(16'h56B1,4);
TASK_PP(16'h56B2,4);
TASK_PP(16'h56B3,4);
TASK_PP(16'h56B4,4);
TASK_PP(16'h56B5,4);
TASK_PP(16'h56B6,4);
TASK_PP(16'h56B7,4);
TASK_PP(16'h56B8,4);
TASK_PP(16'h56B9,4);
TASK_PP(16'h56BA,4);
TASK_PP(16'h56BB,4);
TASK_PP(16'h56BC,4);
TASK_PP(16'h56BD,4);
TASK_PP(16'h56BE,4);
TASK_PP(16'h56BF,4);
TASK_PP(16'h56C0,4);
TASK_PP(16'h56C1,4);
TASK_PP(16'h56C2,4);
TASK_PP(16'h56C3,4);
TASK_PP(16'h56C4,4);
TASK_PP(16'h56C5,4);
TASK_PP(16'h56C6,4);
TASK_PP(16'h56C7,4);
TASK_PP(16'h56C8,4);
TASK_PP(16'h56C9,4);
TASK_PP(16'h56CA,4);
TASK_PP(16'h56CB,4);
TASK_PP(16'h56CC,4);
TASK_PP(16'h56CD,4);
TASK_PP(16'h56CE,4);
TASK_PP(16'h56CF,4);
TASK_PP(16'h56D0,4);
TASK_PP(16'h56D1,4);
TASK_PP(16'h56D2,4);
TASK_PP(16'h56D3,4);
TASK_PP(16'h56D4,4);
TASK_PP(16'h56D5,4);
TASK_PP(16'h56D6,4);
TASK_PP(16'h56D7,4);
TASK_PP(16'h56D8,4);
TASK_PP(16'h56D9,4);
TASK_PP(16'h56DA,4);
TASK_PP(16'h56DB,4);
TASK_PP(16'h56DC,4);
TASK_PP(16'h56DD,4);
TASK_PP(16'h56DE,4);
TASK_PP(16'h56DF,4);
TASK_PP(16'h56E0,4);
TASK_PP(16'h56E1,4);
TASK_PP(16'h56E2,4);
TASK_PP(16'h56E3,4);
TASK_PP(16'h56E4,4);
TASK_PP(16'h56E5,4);
TASK_PP(16'h56E6,4);
TASK_PP(16'h56E7,4);
TASK_PP(16'h56E8,4);
TASK_PP(16'h56E9,4);
TASK_PP(16'h56EA,4);
TASK_PP(16'h56EB,4);
TASK_PP(16'h56EC,4);
TASK_PP(16'h56ED,4);
TASK_PP(16'h56EE,4);
TASK_PP(16'h56EF,4);
TASK_PP(16'h56F0,4);
TASK_PP(16'h56F1,4);
TASK_PP(16'h56F2,4);
TASK_PP(16'h56F3,4);
TASK_PP(16'h56F4,4);
TASK_PP(16'h56F5,4);
TASK_PP(16'h56F6,4);
TASK_PP(16'h56F7,4);
TASK_PP(16'h56F8,4);
TASK_PP(16'h56F9,4);
TASK_PP(16'h56FA,4);
TASK_PP(16'h56FB,4);
TASK_PP(16'h56FC,4);
TASK_PP(16'h56FD,4);
TASK_PP(16'h56FE,4);
TASK_PP(16'h56FF,4);
TASK_PP(16'h5700,4);
TASK_PP(16'h5701,4);
TASK_PP(16'h5702,4);
TASK_PP(16'h5703,4);
TASK_PP(16'h5704,4);
TASK_PP(16'h5705,4);
TASK_PP(16'h5706,4);
TASK_PP(16'h5707,4);
TASK_PP(16'h5708,4);
TASK_PP(16'h5709,4);
TASK_PP(16'h570A,4);
TASK_PP(16'h570B,4);
TASK_PP(16'h570C,4);
TASK_PP(16'h570D,4);
TASK_PP(16'h570E,4);
TASK_PP(16'h570F,4);
TASK_PP(16'h5710,4);
TASK_PP(16'h5711,4);
TASK_PP(16'h5712,4);
TASK_PP(16'h5713,4);
TASK_PP(16'h5714,4);
TASK_PP(16'h5715,4);
TASK_PP(16'h5716,4);
TASK_PP(16'h5717,4);
TASK_PP(16'h5718,4);
TASK_PP(16'h5719,4);
TASK_PP(16'h571A,4);
TASK_PP(16'h571B,4);
TASK_PP(16'h571C,4);
TASK_PP(16'h571D,4);
TASK_PP(16'h571E,4);
TASK_PP(16'h571F,4);
TASK_PP(16'h5720,4);
TASK_PP(16'h5721,4);
TASK_PP(16'h5722,4);
TASK_PP(16'h5723,4);
TASK_PP(16'h5724,4);
TASK_PP(16'h5725,4);
TASK_PP(16'h5726,4);
TASK_PP(16'h5727,4);
TASK_PP(16'h5728,4);
TASK_PP(16'h5729,4);
TASK_PP(16'h572A,4);
TASK_PP(16'h572B,4);
TASK_PP(16'h572C,4);
TASK_PP(16'h572D,4);
TASK_PP(16'h572E,4);
TASK_PP(16'h572F,4);
TASK_PP(16'h5730,4);
TASK_PP(16'h5731,4);
TASK_PP(16'h5732,4);
TASK_PP(16'h5733,4);
TASK_PP(16'h5734,4);
TASK_PP(16'h5735,4);
TASK_PP(16'h5736,4);
TASK_PP(16'h5737,4);
TASK_PP(16'h5738,4);
TASK_PP(16'h5739,4);
TASK_PP(16'h573A,4);
TASK_PP(16'h573B,4);
TASK_PP(16'h573C,4);
TASK_PP(16'h573D,4);
TASK_PP(16'h573E,4);
TASK_PP(16'h573F,4);
TASK_PP(16'h5740,4);
TASK_PP(16'h5741,4);
TASK_PP(16'h5742,4);
TASK_PP(16'h5743,4);
TASK_PP(16'h5744,4);
TASK_PP(16'h5745,4);
TASK_PP(16'h5746,4);
TASK_PP(16'h5747,4);
TASK_PP(16'h5748,4);
TASK_PP(16'h5749,4);
TASK_PP(16'h574A,4);
TASK_PP(16'h574B,4);
TASK_PP(16'h574C,4);
TASK_PP(16'h574D,4);
TASK_PP(16'h574E,4);
TASK_PP(16'h574F,4);
TASK_PP(16'h5750,4);
TASK_PP(16'h5751,4);
TASK_PP(16'h5752,4);
TASK_PP(16'h5753,4);
TASK_PP(16'h5754,4);
TASK_PP(16'h5755,4);
TASK_PP(16'h5756,4);
TASK_PP(16'h5757,4);
TASK_PP(16'h5758,4);
TASK_PP(16'h5759,4);
TASK_PP(16'h575A,4);
TASK_PP(16'h575B,4);
TASK_PP(16'h575C,4);
TASK_PP(16'h575D,4);
TASK_PP(16'h575E,4);
TASK_PP(16'h575F,4);
TASK_PP(16'h5760,4);
TASK_PP(16'h5761,4);
TASK_PP(16'h5762,4);
TASK_PP(16'h5763,4);
TASK_PP(16'h5764,4);
TASK_PP(16'h5765,4);
TASK_PP(16'h5766,4);
TASK_PP(16'h5767,4);
TASK_PP(16'h5768,4);
TASK_PP(16'h5769,4);
TASK_PP(16'h576A,4);
TASK_PP(16'h576B,4);
TASK_PP(16'h576C,4);
TASK_PP(16'h576D,4);
TASK_PP(16'h576E,4);
TASK_PP(16'h576F,4);
TASK_PP(16'h5770,4);
TASK_PP(16'h5771,4);
TASK_PP(16'h5772,4);
TASK_PP(16'h5773,4);
TASK_PP(16'h5774,4);
TASK_PP(16'h5775,4);
TASK_PP(16'h5776,4);
TASK_PP(16'h5777,4);
TASK_PP(16'h5778,4);
TASK_PP(16'h5779,4);
TASK_PP(16'h577A,4);
TASK_PP(16'h577B,4);
TASK_PP(16'h577C,4);
TASK_PP(16'h577D,4);
TASK_PP(16'h577E,4);
TASK_PP(16'h577F,4);
TASK_PP(16'h5780,4);
TASK_PP(16'h5781,4);
TASK_PP(16'h5782,4);
TASK_PP(16'h5783,4);
TASK_PP(16'h5784,4);
TASK_PP(16'h5785,4);
TASK_PP(16'h5786,4);
TASK_PP(16'h5787,4);
TASK_PP(16'h5788,4);
TASK_PP(16'h5789,4);
TASK_PP(16'h578A,4);
TASK_PP(16'h578B,4);
TASK_PP(16'h578C,4);
TASK_PP(16'h578D,4);
TASK_PP(16'h578E,4);
TASK_PP(16'h578F,4);
TASK_PP(16'h5790,4);
TASK_PP(16'h5791,4);
TASK_PP(16'h5792,4);
TASK_PP(16'h5793,4);
TASK_PP(16'h5794,4);
TASK_PP(16'h5795,4);
TASK_PP(16'h5796,4);
TASK_PP(16'h5797,4);
TASK_PP(16'h5798,4);
TASK_PP(16'h5799,4);
TASK_PP(16'h579A,4);
TASK_PP(16'h579B,4);
TASK_PP(16'h579C,4);
TASK_PP(16'h579D,4);
TASK_PP(16'h579E,4);
TASK_PP(16'h579F,4);
TASK_PP(16'h57A0,4);
TASK_PP(16'h57A1,4);
TASK_PP(16'h57A2,4);
TASK_PP(16'h57A3,4);
TASK_PP(16'h57A4,4);
TASK_PP(16'h57A5,4);
TASK_PP(16'h57A6,4);
TASK_PP(16'h57A7,4);
TASK_PP(16'h57A8,4);
TASK_PP(16'h57A9,4);
TASK_PP(16'h57AA,4);
TASK_PP(16'h57AB,4);
TASK_PP(16'h57AC,4);
TASK_PP(16'h57AD,4);
TASK_PP(16'h57AE,4);
TASK_PP(16'h57AF,4);
TASK_PP(16'h57B0,4);
TASK_PP(16'h57B1,4);
TASK_PP(16'h57B2,4);
TASK_PP(16'h57B3,4);
TASK_PP(16'h57B4,4);
TASK_PP(16'h57B5,4);
TASK_PP(16'h57B6,4);
TASK_PP(16'h57B7,4);
TASK_PP(16'h57B8,4);
TASK_PP(16'h57B9,4);
TASK_PP(16'h57BA,4);
TASK_PP(16'h57BB,4);
TASK_PP(16'h57BC,4);
TASK_PP(16'h57BD,4);
TASK_PP(16'h57BE,4);
TASK_PP(16'h57BF,4);
TASK_PP(16'h57C0,4);
TASK_PP(16'h57C1,4);
TASK_PP(16'h57C2,4);
TASK_PP(16'h57C3,4);
TASK_PP(16'h57C4,4);
TASK_PP(16'h57C5,4);
TASK_PP(16'h57C6,4);
TASK_PP(16'h57C7,4);
TASK_PP(16'h57C8,4);
TASK_PP(16'h57C9,4);
TASK_PP(16'h57CA,4);
TASK_PP(16'h57CB,4);
TASK_PP(16'h57CC,4);
TASK_PP(16'h57CD,4);
TASK_PP(16'h57CE,4);
TASK_PP(16'h57CF,4);
TASK_PP(16'h57D0,4);
TASK_PP(16'h57D1,4);
TASK_PP(16'h57D2,4);
TASK_PP(16'h57D3,4);
TASK_PP(16'h57D4,4);
TASK_PP(16'h57D5,4);
TASK_PP(16'h57D6,4);
TASK_PP(16'h57D7,4);
TASK_PP(16'h57D8,4);
TASK_PP(16'h57D9,4);
TASK_PP(16'h57DA,4);
TASK_PP(16'h57DB,4);
TASK_PP(16'h57DC,4);
TASK_PP(16'h57DD,4);
TASK_PP(16'h57DE,4);
TASK_PP(16'h57DF,4);
TASK_PP(16'h57E0,4);
TASK_PP(16'h57E1,4);
TASK_PP(16'h57E2,4);
TASK_PP(16'h57E3,4);
TASK_PP(16'h57E4,4);
TASK_PP(16'h57E5,4);
TASK_PP(16'h57E6,4);
TASK_PP(16'h57E7,4);
TASK_PP(16'h57E8,4);
TASK_PP(16'h57E9,4);
TASK_PP(16'h57EA,4);
TASK_PP(16'h57EB,4);
TASK_PP(16'h57EC,4);
TASK_PP(16'h57ED,4);
TASK_PP(16'h57EE,4);
TASK_PP(16'h57EF,4);
TASK_PP(16'h57F0,4);
TASK_PP(16'h57F1,4);
TASK_PP(16'h57F2,4);
TASK_PP(16'h57F3,4);
TASK_PP(16'h57F4,4);
TASK_PP(16'h57F5,4);
TASK_PP(16'h57F6,4);
TASK_PP(16'h57F7,4);
TASK_PP(16'h57F8,4);
TASK_PP(16'h57F9,4);
TASK_PP(16'h57FA,4);
TASK_PP(16'h57FB,4);
TASK_PP(16'h57FC,4);
TASK_PP(16'h57FD,4);
TASK_PP(16'h57FE,4);
TASK_PP(16'h57FF,4);
TASK_PP(16'h5800,4);
TASK_PP(16'h5801,4);
TASK_PP(16'h5802,4);
TASK_PP(16'h5803,4);
TASK_PP(16'h5804,4);
TASK_PP(16'h5805,4);
TASK_PP(16'h5806,4);
TASK_PP(16'h5807,4);
TASK_PP(16'h5808,4);
TASK_PP(16'h5809,4);
TASK_PP(16'h580A,4);
TASK_PP(16'h580B,4);
TASK_PP(16'h580C,4);
TASK_PP(16'h580D,4);
TASK_PP(16'h580E,4);
TASK_PP(16'h580F,4);
TASK_PP(16'h5810,4);
TASK_PP(16'h5811,4);
TASK_PP(16'h5812,4);
TASK_PP(16'h5813,4);
TASK_PP(16'h5814,4);
TASK_PP(16'h5815,4);
TASK_PP(16'h5816,4);
TASK_PP(16'h5817,4);
TASK_PP(16'h5818,4);
TASK_PP(16'h5819,4);
TASK_PP(16'h581A,4);
TASK_PP(16'h581B,4);
TASK_PP(16'h581C,4);
TASK_PP(16'h581D,4);
TASK_PP(16'h581E,4);
TASK_PP(16'h581F,4);
TASK_PP(16'h5820,4);
TASK_PP(16'h5821,4);
TASK_PP(16'h5822,4);
TASK_PP(16'h5823,4);
TASK_PP(16'h5824,4);
TASK_PP(16'h5825,4);
TASK_PP(16'h5826,4);
TASK_PP(16'h5827,4);
TASK_PP(16'h5828,4);
TASK_PP(16'h5829,4);
TASK_PP(16'h582A,4);
TASK_PP(16'h582B,4);
TASK_PP(16'h582C,4);
TASK_PP(16'h582D,4);
TASK_PP(16'h582E,4);
TASK_PP(16'h582F,4);
TASK_PP(16'h5830,4);
TASK_PP(16'h5831,4);
TASK_PP(16'h5832,4);
TASK_PP(16'h5833,4);
TASK_PP(16'h5834,4);
TASK_PP(16'h5835,4);
TASK_PP(16'h5836,4);
TASK_PP(16'h5837,4);
TASK_PP(16'h5838,4);
TASK_PP(16'h5839,4);
TASK_PP(16'h583A,4);
TASK_PP(16'h583B,4);
TASK_PP(16'h583C,4);
TASK_PP(16'h583D,4);
TASK_PP(16'h583E,4);
TASK_PP(16'h583F,4);
TASK_PP(16'h5840,4);
TASK_PP(16'h5841,4);
TASK_PP(16'h5842,4);
TASK_PP(16'h5843,4);
TASK_PP(16'h5844,4);
TASK_PP(16'h5845,4);
TASK_PP(16'h5846,4);
TASK_PP(16'h5847,4);
TASK_PP(16'h5848,4);
TASK_PP(16'h5849,4);
TASK_PP(16'h584A,4);
TASK_PP(16'h584B,4);
TASK_PP(16'h584C,4);
TASK_PP(16'h584D,4);
TASK_PP(16'h584E,4);
TASK_PP(16'h584F,4);
TASK_PP(16'h5850,4);
TASK_PP(16'h5851,4);
TASK_PP(16'h5852,4);
TASK_PP(16'h5853,4);
TASK_PP(16'h5854,4);
TASK_PP(16'h5855,4);
TASK_PP(16'h5856,4);
TASK_PP(16'h5857,4);
TASK_PP(16'h5858,4);
TASK_PP(16'h5859,4);
TASK_PP(16'h585A,4);
TASK_PP(16'h585B,4);
TASK_PP(16'h585C,4);
TASK_PP(16'h585D,4);
TASK_PP(16'h585E,4);
TASK_PP(16'h585F,4);
TASK_PP(16'h5860,4);
TASK_PP(16'h5861,4);
TASK_PP(16'h5862,4);
TASK_PP(16'h5863,4);
TASK_PP(16'h5864,4);
TASK_PP(16'h5865,4);
TASK_PP(16'h5866,4);
TASK_PP(16'h5867,4);
TASK_PP(16'h5868,4);
TASK_PP(16'h5869,4);
TASK_PP(16'h586A,4);
TASK_PP(16'h586B,4);
TASK_PP(16'h586C,4);
TASK_PP(16'h586D,4);
TASK_PP(16'h586E,4);
TASK_PP(16'h586F,4);
TASK_PP(16'h5870,4);
TASK_PP(16'h5871,4);
TASK_PP(16'h5872,4);
TASK_PP(16'h5873,4);
TASK_PP(16'h5874,4);
TASK_PP(16'h5875,4);
TASK_PP(16'h5876,4);
TASK_PP(16'h5877,4);
TASK_PP(16'h5878,4);
TASK_PP(16'h5879,4);
TASK_PP(16'h587A,4);
TASK_PP(16'h587B,4);
TASK_PP(16'h587C,4);
TASK_PP(16'h587D,4);
TASK_PP(16'h587E,4);
TASK_PP(16'h587F,4);
TASK_PP(16'h5880,4);
TASK_PP(16'h5881,4);
TASK_PP(16'h5882,4);
TASK_PP(16'h5883,4);
TASK_PP(16'h5884,4);
TASK_PP(16'h5885,4);
TASK_PP(16'h5886,4);
TASK_PP(16'h5887,4);
TASK_PP(16'h5888,4);
TASK_PP(16'h5889,4);
TASK_PP(16'h588A,4);
TASK_PP(16'h588B,4);
TASK_PP(16'h588C,4);
TASK_PP(16'h588D,4);
TASK_PP(16'h588E,4);
TASK_PP(16'h588F,4);
TASK_PP(16'h5890,4);
TASK_PP(16'h5891,4);
TASK_PP(16'h5892,4);
TASK_PP(16'h5893,4);
TASK_PP(16'h5894,4);
TASK_PP(16'h5895,4);
TASK_PP(16'h5896,4);
TASK_PP(16'h5897,4);
TASK_PP(16'h5898,4);
TASK_PP(16'h5899,4);
TASK_PP(16'h589A,4);
TASK_PP(16'h589B,4);
TASK_PP(16'h589C,4);
TASK_PP(16'h589D,4);
TASK_PP(16'h589E,4);
TASK_PP(16'h589F,4);
TASK_PP(16'h58A0,4);
TASK_PP(16'h58A1,4);
TASK_PP(16'h58A2,4);
TASK_PP(16'h58A3,4);
TASK_PP(16'h58A4,4);
TASK_PP(16'h58A5,4);
TASK_PP(16'h58A6,4);
TASK_PP(16'h58A7,4);
TASK_PP(16'h58A8,4);
TASK_PP(16'h58A9,4);
TASK_PP(16'h58AA,4);
TASK_PP(16'h58AB,4);
TASK_PP(16'h58AC,4);
TASK_PP(16'h58AD,4);
TASK_PP(16'h58AE,4);
TASK_PP(16'h58AF,4);
TASK_PP(16'h58B0,4);
TASK_PP(16'h58B1,4);
TASK_PP(16'h58B2,4);
TASK_PP(16'h58B3,4);
TASK_PP(16'h58B4,4);
TASK_PP(16'h58B5,4);
TASK_PP(16'h58B6,4);
TASK_PP(16'h58B7,4);
TASK_PP(16'h58B8,4);
TASK_PP(16'h58B9,4);
TASK_PP(16'h58BA,4);
TASK_PP(16'h58BB,4);
TASK_PP(16'h58BC,4);
TASK_PP(16'h58BD,4);
TASK_PP(16'h58BE,4);
TASK_PP(16'h58BF,4);
TASK_PP(16'h58C0,4);
TASK_PP(16'h58C1,4);
TASK_PP(16'h58C2,4);
TASK_PP(16'h58C3,4);
TASK_PP(16'h58C4,4);
TASK_PP(16'h58C5,4);
TASK_PP(16'h58C6,4);
TASK_PP(16'h58C7,4);
TASK_PP(16'h58C8,4);
TASK_PP(16'h58C9,4);
TASK_PP(16'h58CA,4);
TASK_PP(16'h58CB,4);
TASK_PP(16'h58CC,4);
TASK_PP(16'h58CD,4);
TASK_PP(16'h58CE,4);
TASK_PP(16'h58CF,4);
TASK_PP(16'h58D0,4);
TASK_PP(16'h58D1,4);
TASK_PP(16'h58D2,4);
TASK_PP(16'h58D3,4);
TASK_PP(16'h58D4,4);
TASK_PP(16'h58D5,4);
TASK_PP(16'h58D6,4);
TASK_PP(16'h58D7,4);
TASK_PP(16'h58D8,4);
TASK_PP(16'h58D9,4);
TASK_PP(16'h58DA,4);
TASK_PP(16'h58DB,4);
TASK_PP(16'h58DC,4);
TASK_PP(16'h58DD,4);
TASK_PP(16'h58DE,4);
TASK_PP(16'h58DF,4);
TASK_PP(16'h58E0,4);
TASK_PP(16'h58E1,4);
TASK_PP(16'h58E2,4);
TASK_PP(16'h58E3,4);
TASK_PP(16'h58E4,4);
TASK_PP(16'h58E5,4);
TASK_PP(16'h58E6,4);
TASK_PP(16'h58E7,4);
TASK_PP(16'h58E8,4);
TASK_PP(16'h58E9,4);
TASK_PP(16'h58EA,4);
TASK_PP(16'h58EB,4);
TASK_PP(16'h58EC,4);
TASK_PP(16'h58ED,4);
TASK_PP(16'h58EE,4);
TASK_PP(16'h58EF,4);
TASK_PP(16'h58F0,4);
TASK_PP(16'h58F1,4);
TASK_PP(16'h58F2,4);
TASK_PP(16'h58F3,4);
TASK_PP(16'h58F4,4);
TASK_PP(16'h58F5,4);
TASK_PP(16'h58F6,4);
TASK_PP(16'h58F7,4);
TASK_PP(16'h58F8,4);
TASK_PP(16'h58F9,4);
TASK_PP(16'h58FA,4);
TASK_PP(16'h58FB,4);
TASK_PP(16'h58FC,4);
TASK_PP(16'h58FD,4);
TASK_PP(16'h58FE,4);
TASK_PP(16'h58FF,4);
TASK_PP(16'h5900,4);
TASK_PP(16'h5901,4);
TASK_PP(16'h5902,4);
TASK_PP(16'h5903,4);
TASK_PP(16'h5904,4);
TASK_PP(16'h5905,4);
TASK_PP(16'h5906,4);
TASK_PP(16'h5907,4);
TASK_PP(16'h5908,4);
TASK_PP(16'h5909,4);
TASK_PP(16'h590A,4);
TASK_PP(16'h590B,4);
TASK_PP(16'h590C,4);
TASK_PP(16'h590D,4);
TASK_PP(16'h590E,4);
TASK_PP(16'h590F,4);
TASK_PP(16'h5910,4);
TASK_PP(16'h5911,4);
TASK_PP(16'h5912,4);
TASK_PP(16'h5913,4);
TASK_PP(16'h5914,4);
TASK_PP(16'h5915,4);
TASK_PP(16'h5916,4);
TASK_PP(16'h5917,4);
TASK_PP(16'h5918,4);
TASK_PP(16'h5919,4);
TASK_PP(16'h591A,4);
TASK_PP(16'h591B,4);
TASK_PP(16'h591C,4);
TASK_PP(16'h591D,4);
TASK_PP(16'h591E,4);
TASK_PP(16'h591F,4);
TASK_PP(16'h5920,4);
TASK_PP(16'h5921,4);
TASK_PP(16'h5922,4);
TASK_PP(16'h5923,4);
TASK_PP(16'h5924,4);
TASK_PP(16'h5925,4);
TASK_PP(16'h5926,4);
TASK_PP(16'h5927,4);
TASK_PP(16'h5928,4);
TASK_PP(16'h5929,4);
TASK_PP(16'h592A,4);
TASK_PP(16'h592B,4);
TASK_PP(16'h592C,4);
TASK_PP(16'h592D,4);
TASK_PP(16'h592E,4);
TASK_PP(16'h592F,4);
TASK_PP(16'h5930,4);
TASK_PP(16'h5931,4);
TASK_PP(16'h5932,4);
TASK_PP(16'h5933,4);
TASK_PP(16'h5934,4);
TASK_PP(16'h5935,4);
TASK_PP(16'h5936,4);
TASK_PP(16'h5937,4);
TASK_PP(16'h5938,4);
TASK_PP(16'h5939,4);
TASK_PP(16'h593A,4);
TASK_PP(16'h593B,4);
TASK_PP(16'h593C,4);
TASK_PP(16'h593D,4);
TASK_PP(16'h593E,4);
TASK_PP(16'h593F,4);
TASK_PP(16'h5940,4);
TASK_PP(16'h5941,4);
TASK_PP(16'h5942,4);
TASK_PP(16'h5943,4);
TASK_PP(16'h5944,4);
TASK_PP(16'h5945,4);
TASK_PP(16'h5946,4);
TASK_PP(16'h5947,4);
TASK_PP(16'h5948,4);
TASK_PP(16'h5949,4);
TASK_PP(16'h594A,4);
TASK_PP(16'h594B,4);
TASK_PP(16'h594C,4);
TASK_PP(16'h594D,4);
TASK_PP(16'h594E,4);
TASK_PP(16'h594F,4);
TASK_PP(16'h5950,4);
TASK_PP(16'h5951,4);
TASK_PP(16'h5952,4);
TASK_PP(16'h5953,4);
TASK_PP(16'h5954,4);
TASK_PP(16'h5955,4);
TASK_PP(16'h5956,4);
TASK_PP(16'h5957,4);
TASK_PP(16'h5958,4);
TASK_PP(16'h5959,4);
TASK_PP(16'h595A,4);
TASK_PP(16'h595B,4);
TASK_PP(16'h595C,4);
TASK_PP(16'h595D,4);
TASK_PP(16'h595E,4);
TASK_PP(16'h595F,4);
TASK_PP(16'h5960,4);
TASK_PP(16'h5961,4);
TASK_PP(16'h5962,4);
TASK_PP(16'h5963,4);
TASK_PP(16'h5964,4);
TASK_PP(16'h5965,4);
TASK_PP(16'h5966,4);
TASK_PP(16'h5967,4);
TASK_PP(16'h5968,4);
TASK_PP(16'h5969,4);
TASK_PP(16'h596A,4);
TASK_PP(16'h596B,4);
TASK_PP(16'h596C,4);
TASK_PP(16'h596D,4);
TASK_PP(16'h596E,4);
TASK_PP(16'h596F,4);
TASK_PP(16'h5970,4);
TASK_PP(16'h5971,4);
TASK_PP(16'h5972,4);
TASK_PP(16'h5973,4);
TASK_PP(16'h5974,4);
TASK_PP(16'h5975,4);
TASK_PP(16'h5976,4);
TASK_PP(16'h5977,4);
TASK_PP(16'h5978,4);
TASK_PP(16'h5979,4);
TASK_PP(16'h597A,4);
TASK_PP(16'h597B,4);
TASK_PP(16'h597C,4);
TASK_PP(16'h597D,4);
TASK_PP(16'h597E,4);
TASK_PP(16'h597F,4);
TASK_PP(16'h5980,4);
TASK_PP(16'h5981,4);
TASK_PP(16'h5982,4);
TASK_PP(16'h5983,4);
TASK_PP(16'h5984,4);
TASK_PP(16'h5985,4);
TASK_PP(16'h5986,4);
TASK_PP(16'h5987,4);
TASK_PP(16'h5988,4);
TASK_PP(16'h5989,4);
TASK_PP(16'h598A,4);
TASK_PP(16'h598B,4);
TASK_PP(16'h598C,4);
TASK_PP(16'h598D,4);
TASK_PP(16'h598E,4);
TASK_PP(16'h598F,4);
TASK_PP(16'h5990,4);
TASK_PP(16'h5991,4);
TASK_PP(16'h5992,4);
TASK_PP(16'h5993,4);
TASK_PP(16'h5994,4);
TASK_PP(16'h5995,4);
TASK_PP(16'h5996,4);
TASK_PP(16'h5997,4);
TASK_PP(16'h5998,4);
TASK_PP(16'h5999,4);
TASK_PP(16'h599A,4);
TASK_PP(16'h599B,4);
TASK_PP(16'h599C,4);
TASK_PP(16'h599D,4);
TASK_PP(16'h599E,4);
TASK_PP(16'h599F,4);
TASK_PP(16'h59A0,4);
TASK_PP(16'h59A1,4);
TASK_PP(16'h59A2,4);
TASK_PP(16'h59A3,4);
TASK_PP(16'h59A4,4);
TASK_PP(16'h59A5,4);
TASK_PP(16'h59A6,4);
TASK_PP(16'h59A7,4);
TASK_PP(16'h59A8,4);
TASK_PP(16'h59A9,4);
TASK_PP(16'h59AA,4);
TASK_PP(16'h59AB,4);
TASK_PP(16'h59AC,4);
TASK_PP(16'h59AD,4);
TASK_PP(16'h59AE,4);
TASK_PP(16'h59AF,4);
TASK_PP(16'h59B0,4);
TASK_PP(16'h59B1,4);
TASK_PP(16'h59B2,4);
TASK_PP(16'h59B3,4);
TASK_PP(16'h59B4,4);
TASK_PP(16'h59B5,4);
TASK_PP(16'h59B6,4);
TASK_PP(16'h59B7,4);
TASK_PP(16'h59B8,4);
TASK_PP(16'h59B9,4);
TASK_PP(16'h59BA,4);
TASK_PP(16'h59BB,4);
TASK_PP(16'h59BC,4);
TASK_PP(16'h59BD,4);
TASK_PP(16'h59BE,4);
TASK_PP(16'h59BF,4);
TASK_PP(16'h59C0,4);
TASK_PP(16'h59C1,4);
TASK_PP(16'h59C2,4);
TASK_PP(16'h59C3,4);
TASK_PP(16'h59C4,4);
TASK_PP(16'h59C5,4);
TASK_PP(16'h59C6,4);
TASK_PP(16'h59C7,4);
TASK_PP(16'h59C8,4);
TASK_PP(16'h59C9,4);
TASK_PP(16'h59CA,4);
TASK_PP(16'h59CB,4);
TASK_PP(16'h59CC,4);
TASK_PP(16'h59CD,4);
TASK_PP(16'h59CE,4);
TASK_PP(16'h59CF,4);
TASK_PP(16'h59D0,4);
TASK_PP(16'h59D1,4);
TASK_PP(16'h59D2,4);
TASK_PP(16'h59D3,4);
TASK_PP(16'h59D4,4);
TASK_PP(16'h59D5,4);
TASK_PP(16'h59D6,4);
TASK_PP(16'h59D7,4);
TASK_PP(16'h59D8,4);
TASK_PP(16'h59D9,4);
TASK_PP(16'h59DA,4);
TASK_PP(16'h59DB,4);
TASK_PP(16'h59DC,4);
TASK_PP(16'h59DD,4);
TASK_PP(16'h59DE,4);
TASK_PP(16'h59DF,4);
TASK_PP(16'h59E0,4);
TASK_PP(16'h59E1,4);
TASK_PP(16'h59E2,4);
TASK_PP(16'h59E3,4);
TASK_PP(16'h59E4,4);
TASK_PP(16'h59E5,4);
TASK_PP(16'h59E6,4);
TASK_PP(16'h59E7,4);
TASK_PP(16'h59E8,4);
TASK_PP(16'h59E9,4);
TASK_PP(16'h59EA,4);
TASK_PP(16'h59EB,4);
TASK_PP(16'h59EC,4);
TASK_PP(16'h59ED,4);
TASK_PP(16'h59EE,4);
TASK_PP(16'h59EF,4);
TASK_PP(16'h59F0,4);
TASK_PP(16'h59F1,4);
TASK_PP(16'h59F2,4);
TASK_PP(16'h59F3,4);
TASK_PP(16'h59F4,4);
TASK_PP(16'h59F5,4);
TASK_PP(16'h59F6,4);
TASK_PP(16'h59F7,4);
TASK_PP(16'h59F8,4);
TASK_PP(16'h59F9,4);
TASK_PP(16'h59FA,4);
TASK_PP(16'h59FB,4);
TASK_PP(16'h59FC,4);
TASK_PP(16'h59FD,4);
TASK_PP(16'h59FE,4);
TASK_PP(16'h59FF,4);
TASK_PP(16'h5A00,4);
TASK_PP(16'h5A01,4);
TASK_PP(16'h5A02,4);
TASK_PP(16'h5A03,4);
TASK_PP(16'h5A04,4);
TASK_PP(16'h5A05,4);
TASK_PP(16'h5A06,4);
TASK_PP(16'h5A07,4);
TASK_PP(16'h5A08,4);
TASK_PP(16'h5A09,4);
TASK_PP(16'h5A0A,4);
TASK_PP(16'h5A0B,4);
TASK_PP(16'h5A0C,4);
TASK_PP(16'h5A0D,4);
TASK_PP(16'h5A0E,4);
TASK_PP(16'h5A0F,4);
TASK_PP(16'h5A10,4);
TASK_PP(16'h5A11,4);
TASK_PP(16'h5A12,4);
TASK_PP(16'h5A13,4);
TASK_PP(16'h5A14,4);
TASK_PP(16'h5A15,4);
TASK_PP(16'h5A16,4);
TASK_PP(16'h5A17,4);
TASK_PP(16'h5A18,4);
TASK_PP(16'h5A19,4);
TASK_PP(16'h5A1A,4);
TASK_PP(16'h5A1B,4);
TASK_PP(16'h5A1C,4);
TASK_PP(16'h5A1D,4);
TASK_PP(16'h5A1E,4);
TASK_PP(16'h5A1F,4);
TASK_PP(16'h5A20,4);
TASK_PP(16'h5A21,4);
TASK_PP(16'h5A22,4);
TASK_PP(16'h5A23,4);
TASK_PP(16'h5A24,4);
TASK_PP(16'h5A25,4);
TASK_PP(16'h5A26,4);
TASK_PP(16'h5A27,4);
TASK_PP(16'h5A28,4);
TASK_PP(16'h5A29,4);
TASK_PP(16'h5A2A,4);
TASK_PP(16'h5A2B,4);
TASK_PP(16'h5A2C,4);
TASK_PP(16'h5A2D,4);
TASK_PP(16'h5A2E,4);
TASK_PP(16'h5A2F,4);
TASK_PP(16'h5A30,4);
TASK_PP(16'h5A31,4);
TASK_PP(16'h5A32,4);
TASK_PP(16'h5A33,4);
TASK_PP(16'h5A34,4);
TASK_PP(16'h5A35,4);
TASK_PP(16'h5A36,4);
TASK_PP(16'h5A37,4);
TASK_PP(16'h5A38,4);
TASK_PP(16'h5A39,4);
TASK_PP(16'h5A3A,4);
TASK_PP(16'h5A3B,4);
TASK_PP(16'h5A3C,4);
TASK_PP(16'h5A3D,4);
TASK_PP(16'h5A3E,4);
TASK_PP(16'h5A3F,4);
TASK_PP(16'h5A40,4);
TASK_PP(16'h5A41,4);
TASK_PP(16'h5A42,4);
TASK_PP(16'h5A43,4);
TASK_PP(16'h5A44,4);
TASK_PP(16'h5A45,4);
TASK_PP(16'h5A46,4);
TASK_PP(16'h5A47,4);
TASK_PP(16'h5A48,4);
TASK_PP(16'h5A49,4);
TASK_PP(16'h5A4A,4);
TASK_PP(16'h5A4B,4);
TASK_PP(16'h5A4C,4);
TASK_PP(16'h5A4D,4);
TASK_PP(16'h5A4E,4);
TASK_PP(16'h5A4F,4);
TASK_PP(16'h5A50,4);
TASK_PP(16'h5A51,4);
TASK_PP(16'h5A52,4);
TASK_PP(16'h5A53,4);
TASK_PP(16'h5A54,4);
TASK_PP(16'h5A55,4);
TASK_PP(16'h5A56,4);
TASK_PP(16'h5A57,4);
TASK_PP(16'h5A58,4);
TASK_PP(16'h5A59,4);
TASK_PP(16'h5A5A,4);
TASK_PP(16'h5A5B,4);
TASK_PP(16'h5A5C,4);
TASK_PP(16'h5A5D,4);
TASK_PP(16'h5A5E,4);
TASK_PP(16'h5A5F,4);
TASK_PP(16'h5A60,4);
TASK_PP(16'h5A61,4);
TASK_PP(16'h5A62,4);
TASK_PP(16'h5A63,4);
TASK_PP(16'h5A64,4);
TASK_PP(16'h5A65,4);
TASK_PP(16'h5A66,4);
TASK_PP(16'h5A67,4);
TASK_PP(16'h5A68,4);
TASK_PP(16'h5A69,4);
TASK_PP(16'h5A6A,4);
TASK_PP(16'h5A6B,4);
TASK_PP(16'h5A6C,4);
TASK_PP(16'h5A6D,4);
TASK_PP(16'h5A6E,4);
TASK_PP(16'h5A6F,4);
TASK_PP(16'h5A70,4);
TASK_PP(16'h5A71,4);
TASK_PP(16'h5A72,4);
TASK_PP(16'h5A73,4);
TASK_PP(16'h5A74,4);
TASK_PP(16'h5A75,4);
TASK_PP(16'h5A76,4);
TASK_PP(16'h5A77,4);
TASK_PP(16'h5A78,4);
TASK_PP(16'h5A79,4);
TASK_PP(16'h5A7A,4);
TASK_PP(16'h5A7B,4);
TASK_PP(16'h5A7C,4);
TASK_PP(16'h5A7D,4);
TASK_PP(16'h5A7E,4);
TASK_PP(16'h5A7F,4);
TASK_PP(16'h5A80,4);
TASK_PP(16'h5A81,4);
TASK_PP(16'h5A82,4);
TASK_PP(16'h5A83,4);
TASK_PP(16'h5A84,4);
TASK_PP(16'h5A85,4);
TASK_PP(16'h5A86,4);
TASK_PP(16'h5A87,4);
TASK_PP(16'h5A88,4);
TASK_PP(16'h5A89,4);
TASK_PP(16'h5A8A,4);
TASK_PP(16'h5A8B,4);
TASK_PP(16'h5A8C,4);
TASK_PP(16'h5A8D,4);
TASK_PP(16'h5A8E,4);
TASK_PP(16'h5A8F,4);
TASK_PP(16'h5A90,4);
TASK_PP(16'h5A91,4);
TASK_PP(16'h5A92,4);
TASK_PP(16'h5A93,4);
TASK_PP(16'h5A94,4);
TASK_PP(16'h5A95,4);
TASK_PP(16'h5A96,4);
TASK_PP(16'h5A97,4);
TASK_PP(16'h5A98,4);
TASK_PP(16'h5A99,4);
TASK_PP(16'h5A9A,4);
TASK_PP(16'h5A9B,4);
TASK_PP(16'h5A9C,4);
TASK_PP(16'h5A9D,4);
TASK_PP(16'h5A9E,4);
TASK_PP(16'h5A9F,4);
TASK_PP(16'h5AA0,4);
TASK_PP(16'h5AA1,4);
TASK_PP(16'h5AA2,4);
TASK_PP(16'h5AA3,4);
TASK_PP(16'h5AA4,4);
TASK_PP(16'h5AA5,4);
TASK_PP(16'h5AA6,4);
TASK_PP(16'h5AA7,4);
TASK_PP(16'h5AA8,4);
TASK_PP(16'h5AA9,4);
TASK_PP(16'h5AAA,4);
TASK_PP(16'h5AAB,4);
TASK_PP(16'h5AAC,4);
TASK_PP(16'h5AAD,4);
TASK_PP(16'h5AAE,4);
TASK_PP(16'h5AAF,4);
TASK_PP(16'h5AB0,4);
TASK_PP(16'h5AB1,4);
TASK_PP(16'h5AB2,4);
TASK_PP(16'h5AB3,4);
TASK_PP(16'h5AB4,4);
TASK_PP(16'h5AB5,4);
TASK_PP(16'h5AB6,4);
TASK_PP(16'h5AB7,4);
TASK_PP(16'h5AB8,4);
TASK_PP(16'h5AB9,4);
TASK_PP(16'h5ABA,4);
TASK_PP(16'h5ABB,4);
TASK_PP(16'h5ABC,4);
TASK_PP(16'h5ABD,4);
TASK_PP(16'h5ABE,4);
TASK_PP(16'h5ABF,4);
TASK_PP(16'h5AC0,4);
TASK_PP(16'h5AC1,4);
TASK_PP(16'h5AC2,4);
TASK_PP(16'h5AC3,4);
TASK_PP(16'h5AC4,4);
TASK_PP(16'h5AC5,4);
TASK_PP(16'h5AC6,4);
TASK_PP(16'h5AC7,4);
TASK_PP(16'h5AC8,4);
TASK_PP(16'h5AC9,4);
TASK_PP(16'h5ACA,4);
TASK_PP(16'h5ACB,4);
TASK_PP(16'h5ACC,4);
TASK_PP(16'h5ACD,4);
TASK_PP(16'h5ACE,4);
TASK_PP(16'h5ACF,4);
TASK_PP(16'h5AD0,4);
TASK_PP(16'h5AD1,4);
TASK_PP(16'h5AD2,4);
TASK_PP(16'h5AD3,4);
TASK_PP(16'h5AD4,4);
TASK_PP(16'h5AD5,4);
TASK_PP(16'h5AD6,4);
TASK_PP(16'h5AD7,4);
TASK_PP(16'h5AD8,4);
TASK_PP(16'h5AD9,4);
TASK_PP(16'h5ADA,4);
TASK_PP(16'h5ADB,4);
TASK_PP(16'h5ADC,4);
TASK_PP(16'h5ADD,4);
TASK_PP(16'h5ADE,4);
TASK_PP(16'h5ADF,4);
TASK_PP(16'h5AE0,4);
TASK_PP(16'h5AE1,4);
TASK_PP(16'h5AE2,4);
TASK_PP(16'h5AE3,4);
TASK_PP(16'h5AE4,4);
TASK_PP(16'h5AE5,4);
TASK_PP(16'h5AE6,4);
TASK_PP(16'h5AE7,4);
TASK_PP(16'h5AE8,4);
TASK_PP(16'h5AE9,4);
TASK_PP(16'h5AEA,4);
TASK_PP(16'h5AEB,4);
TASK_PP(16'h5AEC,4);
TASK_PP(16'h5AED,4);
TASK_PP(16'h5AEE,4);
TASK_PP(16'h5AEF,4);
TASK_PP(16'h5AF0,4);
TASK_PP(16'h5AF1,4);
TASK_PP(16'h5AF2,4);
TASK_PP(16'h5AF3,4);
TASK_PP(16'h5AF4,4);
TASK_PP(16'h5AF5,4);
TASK_PP(16'h5AF6,4);
TASK_PP(16'h5AF7,4);
TASK_PP(16'h5AF8,4);
TASK_PP(16'h5AF9,4);
TASK_PP(16'h5AFA,4);
TASK_PP(16'h5AFB,4);
TASK_PP(16'h5AFC,4);
TASK_PP(16'h5AFD,4);
TASK_PP(16'h5AFE,4);
TASK_PP(16'h5AFF,4);
TASK_PP(16'h5B00,4);
TASK_PP(16'h5B01,4);
TASK_PP(16'h5B02,4);
TASK_PP(16'h5B03,4);
TASK_PP(16'h5B04,4);
TASK_PP(16'h5B05,4);
TASK_PP(16'h5B06,4);
TASK_PP(16'h5B07,4);
TASK_PP(16'h5B08,4);
TASK_PP(16'h5B09,4);
TASK_PP(16'h5B0A,4);
TASK_PP(16'h5B0B,4);
TASK_PP(16'h5B0C,4);
TASK_PP(16'h5B0D,4);
TASK_PP(16'h5B0E,4);
TASK_PP(16'h5B0F,4);
TASK_PP(16'h5B10,4);
TASK_PP(16'h5B11,4);
TASK_PP(16'h5B12,4);
TASK_PP(16'h5B13,4);
TASK_PP(16'h5B14,4);
TASK_PP(16'h5B15,4);
TASK_PP(16'h5B16,4);
TASK_PP(16'h5B17,4);
TASK_PP(16'h5B18,4);
TASK_PP(16'h5B19,4);
TASK_PP(16'h5B1A,4);
TASK_PP(16'h5B1B,4);
TASK_PP(16'h5B1C,4);
TASK_PP(16'h5B1D,4);
TASK_PP(16'h5B1E,4);
TASK_PP(16'h5B1F,4);
TASK_PP(16'h5B20,4);
TASK_PP(16'h5B21,4);
TASK_PP(16'h5B22,4);
TASK_PP(16'h5B23,4);
TASK_PP(16'h5B24,4);
TASK_PP(16'h5B25,4);
TASK_PP(16'h5B26,4);
TASK_PP(16'h5B27,4);
TASK_PP(16'h5B28,4);
TASK_PP(16'h5B29,4);
TASK_PP(16'h5B2A,4);
TASK_PP(16'h5B2B,4);
TASK_PP(16'h5B2C,4);
TASK_PP(16'h5B2D,4);
TASK_PP(16'h5B2E,4);
TASK_PP(16'h5B2F,4);
TASK_PP(16'h5B30,4);
TASK_PP(16'h5B31,4);
TASK_PP(16'h5B32,4);
TASK_PP(16'h5B33,4);
TASK_PP(16'h5B34,4);
TASK_PP(16'h5B35,4);
TASK_PP(16'h5B36,4);
TASK_PP(16'h5B37,4);
TASK_PP(16'h5B38,4);
TASK_PP(16'h5B39,4);
TASK_PP(16'h5B3A,4);
TASK_PP(16'h5B3B,4);
TASK_PP(16'h5B3C,4);
TASK_PP(16'h5B3D,4);
TASK_PP(16'h5B3E,4);
TASK_PP(16'h5B3F,4);
TASK_PP(16'h5B40,4);
TASK_PP(16'h5B41,4);
TASK_PP(16'h5B42,4);
TASK_PP(16'h5B43,4);
TASK_PP(16'h5B44,4);
TASK_PP(16'h5B45,4);
TASK_PP(16'h5B46,4);
TASK_PP(16'h5B47,4);
TASK_PP(16'h5B48,4);
TASK_PP(16'h5B49,4);
TASK_PP(16'h5B4A,4);
TASK_PP(16'h5B4B,4);
TASK_PP(16'h5B4C,4);
TASK_PP(16'h5B4D,4);
TASK_PP(16'h5B4E,4);
TASK_PP(16'h5B4F,4);
TASK_PP(16'h5B50,4);
TASK_PP(16'h5B51,4);
TASK_PP(16'h5B52,4);
TASK_PP(16'h5B53,4);
TASK_PP(16'h5B54,4);
TASK_PP(16'h5B55,4);
TASK_PP(16'h5B56,4);
TASK_PP(16'h5B57,4);
TASK_PP(16'h5B58,4);
TASK_PP(16'h5B59,4);
TASK_PP(16'h5B5A,4);
TASK_PP(16'h5B5B,4);
TASK_PP(16'h5B5C,4);
TASK_PP(16'h5B5D,4);
TASK_PP(16'h5B5E,4);
TASK_PP(16'h5B5F,4);
TASK_PP(16'h5B60,4);
TASK_PP(16'h5B61,4);
TASK_PP(16'h5B62,4);
TASK_PP(16'h5B63,4);
TASK_PP(16'h5B64,4);
TASK_PP(16'h5B65,4);
TASK_PP(16'h5B66,4);
TASK_PP(16'h5B67,4);
TASK_PP(16'h5B68,4);
TASK_PP(16'h5B69,4);
TASK_PP(16'h5B6A,4);
TASK_PP(16'h5B6B,4);
TASK_PP(16'h5B6C,4);
TASK_PP(16'h5B6D,4);
TASK_PP(16'h5B6E,4);
TASK_PP(16'h5B6F,4);
TASK_PP(16'h5B70,4);
TASK_PP(16'h5B71,4);
TASK_PP(16'h5B72,4);
TASK_PP(16'h5B73,4);
TASK_PP(16'h5B74,4);
TASK_PP(16'h5B75,4);
TASK_PP(16'h5B76,4);
TASK_PP(16'h5B77,4);
TASK_PP(16'h5B78,4);
TASK_PP(16'h5B79,4);
TASK_PP(16'h5B7A,4);
TASK_PP(16'h5B7B,4);
TASK_PP(16'h5B7C,4);
TASK_PP(16'h5B7D,4);
TASK_PP(16'h5B7E,4);
TASK_PP(16'h5B7F,4);
TASK_PP(16'h5B80,4);
TASK_PP(16'h5B81,4);
TASK_PP(16'h5B82,4);
TASK_PP(16'h5B83,4);
TASK_PP(16'h5B84,4);
TASK_PP(16'h5B85,4);
TASK_PP(16'h5B86,4);
TASK_PP(16'h5B87,4);
TASK_PP(16'h5B88,4);
TASK_PP(16'h5B89,4);
TASK_PP(16'h5B8A,4);
TASK_PP(16'h5B8B,4);
TASK_PP(16'h5B8C,4);
TASK_PP(16'h5B8D,4);
TASK_PP(16'h5B8E,4);
TASK_PP(16'h5B8F,4);
TASK_PP(16'h5B90,4);
TASK_PP(16'h5B91,4);
TASK_PP(16'h5B92,4);
TASK_PP(16'h5B93,4);
TASK_PP(16'h5B94,4);
TASK_PP(16'h5B95,4);
TASK_PP(16'h5B96,4);
TASK_PP(16'h5B97,4);
TASK_PP(16'h5B98,4);
TASK_PP(16'h5B99,4);
TASK_PP(16'h5B9A,4);
TASK_PP(16'h5B9B,4);
TASK_PP(16'h5B9C,4);
TASK_PP(16'h5B9D,4);
TASK_PP(16'h5B9E,4);
TASK_PP(16'h5B9F,4);
TASK_PP(16'h5BA0,4);
TASK_PP(16'h5BA1,4);
TASK_PP(16'h5BA2,4);
TASK_PP(16'h5BA3,4);
TASK_PP(16'h5BA4,4);
TASK_PP(16'h5BA5,4);
TASK_PP(16'h5BA6,4);
TASK_PP(16'h5BA7,4);
TASK_PP(16'h5BA8,4);
TASK_PP(16'h5BA9,4);
TASK_PP(16'h5BAA,4);
TASK_PP(16'h5BAB,4);
TASK_PP(16'h5BAC,4);
TASK_PP(16'h5BAD,4);
TASK_PP(16'h5BAE,4);
TASK_PP(16'h5BAF,4);
TASK_PP(16'h5BB0,4);
TASK_PP(16'h5BB1,4);
TASK_PP(16'h5BB2,4);
TASK_PP(16'h5BB3,4);
TASK_PP(16'h5BB4,4);
TASK_PP(16'h5BB5,4);
TASK_PP(16'h5BB6,4);
TASK_PP(16'h5BB7,4);
TASK_PP(16'h5BB8,4);
TASK_PP(16'h5BB9,4);
TASK_PP(16'h5BBA,4);
TASK_PP(16'h5BBB,4);
TASK_PP(16'h5BBC,4);
TASK_PP(16'h5BBD,4);
TASK_PP(16'h5BBE,4);
TASK_PP(16'h5BBF,4);
TASK_PP(16'h5BC0,4);
TASK_PP(16'h5BC1,4);
TASK_PP(16'h5BC2,4);
TASK_PP(16'h5BC3,4);
TASK_PP(16'h5BC4,4);
TASK_PP(16'h5BC5,4);
TASK_PP(16'h5BC6,4);
TASK_PP(16'h5BC7,4);
TASK_PP(16'h5BC8,4);
TASK_PP(16'h5BC9,4);
TASK_PP(16'h5BCA,4);
TASK_PP(16'h5BCB,4);
TASK_PP(16'h5BCC,4);
TASK_PP(16'h5BCD,4);
TASK_PP(16'h5BCE,4);
TASK_PP(16'h5BCF,4);
TASK_PP(16'h5BD0,4);
TASK_PP(16'h5BD1,4);
TASK_PP(16'h5BD2,4);
TASK_PP(16'h5BD3,4);
TASK_PP(16'h5BD4,4);
TASK_PP(16'h5BD5,4);
TASK_PP(16'h5BD6,4);
TASK_PP(16'h5BD7,4);
TASK_PP(16'h5BD8,4);
TASK_PP(16'h5BD9,4);
TASK_PP(16'h5BDA,4);
TASK_PP(16'h5BDB,4);
TASK_PP(16'h5BDC,4);
TASK_PP(16'h5BDD,4);
TASK_PP(16'h5BDE,4);
TASK_PP(16'h5BDF,4);
TASK_PP(16'h5BE0,4);
TASK_PP(16'h5BE1,4);
TASK_PP(16'h5BE2,4);
TASK_PP(16'h5BE3,4);
TASK_PP(16'h5BE4,4);
TASK_PP(16'h5BE5,4);
TASK_PP(16'h5BE6,4);
TASK_PP(16'h5BE7,4);
TASK_PP(16'h5BE8,4);
TASK_PP(16'h5BE9,4);
TASK_PP(16'h5BEA,4);
TASK_PP(16'h5BEB,4);
TASK_PP(16'h5BEC,4);
TASK_PP(16'h5BED,4);
TASK_PP(16'h5BEE,4);
TASK_PP(16'h5BEF,4);
TASK_PP(16'h5BF0,4);
TASK_PP(16'h5BF1,4);
TASK_PP(16'h5BF2,4);
TASK_PP(16'h5BF3,4);
TASK_PP(16'h5BF4,4);
TASK_PP(16'h5BF5,4);
TASK_PP(16'h5BF6,4);
TASK_PP(16'h5BF7,4);
TASK_PP(16'h5BF8,4);
TASK_PP(16'h5BF9,4);
TASK_PP(16'h5BFA,4);
TASK_PP(16'h5BFB,4);
TASK_PP(16'h5BFC,4);
TASK_PP(16'h5BFD,4);
TASK_PP(16'h5BFE,4);
TASK_PP(16'h5BFF,4);
TASK_PP(16'h5C00,4);
TASK_PP(16'h5C01,4);
TASK_PP(16'h5C02,4);
TASK_PP(16'h5C03,4);
TASK_PP(16'h5C04,4);
TASK_PP(16'h5C05,4);
TASK_PP(16'h5C06,4);
TASK_PP(16'h5C07,4);
TASK_PP(16'h5C08,4);
TASK_PP(16'h5C09,4);
TASK_PP(16'h5C0A,4);
TASK_PP(16'h5C0B,4);
TASK_PP(16'h5C0C,4);
TASK_PP(16'h5C0D,4);
TASK_PP(16'h5C0E,4);
TASK_PP(16'h5C0F,4);
TASK_PP(16'h5C10,4);
TASK_PP(16'h5C11,4);
TASK_PP(16'h5C12,4);
TASK_PP(16'h5C13,4);
TASK_PP(16'h5C14,4);
TASK_PP(16'h5C15,4);
TASK_PP(16'h5C16,4);
TASK_PP(16'h5C17,4);
TASK_PP(16'h5C18,4);
TASK_PP(16'h5C19,4);
TASK_PP(16'h5C1A,4);
TASK_PP(16'h5C1B,4);
TASK_PP(16'h5C1C,4);
TASK_PP(16'h5C1D,4);
TASK_PP(16'h5C1E,4);
TASK_PP(16'h5C1F,4);
TASK_PP(16'h5C20,4);
TASK_PP(16'h5C21,4);
TASK_PP(16'h5C22,4);
TASK_PP(16'h5C23,4);
TASK_PP(16'h5C24,4);
TASK_PP(16'h5C25,4);
TASK_PP(16'h5C26,4);
TASK_PP(16'h5C27,4);
TASK_PP(16'h5C28,4);
TASK_PP(16'h5C29,4);
TASK_PP(16'h5C2A,4);
TASK_PP(16'h5C2B,4);
TASK_PP(16'h5C2C,4);
TASK_PP(16'h5C2D,4);
TASK_PP(16'h5C2E,4);
TASK_PP(16'h5C2F,4);
TASK_PP(16'h5C30,4);
TASK_PP(16'h5C31,4);
TASK_PP(16'h5C32,4);
TASK_PP(16'h5C33,4);
TASK_PP(16'h5C34,4);
TASK_PP(16'h5C35,4);
TASK_PP(16'h5C36,4);
TASK_PP(16'h5C37,4);
TASK_PP(16'h5C38,4);
TASK_PP(16'h5C39,4);
TASK_PP(16'h5C3A,4);
TASK_PP(16'h5C3B,4);
TASK_PP(16'h5C3C,4);
TASK_PP(16'h5C3D,4);
TASK_PP(16'h5C3E,4);
TASK_PP(16'h5C3F,4);
TASK_PP(16'h5C40,4);
TASK_PP(16'h5C41,4);
TASK_PP(16'h5C42,4);
TASK_PP(16'h5C43,4);
TASK_PP(16'h5C44,4);
TASK_PP(16'h5C45,4);
TASK_PP(16'h5C46,4);
TASK_PP(16'h5C47,4);
TASK_PP(16'h5C48,4);
TASK_PP(16'h5C49,4);
TASK_PP(16'h5C4A,4);
TASK_PP(16'h5C4B,4);
TASK_PP(16'h5C4C,4);
TASK_PP(16'h5C4D,4);
TASK_PP(16'h5C4E,4);
TASK_PP(16'h5C4F,4);
TASK_PP(16'h5C50,4);
TASK_PP(16'h5C51,4);
TASK_PP(16'h5C52,4);
TASK_PP(16'h5C53,4);
TASK_PP(16'h5C54,4);
TASK_PP(16'h5C55,4);
TASK_PP(16'h5C56,4);
TASK_PP(16'h5C57,4);
TASK_PP(16'h5C58,4);
TASK_PP(16'h5C59,4);
TASK_PP(16'h5C5A,4);
TASK_PP(16'h5C5B,4);
TASK_PP(16'h5C5C,4);
TASK_PP(16'h5C5D,4);
TASK_PP(16'h5C5E,4);
TASK_PP(16'h5C5F,4);
TASK_PP(16'h5C60,4);
TASK_PP(16'h5C61,4);
TASK_PP(16'h5C62,4);
TASK_PP(16'h5C63,4);
TASK_PP(16'h5C64,4);
TASK_PP(16'h5C65,4);
TASK_PP(16'h5C66,4);
TASK_PP(16'h5C67,4);
TASK_PP(16'h5C68,4);
TASK_PP(16'h5C69,4);
TASK_PP(16'h5C6A,4);
TASK_PP(16'h5C6B,4);
TASK_PP(16'h5C6C,4);
TASK_PP(16'h5C6D,4);
TASK_PP(16'h5C6E,4);
TASK_PP(16'h5C6F,4);
TASK_PP(16'h5C70,4);
TASK_PP(16'h5C71,4);
TASK_PP(16'h5C72,4);
TASK_PP(16'h5C73,4);
TASK_PP(16'h5C74,4);
TASK_PP(16'h5C75,4);
TASK_PP(16'h5C76,4);
TASK_PP(16'h5C77,4);
TASK_PP(16'h5C78,4);
TASK_PP(16'h5C79,4);
TASK_PP(16'h5C7A,4);
TASK_PP(16'h5C7B,4);
TASK_PP(16'h5C7C,4);
TASK_PP(16'h5C7D,4);
TASK_PP(16'h5C7E,4);
TASK_PP(16'h5C7F,4);
TASK_PP(16'h5C80,4);
TASK_PP(16'h5C81,4);
TASK_PP(16'h5C82,4);
TASK_PP(16'h5C83,4);
TASK_PP(16'h5C84,4);
TASK_PP(16'h5C85,4);
TASK_PP(16'h5C86,4);
TASK_PP(16'h5C87,4);
TASK_PP(16'h5C88,4);
TASK_PP(16'h5C89,4);
TASK_PP(16'h5C8A,4);
TASK_PP(16'h5C8B,4);
TASK_PP(16'h5C8C,4);
TASK_PP(16'h5C8D,4);
TASK_PP(16'h5C8E,4);
TASK_PP(16'h5C8F,4);
TASK_PP(16'h5C90,4);
TASK_PP(16'h5C91,4);
TASK_PP(16'h5C92,4);
TASK_PP(16'h5C93,4);
TASK_PP(16'h5C94,4);
TASK_PP(16'h5C95,4);
TASK_PP(16'h5C96,4);
TASK_PP(16'h5C97,4);
TASK_PP(16'h5C98,4);
TASK_PP(16'h5C99,4);
TASK_PP(16'h5C9A,4);
TASK_PP(16'h5C9B,4);
TASK_PP(16'h5C9C,4);
TASK_PP(16'h5C9D,4);
TASK_PP(16'h5C9E,4);
TASK_PP(16'h5C9F,4);
TASK_PP(16'h5CA0,4);
TASK_PP(16'h5CA1,4);
TASK_PP(16'h5CA2,4);
TASK_PP(16'h5CA3,4);
TASK_PP(16'h5CA4,4);
TASK_PP(16'h5CA5,4);
TASK_PP(16'h5CA6,4);
TASK_PP(16'h5CA7,4);
TASK_PP(16'h5CA8,4);
TASK_PP(16'h5CA9,4);
TASK_PP(16'h5CAA,4);
TASK_PP(16'h5CAB,4);
TASK_PP(16'h5CAC,4);
TASK_PP(16'h5CAD,4);
TASK_PP(16'h5CAE,4);
TASK_PP(16'h5CAF,4);
TASK_PP(16'h5CB0,4);
TASK_PP(16'h5CB1,4);
TASK_PP(16'h5CB2,4);
TASK_PP(16'h5CB3,4);
TASK_PP(16'h5CB4,4);
TASK_PP(16'h5CB5,4);
TASK_PP(16'h5CB6,4);
TASK_PP(16'h5CB7,4);
TASK_PP(16'h5CB8,4);
TASK_PP(16'h5CB9,4);
TASK_PP(16'h5CBA,4);
TASK_PP(16'h5CBB,4);
TASK_PP(16'h5CBC,4);
TASK_PP(16'h5CBD,4);
TASK_PP(16'h5CBE,4);
TASK_PP(16'h5CBF,4);
TASK_PP(16'h5CC0,4);
TASK_PP(16'h5CC1,4);
TASK_PP(16'h5CC2,4);
TASK_PP(16'h5CC3,4);
TASK_PP(16'h5CC4,4);
TASK_PP(16'h5CC5,4);
TASK_PP(16'h5CC6,4);
TASK_PP(16'h5CC7,4);
TASK_PP(16'h5CC8,4);
TASK_PP(16'h5CC9,4);
TASK_PP(16'h5CCA,4);
TASK_PP(16'h5CCB,4);
TASK_PP(16'h5CCC,4);
TASK_PP(16'h5CCD,4);
TASK_PP(16'h5CCE,4);
TASK_PP(16'h5CCF,4);
TASK_PP(16'h5CD0,4);
TASK_PP(16'h5CD1,4);
TASK_PP(16'h5CD2,4);
TASK_PP(16'h5CD3,4);
TASK_PP(16'h5CD4,4);
TASK_PP(16'h5CD5,4);
TASK_PP(16'h5CD6,4);
TASK_PP(16'h5CD7,4);
TASK_PP(16'h5CD8,4);
TASK_PP(16'h5CD9,4);
TASK_PP(16'h5CDA,4);
TASK_PP(16'h5CDB,4);
TASK_PP(16'h5CDC,4);
TASK_PP(16'h5CDD,4);
TASK_PP(16'h5CDE,4);
TASK_PP(16'h5CDF,4);
TASK_PP(16'h5CE0,4);
TASK_PP(16'h5CE1,4);
TASK_PP(16'h5CE2,4);
TASK_PP(16'h5CE3,4);
TASK_PP(16'h5CE4,4);
TASK_PP(16'h5CE5,4);
TASK_PP(16'h5CE6,4);
TASK_PP(16'h5CE7,4);
TASK_PP(16'h5CE8,4);
TASK_PP(16'h5CE9,4);
TASK_PP(16'h5CEA,4);
TASK_PP(16'h5CEB,4);
TASK_PP(16'h5CEC,4);
TASK_PP(16'h5CED,4);
TASK_PP(16'h5CEE,4);
TASK_PP(16'h5CEF,4);
TASK_PP(16'h5CF0,4);
TASK_PP(16'h5CF1,4);
TASK_PP(16'h5CF2,4);
TASK_PP(16'h5CF3,4);
TASK_PP(16'h5CF4,4);
TASK_PP(16'h5CF5,4);
TASK_PP(16'h5CF6,4);
TASK_PP(16'h5CF7,4);
TASK_PP(16'h5CF8,4);
TASK_PP(16'h5CF9,4);
TASK_PP(16'h5CFA,4);
TASK_PP(16'h5CFB,4);
TASK_PP(16'h5CFC,4);
TASK_PP(16'h5CFD,4);
TASK_PP(16'h5CFE,4);
TASK_PP(16'h5CFF,4);
TASK_PP(16'h5D00,4);
TASK_PP(16'h5D01,4);
TASK_PP(16'h5D02,4);
TASK_PP(16'h5D03,4);
TASK_PP(16'h5D04,4);
TASK_PP(16'h5D05,4);
TASK_PP(16'h5D06,4);
TASK_PP(16'h5D07,4);
TASK_PP(16'h5D08,4);
TASK_PP(16'h5D09,4);
TASK_PP(16'h5D0A,4);
TASK_PP(16'h5D0B,4);
TASK_PP(16'h5D0C,4);
TASK_PP(16'h5D0D,4);
TASK_PP(16'h5D0E,4);
TASK_PP(16'h5D0F,4);
TASK_PP(16'h5D10,4);
TASK_PP(16'h5D11,4);
TASK_PP(16'h5D12,4);
TASK_PP(16'h5D13,4);
TASK_PP(16'h5D14,4);
TASK_PP(16'h5D15,4);
TASK_PP(16'h5D16,4);
TASK_PP(16'h5D17,4);
TASK_PP(16'h5D18,4);
TASK_PP(16'h5D19,4);
TASK_PP(16'h5D1A,4);
TASK_PP(16'h5D1B,4);
TASK_PP(16'h5D1C,4);
TASK_PP(16'h5D1D,4);
TASK_PP(16'h5D1E,4);
TASK_PP(16'h5D1F,4);
TASK_PP(16'h5D20,4);
TASK_PP(16'h5D21,4);
TASK_PP(16'h5D22,4);
TASK_PP(16'h5D23,4);
TASK_PP(16'h5D24,4);
TASK_PP(16'h5D25,4);
TASK_PP(16'h5D26,4);
TASK_PP(16'h5D27,4);
TASK_PP(16'h5D28,4);
TASK_PP(16'h5D29,4);
TASK_PP(16'h5D2A,4);
TASK_PP(16'h5D2B,4);
TASK_PP(16'h5D2C,4);
TASK_PP(16'h5D2D,4);
TASK_PP(16'h5D2E,4);
TASK_PP(16'h5D2F,4);
TASK_PP(16'h5D30,4);
TASK_PP(16'h5D31,4);
TASK_PP(16'h5D32,4);
TASK_PP(16'h5D33,4);
TASK_PP(16'h5D34,4);
TASK_PP(16'h5D35,4);
TASK_PP(16'h5D36,4);
TASK_PP(16'h5D37,4);
TASK_PP(16'h5D38,4);
TASK_PP(16'h5D39,4);
TASK_PP(16'h5D3A,4);
TASK_PP(16'h5D3B,4);
TASK_PP(16'h5D3C,4);
TASK_PP(16'h5D3D,4);
TASK_PP(16'h5D3E,4);
TASK_PP(16'h5D3F,4);
TASK_PP(16'h5D40,4);
TASK_PP(16'h5D41,4);
TASK_PP(16'h5D42,4);
TASK_PP(16'h5D43,4);
TASK_PP(16'h5D44,4);
TASK_PP(16'h5D45,4);
TASK_PP(16'h5D46,4);
TASK_PP(16'h5D47,4);
TASK_PP(16'h5D48,4);
TASK_PP(16'h5D49,4);
TASK_PP(16'h5D4A,4);
TASK_PP(16'h5D4B,4);
TASK_PP(16'h5D4C,4);
TASK_PP(16'h5D4D,4);
TASK_PP(16'h5D4E,4);
TASK_PP(16'h5D4F,4);
TASK_PP(16'h5D50,4);
TASK_PP(16'h5D51,4);
TASK_PP(16'h5D52,4);
TASK_PP(16'h5D53,4);
TASK_PP(16'h5D54,4);
TASK_PP(16'h5D55,4);
TASK_PP(16'h5D56,4);
TASK_PP(16'h5D57,4);
TASK_PP(16'h5D58,4);
TASK_PP(16'h5D59,4);
TASK_PP(16'h5D5A,4);
TASK_PP(16'h5D5B,4);
TASK_PP(16'h5D5C,4);
TASK_PP(16'h5D5D,4);
TASK_PP(16'h5D5E,4);
TASK_PP(16'h5D5F,4);
TASK_PP(16'h5D60,4);
TASK_PP(16'h5D61,4);
TASK_PP(16'h5D62,4);
TASK_PP(16'h5D63,4);
TASK_PP(16'h5D64,4);
TASK_PP(16'h5D65,4);
TASK_PP(16'h5D66,4);
TASK_PP(16'h5D67,4);
TASK_PP(16'h5D68,4);
TASK_PP(16'h5D69,4);
TASK_PP(16'h5D6A,4);
TASK_PP(16'h5D6B,4);
TASK_PP(16'h5D6C,4);
TASK_PP(16'h5D6D,4);
TASK_PP(16'h5D6E,4);
TASK_PP(16'h5D6F,4);
TASK_PP(16'h5D70,4);
TASK_PP(16'h5D71,4);
TASK_PP(16'h5D72,4);
TASK_PP(16'h5D73,4);
TASK_PP(16'h5D74,4);
TASK_PP(16'h5D75,4);
TASK_PP(16'h5D76,4);
TASK_PP(16'h5D77,4);
TASK_PP(16'h5D78,4);
TASK_PP(16'h5D79,4);
TASK_PP(16'h5D7A,4);
TASK_PP(16'h5D7B,4);
TASK_PP(16'h5D7C,4);
TASK_PP(16'h5D7D,4);
TASK_PP(16'h5D7E,4);
TASK_PP(16'h5D7F,4);
TASK_PP(16'h5D80,4);
TASK_PP(16'h5D81,4);
TASK_PP(16'h5D82,4);
TASK_PP(16'h5D83,4);
TASK_PP(16'h5D84,4);
TASK_PP(16'h5D85,4);
TASK_PP(16'h5D86,4);
TASK_PP(16'h5D87,4);
TASK_PP(16'h5D88,4);
TASK_PP(16'h5D89,4);
TASK_PP(16'h5D8A,4);
TASK_PP(16'h5D8B,4);
TASK_PP(16'h5D8C,4);
TASK_PP(16'h5D8D,4);
TASK_PP(16'h5D8E,4);
TASK_PP(16'h5D8F,4);
TASK_PP(16'h5D90,4);
TASK_PP(16'h5D91,4);
TASK_PP(16'h5D92,4);
TASK_PP(16'h5D93,4);
TASK_PP(16'h5D94,4);
TASK_PP(16'h5D95,4);
TASK_PP(16'h5D96,4);
TASK_PP(16'h5D97,4);
TASK_PP(16'h5D98,4);
TASK_PP(16'h5D99,4);
TASK_PP(16'h5D9A,4);
TASK_PP(16'h5D9B,4);
TASK_PP(16'h5D9C,4);
TASK_PP(16'h5D9D,4);
TASK_PP(16'h5D9E,4);
TASK_PP(16'h5D9F,4);
TASK_PP(16'h5DA0,4);
TASK_PP(16'h5DA1,4);
TASK_PP(16'h5DA2,4);
TASK_PP(16'h5DA3,4);
TASK_PP(16'h5DA4,4);
TASK_PP(16'h5DA5,4);
TASK_PP(16'h5DA6,4);
TASK_PP(16'h5DA7,4);
TASK_PP(16'h5DA8,4);
TASK_PP(16'h5DA9,4);
TASK_PP(16'h5DAA,4);
TASK_PP(16'h5DAB,4);
TASK_PP(16'h5DAC,4);
TASK_PP(16'h5DAD,4);
TASK_PP(16'h5DAE,4);
TASK_PP(16'h5DAF,4);
TASK_PP(16'h5DB0,4);
TASK_PP(16'h5DB1,4);
TASK_PP(16'h5DB2,4);
TASK_PP(16'h5DB3,4);
TASK_PP(16'h5DB4,4);
TASK_PP(16'h5DB5,4);
TASK_PP(16'h5DB6,4);
TASK_PP(16'h5DB7,4);
TASK_PP(16'h5DB8,4);
TASK_PP(16'h5DB9,4);
TASK_PP(16'h5DBA,4);
TASK_PP(16'h5DBB,4);
TASK_PP(16'h5DBC,4);
TASK_PP(16'h5DBD,4);
TASK_PP(16'h5DBE,4);
TASK_PP(16'h5DBF,4);
TASK_PP(16'h5DC0,4);
TASK_PP(16'h5DC1,4);
TASK_PP(16'h5DC2,4);
TASK_PP(16'h5DC3,4);
TASK_PP(16'h5DC4,4);
TASK_PP(16'h5DC5,4);
TASK_PP(16'h5DC6,4);
TASK_PP(16'h5DC7,4);
TASK_PP(16'h5DC8,4);
TASK_PP(16'h5DC9,4);
TASK_PP(16'h5DCA,4);
TASK_PP(16'h5DCB,4);
TASK_PP(16'h5DCC,4);
TASK_PP(16'h5DCD,4);
TASK_PP(16'h5DCE,4);
TASK_PP(16'h5DCF,4);
TASK_PP(16'h5DD0,4);
TASK_PP(16'h5DD1,4);
TASK_PP(16'h5DD2,4);
TASK_PP(16'h5DD3,4);
TASK_PP(16'h5DD4,4);
TASK_PP(16'h5DD5,4);
TASK_PP(16'h5DD6,4);
TASK_PP(16'h5DD7,4);
TASK_PP(16'h5DD8,4);
TASK_PP(16'h5DD9,4);
TASK_PP(16'h5DDA,4);
TASK_PP(16'h5DDB,4);
TASK_PP(16'h5DDC,4);
TASK_PP(16'h5DDD,4);
TASK_PP(16'h5DDE,4);
TASK_PP(16'h5DDF,4);
TASK_PP(16'h5DE0,4);
TASK_PP(16'h5DE1,4);
TASK_PP(16'h5DE2,4);
TASK_PP(16'h5DE3,4);
TASK_PP(16'h5DE4,4);
TASK_PP(16'h5DE5,4);
TASK_PP(16'h5DE6,4);
TASK_PP(16'h5DE7,4);
TASK_PP(16'h5DE8,4);
TASK_PP(16'h5DE9,4);
TASK_PP(16'h5DEA,4);
TASK_PP(16'h5DEB,4);
TASK_PP(16'h5DEC,4);
TASK_PP(16'h5DED,4);
TASK_PP(16'h5DEE,4);
TASK_PP(16'h5DEF,4);
TASK_PP(16'h5DF0,4);
TASK_PP(16'h5DF1,4);
TASK_PP(16'h5DF2,4);
TASK_PP(16'h5DF3,4);
TASK_PP(16'h5DF4,4);
TASK_PP(16'h5DF5,4);
TASK_PP(16'h5DF6,4);
TASK_PP(16'h5DF7,4);
TASK_PP(16'h5DF8,4);
TASK_PP(16'h5DF9,4);
TASK_PP(16'h5DFA,4);
TASK_PP(16'h5DFB,4);
TASK_PP(16'h5DFC,4);
TASK_PP(16'h5DFD,4);
TASK_PP(16'h5DFE,4);
TASK_PP(16'h5DFF,4);
TASK_PP(16'h5E00,4);
TASK_PP(16'h5E01,4);
TASK_PP(16'h5E02,4);
TASK_PP(16'h5E03,4);
TASK_PP(16'h5E04,4);
TASK_PP(16'h5E05,4);
TASK_PP(16'h5E06,4);
TASK_PP(16'h5E07,4);
TASK_PP(16'h5E08,4);
TASK_PP(16'h5E09,4);
TASK_PP(16'h5E0A,4);
TASK_PP(16'h5E0B,4);
TASK_PP(16'h5E0C,4);
TASK_PP(16'h5E0D,4);
TASK_PP(16'h5E0E,4);
TASK_PP(16'h5E0F,4);
TASK_PP(16'h5E10,4);
TASK_PP(16'h5E11,4);
TASK_PP(16'h5E12,4);
TASK_PP(16'h5E13,4);
TASK_PP(16'h5E14,4);
TASK_PP(16'h5E15,4);
TASK_PP(16'h5E16,4);
TASK_PP(16'h5E17,4);
TASK_PP(16'h5E18,4);
TASK_PP(16'h5E19,4);
TASK_PP(16'h5E1A,4);
TASK_PP(16'h5E1B,4);
TASK_PP(16'h5E1C,4);
TASK_PP(16'h5E1D,4);
TASK_PP(16'h5E1E,4);
TASK_PP(16'h5E1F,4);
TASK_PP(16'h5E20,4);
TASK_PP(16'h5E21,4);
TASK_PP(16'h5E22,4);
TASK_PP(16'h5E23,4);
TASK_PP(16'h5E24,4);
TASK_PP(16'h5E25,4);
TASK_PP(16'h5E26,4);
TASK_PP(16'h5E27,4);
TASK_PP(16'h5E28,4);
TASK_PP(16'h5E29,4);
TASK_PP(16'h5E2A,4);
TASK_PP(16'h5E2B,4);
TASK_PP(16'h5E2C,4);
TASK_PP(16'h5E2D,4);
TASK_PP(16'h5E2E,4);
TASK_PP(16'h5E2F,4);
TASK_PP(16'h5E30,4);
TASK_PP(16'h5E31,4);
TASK_PP(16'h5E32,4);
TASK_PP(16'h5E33,4);
TASK_PP(16'h5E34,4);
TASK_PP(16'h5E35,4);
TASK_PP(16'h5E36,4);
TASK_PP(16'h5E37,4);
TASK_PP(16'h5E38,4);
TASK_PP(16'h5E39,4);
TASK_PP(16'h5E3A,4);
TASK_PP(16'h5E3B,4);
TASK_PP(16'h5E3C,4);
TASK_PP(16'h5E3D,4);
TASK_PP(16'h5E3E,4);
TASK_PP(16'h5E3F,4);
TASK_PP(16'h5E40,4);
TASK_PP(16'h5E41,4);
TASK_PP(16'h5E42,4);
TASK_PP(16'h5E43,4);
TASK_PP(16'h5E44,4);
TASK_PP(16'h5E45,4);
TASK_PP(16'h5E46,4);
TASK_PP(16'h5E47,4);
TASK_PP(16'h5E48,4);
TASK_PP(16'h5E49,4);
TASK_PP(16'h5E4A,4);
TASK_PP(16'h5E4B,4);
TASK_PP(16'h5E4C,4);
TASK_PP(16'h5E4D,4);
TASK_PP(16'h5E4E,4);
TASK_PP(16'h5E4F,4);
TASK_PP(16'h5E50,4);
TASK_PP(16'h5E51,4);
TASK_PP(16'h5E52,4);
TASK_PP(16'h5E53,4);
TASK_PP(16'h5E54,4);
TASK_PP(16'h5E55,4);
TASK_PP(16'h5E56,4);
TASK_PP(16'h5E57,4);
TASK_PP(16'h5E58,4);
TASK_PP(16'h5E59,4);
TASK_PP(16'h5E5A,4);
TASK_PP(16'h5E5B,4);
TASK_PP(16'h5E5C,4);
TASK_PP(16'h5E5D,4);
TASK_PP(16'h5E5E,4);
TASK_PP(16'h5E5F,4);
TASK_PP(16'h5E60,4);
TASK_PP(16'h5E61,4);
TASK_PP(16'h5E62,4);
TASK_PP(16'h5E63,4);
TASK_PP(16'h5E64,4);
TASK_PP(16'h5E65,4);
TASK_PP(16'h5E66,4);
TASK_PP(16'h5E67,4);
TASK_PP(16'h5E68,4);
TASK_PP(16'h5E69,4);
TASK_PP(16'h5E6A,4);
TASK_PP(16'h5E6B,4);
TASK_PP(16'h5E6C,4);
TASK_PP(16'h5E6D,4);
TASK_PP(16'h5E6E,4);
TASK_PP(16'h5E6F,4);
TASK_PP(16'h5E70,4);
TASK_PP(16'h5E71,4);
TASK_PP(16'h5E72,4);
TASK_PP(16'h5E73,4);
TASK_PP(16'h5E74,4);
TASK_PP(16'h5E75,4);
TASK_PP(16'h5E76,4);
TASK_PP(16'h5E77,4);
TASK_PP(16'h5E78,4);
TASK_PP(16'h5E79,4);
TASK_PP(16'h5E7A,4);
TASK_PP(16'h5E7B,4);
TASK_PP(16'h5E7C,4);
TASK_PP(16'h5E7D,4);
TASK_PP(16'h5E7E,4);
TASK_PP(16'h5E7F,4);
TASK_PP(16'h5E80,4);
TASK_PP(16'h5E81,4);
TASK_PP(16'h5E82,4);
TASK_PP(16'h5E83,4);
TASK_PP(16'h5E84,4);
TASK_PP(16'h5E85,4);
TASK_PP(16'h5E86,4);
TASK_PP(16'h5E87,4);
TASK_PP(16'h5E88,4);
TASK_PP(16'h5E89,4);
TASK_PP(16'h5E8A,4);
TASK_PP(16'h5E8B,4);
TASK_PP(16'h5E8C,4);
TASK_PP(16'h5E8D,4);
TASK_PP(16'h5E8E,4);
TASK_PP(16'h5E8F,4);
TASK_PP(16'h5E90,4);
TASK_PP(16'h5E91,4);
TASK_PP(16'h5E92,4);
TASK_PP(16'h5E93,4);
TASK_PP(16'h5E94,4);
TASK_PP(16'h5E95,4);
TASK_PP(16'h5E96,4);
TASK_PP(16'h5E97,4);
TASK_PP(16'h5E98,4);
TASK_PP(16'h5E99,4);
TASK_PP(16'h5E9A,4);
TASK_PP(16'h5E9B,4);
TASK_PP(16'h5E9C,4);
TASK_PP(16'h5E9D,4);
TASK_PP(16'h5E9E,4);
TASK_PP(16'h5E9F,4);
TASK_PP(16'h5EA0,4);
TASK_PP(16'h5EA1,4);
TASK_PP(16'h5EA2,4);
TASK_PP(16'h5EA3,4);
TASK_PP(16'h5EA4,4);
TASK_PP(16'h5EA5,4);
TASK_PP(16'h5EA6,4);
TASK_PP(16'h5EA7,4);
TASK_PP(16'h5EA8,4);
TASK_PP(16'h5EA9,4);
TASK_PP(16'h5EAA,4);
TASK_PP(16'h5EAB,4);
TASK_PP(16'h5EAC,4);
TASK_PP(16'h5EAD,4);
TASK_PP(16'h5EAE,4);
TASK_PP(16'h5EAF,4);
TASK_PP(16'h5EB0,4);
TASK_PP(16'h5EB1,4);
TASK_PP(16'h5EB2,4);
TASK_PP(16'h5EB3,4);
TASK_PP(16'h5EB4,4);
TASK_PP(16'h5EB5,4);
TASK_PP(16'h5EB6,4);
TASK_PP(16'h5EB7,4);
TASK_PP(16'h5EB8,4);
TASK_PP(16'h5EB9,4);
TASK_PP(16'h5EBA,4);
TASK_PP(16'h5EBB,4);
TASK_PP(16'h5EBC,4);
TASK_PP(16'h5EBD,4);
TASK_PP(16'h5EBE,4);
TASK_PP(16'h5EBF,4);
TASK_PP(16'h5EC0,4);
TASK_PP(16'h5EC1,4);
TASK_PP(16'h5EC2,4);
TASK_PP(16'h5EC3,4);
TASK_PP(16'h5EC4,4);
TASK_PP(16'h5EC5,4);
TASK_PP(16'h5EC6,4);
TASK_PP(16'h5EC7,4);
TASK_PP(16'h5EC8,4);
TASK_PP(16'h5EC9,4);
TASK_PP(16'h5ECA,4);
TASK_PP(16'h5ECB,4);
TASK_PP(16'h5ECC,4);
TASK_PP(16'h5ECD,4);
TASK_PP(16'h5ECE,4);
TASK_PP(16'h5ECF,4);
TASK_PP(16'h5ED0,4);
TASK_PP(16'h5ED1,4);
TASK_PP(16'h5ED2,4);
TASK_PP(16'h5ED3,4);
TASK_PP(16'h5ED4,4);
TASK_PP(16'h5ED5,4);
TASK_PP(16'h5ED6,4);
TASK_PP(16'h5ED7,4);
TASK_PP(16'h5ED8,4);
TASK_PP(16'h5ED9,4);
TASK_PP(16'h5EDA,4);
TASK_PP(16'h5EDB,4);
TASK_PP(16'h5EDC,4);
TASK_PP(16'h5EDD,4);
TASK_PP(16'h5EDE,4);
TASK_PP(16'h5EDF,4);
TASK_PP(16'h5EE0,4);
TASK_PP(16'h5EE1,4);
TASK_PP(16'h5EE2,4);
TASK_PP(16'h5EE3,4);
TASK_PP(16'h5EE4,4);
TASK_PP(16'h5EE5,4);
TASK_PP(16'h5EE6,4);
TASK_PP(16'h5EE7,4);
TASK_PP(16'h5EE8,4);
TASK_PP(16'h5EE9,4);
TASK_PP(16'h5EEA,4);
TASK_PP(16'h5EEB,4);
TASK_PP(16'h5EEC,4);
TASK_PP(16'h5EED,4);
TASK_PP(16'h5EEE,4);
TASK_PP(16'h5EEF,4);
TASK_PP(16'h5EF0,4);
TASK_PP(16'h5EF1,4);
TASK_PP(16'h5EF2,4);
TASK_PP(16'h5EF3,4);
TASK_PP(16'h5EF4,4);
TASK_PP(16'h5EF5,4);
TASK_PP(16'h5EF6,4);
TASK_PP(16'h5EF7,4);
TASK_PP(16'h5EF8,4);
TASK_PP(16'h5EF9,4);
TASK_PP(16'h5EFA,4);
TASK_PP(16'h5EFB,4);
TASK_PP(16'h5EFC,4);
TASK_PP(16'h5EFD,4);
TASK_PP(16'h5EFE,4);
TASK_PP(16'h5EFF,4);
TASK_PP(16'h5F00,4);
TASK_PP(16'h5F01,4);
TASK_PP(16'h5F02,4);
TASK_PP(16'h5F03,4);
TASK_PP(16'h5F04,4);
TASK_PP(16'h5F05,4);
TASK_PP(16'h5F06,4);
TASK_PP(16'h5F07,4);
TASK_PP(16'h5F08,4);
TASK_PP(16'h5F09,4);
TASK_PP(16'h5F0A,4);
TASK_PP(16'h5F0B,4);
TASK_PP(16'h5F0C,4);
TASK_PP(16'h5F0D,4);
TASK_PP(16'h5F0E,4);
TASK_PP(16'h5F0F,4);
TASK_PP(16'h5F10,4);
TASK_PP(16'h5F11,4);
TASK_PP(16'h5F12,4);
TASK_PP(16'h5F13,4);
TASK_PP(16'h5F14,4);
TASK_PP(16'h5F15,4);
TASK_PP(16'h5F16,4);
TASK_PP(16'h5F17,4);
TASK_PP(16'h5F18,4);
TASK_PP(16'h5F19,4);
TASK_PP(16'h5F1A,4);
TASK_PP(16'h5F1B,4);
TASK_PP(16'h5F1C,4);
TASK_PP(16'h5F1D,4);
TASK_PP(16'h5F1E,4);
TASK_PP(16'h5F1F,4);
TASK_PP(16'h5F20,4);
TASK_PP(16'h5F21,4);
TASK_PP(16'h5F22,4);
TASK_PP(16'h5F23,4);
TASK_PP(16'h5F24,4);
TASK_PP(16'h5F25,4);
TASK_PP(16'h5F26,4);
TASK_PP(16'h5F27,4);
TASK_PP(16'h5F28,4);
TASK_PP(16'h5F29,4);
TASK_PP(16'h5F2A,4);
TASK_PP(16'h5F2B,4);
TASK_PP(16'h5F2C,4);
TASK_PP(16'h5F2D,4);
TASK_PP(16'h5F2E,4);
TASK_PP(16'h5F2F,4);
TASK_PP(16'h5F30,4);
TASK_PP(16'h5F31,4);
TASK_PP(16'h5F32,4);
TASK_PP(16'h5F33,4);
TASK_PP(16'h5F34,4);
TASK_PP(16'h5F35,4);
TASK_PP(16'h5F36,4);
TASK_PP(16'h5F37,4);
TASK_PP(16'h5F38,4);
TASK_PP(16'h5F39,4);
TASK_PP(16'h5F3A,4);
TASK_PP(16'h5F3B,4);
TASK_PP(16'h5F3C,4);
TASK_PP(16'h5F3D,4);
TASK_PP(16'h5F3E,4);
TASK_PP(16'h5F3F,4);
TASK_PP(16'h5F40,4);
TASK_PP(16'h5F41,4);
TASK_PP(16'h5F42,4);
TASK_PP(16'h5F43,4);
TASK_PP(16'h5F44,4);
TASK_PP(16'h5F45,4);
TASK_PP(16'h5F46,4);
TASK_PP(16'h5F47,4);
TASK_PP(16'h5F48,4);
TASK_PP(16'h5F49,4);
TASK_PP(16'h5F4A,4);
TASK_PP(16'h5F4B,4);
TASK_PP(16'h5F4C,4);
TASK_PP(16'h5F4D,4);
TASK_PP(16'h5F4E,4);
TASK_PP(16'h5F4F,4);
TASK_PP(16'h5F50,4);
TASK_PP(16'h5F51,4);
TASK_PP(16'h5F52,4);
TASK_PP(16'h5F53,4);
TASK_PP(16'h5F54,4);
TASK_PP(16'h5F55,4);
TASK_PP(16'h5F56,4);
TASK_PP(16'h5F57,4);
TASK_PP(16'h5F58,4);
TASK_PP(16'h5F59,4);
TASK_PP(16'h5F5A,4);
TASK_PP(16'h5F5B,4);
TASK_PP(16'h5F5C,4);
TASK_PP(16'h5F5D,4);
TASK_PP(16'h5F5E,4);
TASK_PP(16'h5F5F,4);
TASK_PP(16'h5F60,4);
TASK_PP(16'h5F61,4);
TASK_PP(16'h5F62,4);
TASK_PP(16'h5F63,4);
TASK_PP(16'h5F64,4);
TASK_PP(16'h5F65,4);
TASK_PP(16'h5F66,4);
TASK_PP(16'h5F67,4);
TASK_PP(16'h5F68,4);
TASK_PP(16'h5F69,4);
TASK_PP(16'h5F6A,4);
TASK_PP(16'h5F6B,4);
TASK_PP(16'h5F6C,4);
TASK_PP(16'h5F6D,4);
TASK_PP(16'h5F6E,4);
TASK_PP(16'h5F6F,4);
TASK_PP(16'h5F70,4);
TASK_PP(16'h5F71,4);
TASK_PP(16'h5F72,4);
TASK_PP(16'h5F73,4);
TASK_PP(16'h5F74,4);
TASK_PP(16'h5F75,4);
TASK_PP(16'h5F76,4);
TASK_PP(16'h5F77,4);
TASK_PP(16'h5F78,4);
TASK_PP(16'h5F79,4);
TASK_PP(16'h5F7A,4);
TASK_PP(16'h5F7B,4);
TASK_PP(16'h5F7C,4);
TASK_PP(16'h5F7D,4);
TASK_PP(16'h5F7E,4);
TASK_PP(16'h5F7F,4);
TASK_PP(16'h5F80,4);
TASK_PP(16'h5F81,4);
TASK_PP(16'h5F82,4);
TASK_PP(16'h5F83,4);
TASK_PP(16'h5F84,4);
TASK_PP(16'h5F85,4);
TASK_PP(16'h5F86,4);
TASK_PP(16'h5F87,4);
TASK_PP(16'h5F88,4);
TASK_PP(16'h5F89,4);
TASK_PP(16'h5F8A,4);
TASK_PP(16'h5F8B,4);
TASK_PP(16'h5F8C,4);
TASK_PP(16'h5F8D,4);
TASK_PP(16'h5F8E,4);
TASK_PP(16'h5F8F,4);
TASK_PP(16'h5F90,4);
TASK_PP(16'h5F91,4);
TASK_PP(16'h5F92,4);
TASK_PP(16'h5F93,4);
TASK_PP(16'h5F94,4);
TASK_PP(16'h5F95,4);
TASK_PP(16'h5F96,4);
TASK_PP(16'h5F97,4);
TASK_PP(16'h5F98,4);
TASK_PP(16'h5F99,4);
TASK_PP(16'h5F9A,4);
TASK_PP(16'h5F9B,4);
TASK_PP(16'h5F9C,4);
TASK_PP(16'h5F9D,4);
TASK_PP(16'h5F9E,4);
TASK_PP(16'h5F9F,4);
TASK_PP(16'h5FA0,4);
TASK_PP(16'h5FA1,4);
TASK_PP(16'h5FA2,4);
TASK_PP(16'h5FA3,4);
TASK_PP(16'h5FA4,4);
TASK_PP(16'h5FA5,4);
TASK_PP(16'h5FA6,4);
TASK_PP(16'h5FA7,4);
TASK_PP(16'h5FA8,4);
TASK_PP(16'h5FA9,4);
TASK_PP(16'h5FAA,4);
TASK_PP(16'h5FAB,4);
TASK_PP(16'h5FAC,4);
TASK_PP(16'h5FAD,4);
TASK_PP(16'h5FAE,4);
TASK_PP(16'h5FAF,4);
TASK_PP(16'h5FB0,4);
TASK_PP(16'h5FB1,4);
TASK_PP(16'h5FB2,4);
TASK_PP(16'h5FB3,4);
TASK_PP(16'h5FB4,4);
TASK_PP(16'h5FB5,4);
TASK_PP(16'h5FB6,4);
TASK_PP(16'h5FB7,4);
TASK_PP(16'h5FB8,4);
TASK_PP(16'h5FB9,4);
TASK_PP(16'h5FBA,4);
TASK_PP(16'h5FBB,4);
TASK_PP(16'h5FBC,4);
TASK_PP(16'h5FBD,4);
TASK_PP(16'h5FBE,4);
TASK_PP(16'h5FBF,4);
TASK_PP(16'h5FC0,4);
TASK_PP(16'h5FC1,4);
TASK_PP(16'h5FC2,4);
TASK_PP(16'h5FC3,4);
TASK_PP(16'h5FC4,4);
TASK_PP(16'h5FC5,4);
TASK_PP(16'h5FC6,4);
TASK_PP(16'h5FC7,4);
TASK_PP(16'h5FC8,4);
TASK_PP(16'h5FC9,4);
TASK_PP(16'h5FCA,4);
TASK_PP(16'h5FCB,4);
TASK_PP(16'h5FCC,4);
TASK_PP(16'h5FCD,4);
TASK_PP(16'h5FCE,4);
TASK_PP(16'h5FCF,4);
TASK_PP(16'h5FD0,4);
TASK_PP(16'h5FD1,4);
TASK_PP(16'h5FD2,4);
TASK_PP(16'h5FD3,4);
TASK_PP(16'h5FD4,4);
TASK_PP(16'h5FD5,4);
TASK_PP(16'h5FD6,4);
TASK_PP(16'h5FD7,4);
TASK_PP(16'h5FD8,4);
TASK_PP(16'h5FD9,4);
TASK_PP(16'h5FDA,4);
TASK_PP(16'h5FDB,4);
TASK_PP(16'h5FDC,4);
TASK_PP(16'h5FDD,4);
TASK_PP(16'h5FDE,4);
TASK_PP(16'h5FDF,4);
TASK_PP(16'h5FE0,4);
TASK_PP(16'h5FE1,4);
TASK_PP(16'h5FE2,4);
TASK_PP(16'h5FE3,4);
TASK_PP(16'h5FE4,4);
TASK_PP(16'h5FE5,4);
TASK_PP(16'h5FE6,4);
TASK_PP(16'h5FE7,4);
TASK_PP(16'h5FE8,4);
TASK_PP(16'h5FE9,4);
TASK_PP(16'h5FEA,4);
TASK_PP(16'h5FEB,4);
TASK_PP(16'h5FEC,4);
TASK_PP(16'h5FED,4);
TASK_PP(16'h5FEE,4);
TASK_PP(16'h5FEF,4);
TASK_PP(16'h5FF0,4);
TASK_PP(16'h5FF1,4);
TASK_PP(16'h5FF2,4);
TASK_PP(16'h5FF3,4);
TASK_PP(16'h5FF4,4);
TASK_PP(16'h5FF5,4);
TASK_PP(16'h5FF6,4);
TASK_PP(16'h5FF7,4);
TASK_PP(16'h5FF8,4);
TASK_PP(16'h5FF9,4);
TASK_PP(16'h5FFA,4);
TASK_PP(16'h5FFB,4);
TASK_PP(16'h5FFC,4);
TASK_PP(16'h5FFD,4);
TASK_PP(16'h5FFE,4);
TASK_PP(16'h5FFF,4);
TASK_PP(16'h6000,4);
TASK_PP(16'h6001,4);
TASK_PP(16'h6002,4);
TASK_PP(16'h6003,4);
TASK_PP(16'h6004,4);
TASK_PP(16'h6005,4);
TASK_PP(16'h6006,4);
TASK_PP(16'h6007,4);
TASK_PP(16'h6008,4);
TASK_PP(16'h6009,4);
TASK_PP(16'h600A,4);
TASK_PP(16'h600B,4);
TASK_PP(16'h600C,4);
TASK_PP(16'h600D,4);
TASK_PP(16'h600E,4);
TASK_PP(16'h600F,4);
TASK_PP(16'h6010,4);
TASK_PP(16'h6011,4);
TASK_PP(16'h6012,4);
TASK_PP(16'h6013,4);
TASK_PP(16'h6014,4);
TASK_PP(16'h6015,4);
TASK_PP(16'h6016,4);
TASK_PP(16'h6017,4);
TASK_PP(16'h6018,4);
TASK_PP(16'h6019,4);
TASK_PP(16'h601A,4);
TASK_PP(16'h601B,4);
TASK_PP(16'h601C,4);
TASK_PP(16'h601D,4);
TASK_PP(16'h601E,4);
TASK_PP(16'h601F,4);
TASK_PP(16'h6020,4);
TASK_PP(16'h6021,4);
TASK_PP(16'h6022,4);
TASK_PP(16'h6023,4);
TASK_PP(16'h6024,4);
TASK_PP(16'h6025,4);
TASK_PP(16'h6026,4);
TASK_PP(16'h6027,4);
TASK_PP(16'h6028,4);
TASK_PP(16'h6029,4);
TASK_PP(16'h602A,4);
TASK_PP(16'h602B,4);
TASK_PP(16'h602C,4);
TASK_PP(16'h602D,4);
TASK_PP(16'h602E,4);
TASK_PP(16'h602F,4);
TASK_PP(16'h6030,4);
TASK_PP(16'h6031,4);
TASK_PP(16'h6032,4);
TASK_PP(16'h6033,4);
TASK_PP(16'h6034,4);
TASK_PP(16'h6035,4);
TASK_PP(16'h6036,4);
TASK_PP(16'h6037,4);
TASK_PP(16'h6038,4);
TASK_PP(16'h6039,4);
TASK_PP(16'h603A,4);
TASK_PP(16'h603B,4);
TASK_PP(16'h603C,4);
TASK_PP(16'h603D,4);
TASK_PP(16'h603E,4);
TASK_PP(16'h603F,4);
TASK_PP(16'h6040,4);
TASK_PP(16'h6041,4);
TASK_PP(16'h6042,4);
TASK_PP(16'h6043,4);
TASK_PP(16'h6044,4);
TASK_PP(16'h6045,4);
TASK_PP(16'h6046,4);
TASK_PP(16'h6047,4);
TASK_PP(16'h6048,4);
TASK_PP(16'h6049,4);
TASK_PP(16'h604A,4);
TASK_PP(16'h604B,4);
TASK_PP(16'h604C,4);
TASK_PP(16'h604D,4);
TASK_PP(16'h604E,4);
TASK_PP(16'h604F,4);
TASK_PP(16'h6050,4);
TASK_PP(16'h6051,4);
TASK_PP(16'h6052,4);
TASK_PP(16'h6053,4);
TASK_PP(16'h6054,4);
TASK_PP(16'h6055,4);
TASK_PP(16'h6056,4);
TASK_PP(16'h6057,4);
TASK_PP(16'h6058,4);
TASK_PP(16'h6059,4);
TASK_PP(16'h605A,4);
TASK_PP(16'h605B,4);
TASK_PP(16'h605C,4);
TASK_PP(16'h605D,4);
TASK_PP(16'h605E,4);
TASK_PP(16'h605F,4);
TASK_PP(16'h6060,4);
TASK_PP(16'h6061,4);
TASK_PP(16'h6062,4);
TASK_PP(16'h6063,4);
TASK_PP(16'h6064,4);
TASK_PP(16'h6065,4);
TASK_PP(16'h6066,4);
TASK_PP(16'h6067,4);
TASK_PP(16'h6068,4);
TASK_PP(16'h6069,4);
TASK_PP(16'h606A,4);
TASK_PP(16'h606B,4);
TASK_PP(16'h606C,4);
TASK_PP(16'h606D,4);
TASK_PP(16'h606E,4);
TASK_PP(16'h606F,4);
TASK_PP(16'h6070,4);
TASK_PP(16'h6071,4);
TASK_PP(16'h6072,4);
TASK_PP(16'h6073,4);
TASK_PP(16'h6074,4);
TASK_PP(16'h6075,4);
TASK_PP(16'h6076,4);
TASK_PP(16'h6077,4);
TASK_PP(16'h6078,4);
TASK_PP(16'h6079,4);
TASK_PP(16'h607A,4);
TASK_PP(16'h607B,4);
TASK_PP(16'h607C,4);
TASK_PP(16'h607D,4);
TASK_PP(16'h607E,4);
TASK_PP(16'h607F,4);
TASK_PP(16'h6080,4);
TASK_PP(16'h6081,4);
TASK_PP(16'h6082,4);
TASK_PP(16'h6083,4);
TASK_PP(16'h6084,4);
TASK_PP(16'h6085,4);
TASK_PP(16'h6086,4);
TASK_PP(16'h6087,4);
TASK_PP(16'h6088,4);
TASK_PP(16'h6089,4);
TASK_PP(16'h608A,4);
TASK_PP(16'h608B,4);
TASK_PP(16'h608C,4);
TASK_PP(16'h608D,4);
TASK_PP(16'h608E,4);
TASK_PP(16'h608F,4);
TASK_PP(16'h6090,4);
TASK_PP(16'h6091,4);
TASK_PP(16'h6092,4);
TASK_PP(16'h6093,4);
TASK_PP(16'h6094,4);
TASK_PP(16'h6095,4);
TASK_PP(16'h6096,4);
TASK_PP(16'h6097,4);
TASK_PP(16'h6098,4);
TASK_PP(16'h6099,4);
TASK_PP(16'h609A,4);
TASK_PP(16'h609B,4);
TASK_PP(16'h609C,4);
TASK_PP(16'h609D,4);
TASK_PP(16'h609E,4);
TASK_PP(16'h609F,4);
TASK_PP(16'h60A0,4);
TASK_PP(16'h60A1,4);
TASK_PP(16'h60A2,4);
TASK_PP(16'h60A3,4);
TASK_PP(16'h60A4,4);
TASK_PP(16'h60A5,4);
TASK_PP(16'h60A6,4);
TASK_PP(16'h60A7,4);
TASK_PP(16'h60A8,4);
TASK_PP(16'h60A9,4);
TASK_PP(16'h60AA,4);
TASK_PP(16'h60AB,4);
TASK_PP(16'h60AC,4);
TASK_PP(16'h60AD,4);
TASK_PP(16'h60AE,4);
TASK_PP(16'h60AF,4);
TASK_PP(16'h60B0,4);
TASK_PP(16'h60B1,4);
TASK_PP(16'h60B2,4);
TASK_PP(16'h60B3,4);
TASK_PP(16'h60B4,4);
TASK_PP(16'h60B5,4);
TASK_PP(16'h60B6,4);
TASK_PP(16'h60B7,4);
TASK_PP(16'h60B8,4);
TASK_PP(16'h60B9,4);
TASK_PP(16'h60BA,4);
TASK_PP(16'h60BB,4);
TASK_PP(16'h60BC,4);
TASK_PP(16'h60BD,4);
TASK_PP(16'h60BE,4);
TASK_PP(16'h60BF,4);
TASK_PP(16'h60C0,4);
TASK_PP(16'h60C1,4);
TASK_PP(16'h60C2,4);
TASK_PP(16'h60C3,4);
TASK_PP(16'h60C4,4);
TASK_PP(16'h60C5,4);
TASK_PP(16'h60C6,4);
TASK_PP(16'h60C7,4);
TASK_PP(16'h60C8,4);
TASK_PP(16'h60C9,4);
TASK_PP(16'h60CA,4);
TASK_PP(16'h60CB,4);
TASK_PP(16'h60CC,4);
TASK_PP(16'h60CD,4);
TASK_PP(16'h60CE,4);
TASK_PP(16'h60CF,4);
TASK_PP(16'h60D0,4);
TASK_PP(16'h60D1,4);
TASK_PP(16'h60D2,4);
TASK_PP(16'h60D3,4);
TASK_PP(16'h60D4,4);
TASK_PP(16'h60D5,4);
TASK_PP(16'h60D6,4);
TASK_PP(16'h60D7,4);
TASK_PP(16'h60D8,4);
TASK_PP(16'h60D9,4);
TASK_PP(16'h60DA,4);
TASK_PP(16'h60DB,4);
TASK_PP(16'h60DC,4);
TASK_PP(16'h60DD,4);
TASK_PP(16'h60DE,4);
TASK_PP(16'h60DF,4);
TASK_PP(16'h60E0,4);
TASK_PP(16'h60E1,4);
TASK_PP(16'h60E2,4);
TASK_PP(16'h60E3,4);
TASK_PP(16'h60E4,4);
TASK_PP(16'h60E5,4);
TASK_PP(16'h60E6,4);
TASK_PP(16'h60E7,4);
TASK_PP(16'h60E8,4);
TASK_PP(16'h60E9,4);
TASK_PP(16'h60EA,4);
TASK_PP(16'h60EB,4);
TASK_PP(16'h60EC,4);
TASK_PP(16'h60ED,4);
TASK_PP(16'h60EE,4);
TASK_PP(16'h60EF,4);
TASK_PP(16'h60F0,4);
TASK_PP(16'h60F1,4);
TASK_PP(16'h60F2,4);
TASK_PP(16'h60F3,4);
TASK_PP(16'h60F4,4);
TASK_PP(16'h60F5,4);
TASK_PP(16'h60F6,4);
TASK_PP(16'h60F7,4);
TASK_PP(16'h60F8,4);
TASK_PP(16'h60F9,4);
TASK_PP(16'h60FA,4);
TASK_PP(16'h60FB,4);
TASK_PP(16'h60FC,4);
TASK_PP(16'h60FD,4);
TASK_PP(16'h60FE,4);
TASK_PP(16'h60FF,4);
TASK_PP(16'h6100,4);
TASK_PP(16'h6101,4);
TASK_PP(16'h6102,4);
TASK_PP(16'h6103,4);
TASK_PP(16'h6104,4);
TASK_PP(16'h6105,4);
TASK_PP(16'h6106,4);
TASK_PP(16'h6107,4);
TASK_PP(16'h6108,4);
TASK_PP(16'h6109,4);
TASK_PP(16'h610A,4);
TASK_PP(16'h610B,4);
TASK_PP(16'h610C,4);
TASK_PP(16'h610D,4);
TASK_PP(16'h610E,4);
TASK_PP(16'h610F,4);
TASK_PP(16'h6110,4);
TASK_PP(16'h6111,4);
TASK_PP(16'h6112,4);
TASK_PP(16'h6113,4);
TASK_PP(16'h6114,4);
TASK_PP(16'h6115,4);
TASK_PP(16'h6116,4);
TASK_PP(16'h6117,4);
TASK_PP(16'h6118,4);
TASK_PP(16'h6119,4);
TASK_PP(16'h611A,4);
TASK_PP(16'h611B,4);
TASK_PP(16'h611C,4);
TASK_PP(16'h611D,4);
TASK_PP(16'h611E,4);
TASK_PP(16'h611F,4);
TASK_PP(16'h6120,4);
TASK_PP(16'h6121,4);
TASK_PP(16'h6122,4);
TASK_PP(16'h6123,4);
TASK_PP(16'h6124,4);
TASK_PP(16'h6125,4);
TASK_PP(16'h6126,4);
TASK_PP(16'h6127,4);
TASK_PP(16'h6128,4);
TASK_PP(16'h6129,4);
TASK_PP(16'h612A,4);
TASK_PP(16'h612B,4);
TASK_PP(16'h612C,4);
TASK_PP(16'h612D,4);
TASK_PP(16'h612E,4);
TASK_PP(16'h612F,4);
TASK_PP(16'h6130,4);
TASK_PP(16'h6131,4);
TASK_PP(16'h6132,4);
TASK_PP(16'h6133,4);
TASK_PP(16'h6134,4);
TASK_PP(16'h6135,4);
TASK_PP(16'h6136,4);
TASK_PP(16'h6137,4);
TASK_PP(16'h6138,4);
TASK_PP(16'h6139,4);
TASK_PP(16'h613A,4);
TASK_PP(16'h613B,4);
TASK_PP(16'h613C,4);
TASK_PP(16'h613D,4);
TASK_PP(16'h613E,4);
TASK_PP(16'h613F,4);
TASK_PP(16'h6140,4);
TASK_PP(16'h6141,4);
TASK_PP(16'h6142,4);
TASK_PP(16'h6143,4);
TASK_PP(16'h6144,4);
TASK_PP(16'h6145,4);
TASK_PP(16'h6146,4);
TASK_PP(16'h6147,4);
TASK_PP(16'h6148,4);
TASK_PP(16'h6149,4);
TASK_PP(16'h614A,4);
TASK_PP(16'h614B,4);
TASK_PP(16'h614C,4);
TASK_PP(16'h614D,4);
TASK_PP(16'h614E,4);
TASK_PP(16'h614F,4);
TASK_PP(16'h6150,4);
TASK_PP(16'h6151,4);
TASK_PP(16'h6152,4);
TASK_PP(16'h6153,4);
TASK_PP(16'h6154,4);
TASK_PP(16'h6155,4);
TASK_PP(16'h6156,4);
TASK_PP(16'h6157,4);
TASK_PP(16'h6158,4);
TASK_PP(16'h6159,4);
TASK_PP(16'h615A,4);
TASK_PP(16'h615B,4);
TASK_PP(16'h615C,4);
TASK_PP(16'h615D,4);
TASK_PP(16'h615E,4);
TASK_PP(16'h615F,4);
TASK_PP(16'h6160,4);
TASK_PP(16'h6161,4);
TASK_PP(16'h6162,4);
TASK_PP(16'h6163,4);
TASK_PP(16'h6164,4);
TASK_PP(16'h6165,4);
TASK_PP(16'h6166,4);
TASK_PP(16'h6167,4);
TASK_PP(16'h6168,4);
TASK_PP(16'h6169,4);
TASK_PP(16'h616A,4);
TASK_PP(16'h616B,4);
TASK_PP(16'h616C,4);
TASK_PP(16'h616D,4);
TASK_PP(16'h616E,4);
TASK_PP(16'h616F,4);
TASK_PP(16'h6170,4);
TASK_PP(16'h6171,4);
TASK_PP(16'h6172,4);
TASK_PP(16'h6173,4);
TASK_PP(16'h6174,4);
TASK_PP(16'h6175,4);
TASK_PP(16'h6176,4);
TASK_PP(16'h6177,4);
TASK_PP(16'h6178,4);
TASK_PP(16'h6179,4);
TASK_PP(16'h617A,4);
TASK_PP(16'h617B,4);
TASK_PP(16'h617C,4);
TASK_PP(16'h617D,4);
TASK_PP(16'h617E,4);
TASK_PP(16'h617F,4);
TASK_PP(16'h6180,4);
TASK_PP(16'h6181,4);
TASK_PP(16'h6182,4);
TASK_PP(16'h6183,4);
TASK_PP(16'h6184,4);
TASK_PP(16'h6185,4);
TASK_PP(16'h6186,4);
TASK_PP(16'h6187,4);
TASK_PP(16'h6188,4);
TASK_PP(16'h6189,4);
TASK_PP(16'h618A,4);
TASK_PP(16'h618B,4);
TASK_PP(16'h618C,4);
TASK_PP(16'h618D,4);
TASK_PP(16'h618E,4);
TASK_PP(16'h618F,4);
TASK_PP(16'h6190,4);
TASK_PP(16'h6191,4);
TASK_PP(16'h6192,4);
TASK_PP(16'h6193,4);
TASK_PP(16'h6194,4);
TASK_PP(16'h6195,4);
TASK_PP(16'h6196,4);
TASK_PP(16'h6197,4);
TASK_PP(16'h6198,4);
TASK_PP(16'h6199,4);
TASK_PP(16'h619A,4);
TASK_PP(16'h619B,4);
TASK_PP(16'h619C,4);
TASK_PP(16'h619D,4);
TASK_PP(16'h619E,4);
TASK_PP(16'h619F,4);
TASK_PP(16'h61A0,4);
TASK_PP(16'h61A1,4);
TASK_PP(16'h61A2,4);
TASK_PP(16'h61A3,4);
TASK_PP(16'h61A4,4);
TASK_PP(16'h61A5,4);
TASK_PP(16'h61A6,4);
TASK_PP(16'h61A7,4);
TASK_PP(16'h61A8,4);
TASK_PP(16'h61A9,4);
TASK_PP(16'h61AA,4);
TASK_PP(16'h61AB,4);
TASK_PP(16'h61AC,4);
TASK_PP(16'h61AD,4);
TASK_PP(16'h61AE,4);
TASK_PP(16'h61AF,4);
TASK_PP(16'h61B0,4);
TASK_PP(16'h61B1,4);
TASK_PP(16'h61B2,4);
TASK_PP(16'h61B3,4);
TASK_PP(16'h61B4,4);
TASK_PP(16'h61B5,4);
TASK_PP(16'h61B6,4);
TASK_PP(16'h61B7,4);
TASK_PP(16'h61B8,4);
TASK_PP(16'h61B9,4);
TASK_PP(16'h61BA,4);
TASK_PP(16'h61BB,4);
TASK_PP(16'h61BC,4);
TASK_PP(16'h61BD,4);
TASK_PP(16'h61BE,4);
TASK_PP(16'h61BF,4);
TASK_PP(16'h61C0,4);
TASK_PP(16'h61C1,4);
TASK_PP(16'h61C2,4);
TASK_PP(16'h61C3,4);
TASK_PP(16'h61C4,4);
TASK_PP(16'h61C5,4);
TASK_PP(16'h61C6,4);
TASK_PP(16'h61C7,4);
TASK_PP(16'h61C8,4);
TASK_PP(16'h61C9,4);
TASK_PP(16'h61CA,4);
TASK_PP(16'h61CB,4);
TASK_PP(16'h61CC,4);
TASK_PP(16'h61CD,4);
TASK_PP(16'h61CE,4);
TASK_PP(16'h61CF,4);
TASK_PP(16'h61D0,4);
TASK_PP(16'h61D1,4);
TASK_PP(16'h61D2,4);
TASK_PP(16'h61D3,4);
TASK_PP(16'h61D4,4);
TASK_PP(16'h61D5,4);
TASK_PP(16'h61D6,4);
TASK_PP(16'h61D7,4);
TASK_PP(16'h61D8,4);
TASK_PP(16'h61D9,4);
TASK_PP(16'h61DA,4);
TASK_PP(16'h61DB,4);
TASK_PP(16'h61DC,4);
TASK_PP(16'h61DD,4);
TASK_PP(16'h61DE,4);
TASK_PP(16'h61DF,4);
TASK_PP(16'h61E0,4);
TASK_PP(16'h61E1,4);
TASK_PP(16'h61E2,4);
TASK_PP(16'h61E3,4);
TASK_PP(16'h61E4,4);
TASK_PP(16'h61E5,4);
TASK_PP(16'h61E6,4);
TASK_PP(16'h61E7,4);
TASK_PP(16'h61E8,4);
TASK_PP(16'h61E9,4);
TASK_PP(16'h61EA,4);
TASK_PP(16'h61EB,4);
TASK_PP(16'h61EC,4);
TASK_PP(16'h61ED,4);
TASK_PP(16'h61EE,4);
TASK_PP(16'h61EF,4);
TASK_PP(16'h61F0,4);
TASK_PP(16'h61F1,4);
TASK_PP(16'h61F2,4);
TASK_PP(16'h61F3,4);
TASK_PP(16'h61F4,4);
TASK_PP(16'h61F5,4);
TASK_PP(16'h61F6,4);
TASK_PP(16'h61F7,4);
TASK_PP(16'h61F8,4);
TASK_PP(16'h61F9,4);
TASK_PP(16'h61FA,4);
TASK_PP(16'h61FB,4);
TASK_PP(16'h61FC,4);
TASK_PP(16'h61FD,4);
TASK_PP(16'h61FE,4);
TASK_PP(16'h61FF,4);
TASK_PP(16'h6200,4);
TASK_PP(16'h6201,4);
TASK_PP(16'h6202,4);
TASK_PP(16'h6203,4);
TASK_PP(16'h6204,4);
TASK_PP(16'h6205,4);
TASK_PP(16'h6206,4);
TASK_PP(16'h6207,4);
TASK_PP(16'h6208,4);
TASK_PP(16'h6209,4);
TASK_PP(16'h620A,4);
TASK_PP(16'h620B,4);
TASK_PP(16'h620C,4);
TASK_PP(16'h620D,4);
TASK_PP(16'h620E,4);
TASK_PP(16'h620F,4);
TASK_PP(16'h6210,4);
TASK_PP(16'h6211,4);
TASK_PP(16'h6212,4);
TASK_PP(16'h6213,4);
TASK_PP(16'h6214,4);
TASK_PP(16'h6215,4);
TASK_PP(16'h6216,4);
TASK_PP(16'h6217,4);
TASK_PP(16'h6218,4);
TASK_PP(16'h6219,4);
TASK_PP(16'h621A,4);
TASK_PP(16'h621B,4);
TASK_PP(16'h621C,4);
TASK_PP(16'h621D,4);
TASK_PP(16'h621E,4);
TASK_PP(16'h621F,4);
TASK_PP(16'h6220,4);
TASK_PP(16'h6221,4);
TASK_PP(16'h6222,4);
TASK_PP(16'h6223,4);
TASK_PP(16'h6224,4);
TASK_PP(16'h6225,4);
TASK_PP(16'h6226,4);
TASK_PP(16'h6227,4);
TASK_PP(16'h6228,4);
TASK_PP(16'h6229,4);
TASK_PP(16'h622A,4);
TASK_PP(16'h622B,4);
TASK_PP(16'h622C,4);
TASK_PP(16'h622D,4);
TASK_PP(16'h622E,4);
TASK_PP(16'h622F,4);
TASK_PP(16'h6230,4);
TASK_PP(16'h6231,4);
TASK_PP(16'h6232,4);
TASK_PP(16'h6233,4);
TASK_PP(16'h6234,4);
TASK_PP(16'h6235,4);
TASK_PP(16'h6236,4);
TASK_PP(16'h6237,4);
TASK_PP(16'h6238,4);
TASK_PP(16'h6239,4);
TASK_PP(16'h623A,4);
TASK_PP(16'h623B,4);
TASK_PP(16'h623C,4);
TASK_PP(16'h623D,4);
TASK_PP(16'h623E,4);
TASK_PP(16'h623F,4);
TASK_PP(16'h6240,4);
TASK_PP(16'h6241,4);
TASK_PP(16'h6242,4);
TASK_PP(16'h6243,4);
TASK_PP(16'h6244,4);
TASK_PP(16'h6245,4);
TASK_PP(16'h6246,4);
TASK_PP(16'h6247,4);
TASK_PP(16'h6248,4);
TASK_PP(16'h6249,4);
TASK_PP(16'h624A,4);
TASK_PP(16'h624B,4);
TASK_PP(16'h624C,4);
TASK_PP(16'h624D,4);
TASK_PP(16'h624E,4);
TASK_PP(16'h624F,4);
TASK_PP(16'h6250,4);
TASK_PP(16'h6251,4);
TASK_PP(16'h6252,4);
TASK_PP(16'h6253,4);
TASK_PP(16'h6254,4);
TASK_PP(16'h6255,4);
TASK_PP(16'h6256,4);
TASK_PP(16'h6257,4);
TASK_PP(16'h6258,4);
TASK_PP(16'h6259,4);
TASK_PP(16'h625A,4);
TASK_PP(16'h625B,4);
TASK_PP(16'h625C,4);
TASK_PP(16'h625D,4);
TASK_PP(16'h625E,4);
TASK_PP(16'h625F,4);
TASK_PP(16'h6260,4);
TASK_PP(16'h6261,4);
TASK_PP(16'h6262,4);
TASK_PP(16'h6263,4);
TASK_PP(16'h6264,4);
TASK_PP(16'h6265,4);
TASK_PP(16'h6266,4);
TASK_PP(16'h6267,4);
TASK_PP(16'h6268,4);
TASK_PP(16'h6269,4);
TASK_PP(16'h626A,4);
TASK_PP(16'h626B,4);
TASK_PP(16'h626C,4);
TASK_PP(16'h626D,4);
TASK_PP(16'h626E,4);
TASK_PP(16'h626F,4);
TASK_PP(16'h6270,4);
TASK_PP(16'h6271,4);
TASK_PP(16'h6272,4);
TASK_PP(16'h6273,4);
TASK_PP(16'h6274,4);
TASK_PP(16'h6275,4);
TASK_PP(16'h6276,4);
TASK_PP(16'h6277,4);
TASK_PP(16'h6278,4);
TASK_PP(16'h6279,4);
TASK_PP(16'h627A,4);
TASK_PP(16'h627B,4);
TASK_PP(16'h627C,4);
TASK_PP(16'h627D,4);
TASK_PP(16'h627E,4);
TASK_PP(16'h627F,4);
TASK_PP(16'h6280,4);
TASK_PP(16'h6281,4);
TASK_PP(16'h6282,4);
TASK_PP(16'h6283,4);
TASK_PP(16'h6284,4);
TASK_PP(16'h6285,4);
TASK_PP(16'h6286,4);
TASK_PP(16'h6287,4);
TASK_PP(16'h6288,4);
TASK_PP(16'h6289,4);
TASK_PP(16'h628A,4);
TASK_PP(16'h628B,4);
TASK_PP(16'h628C,4);
TASK_PP(16'h628D,4);
TASK_PP(16'h628E,4);
TASK_PP(16'h628F,4);
TASK_PP(16'h6290,4);
TASK_PP(16'h6291,4);
TASK_PP(16'h6292,4);
TASK_PP(16'h6293,4);
TASK_PP(16'h6294,4);
TASK_PP(16'h6295,4);
TASK_PP(16'h6296,4);
TASK_PP(16'h6297,4);
TASK_PP(16'h6298,4);
TASK_PP(16'h6299,4);
TASK_PP(16'h629A,4);
TASK_PP(16'h629B,4);
TASK_PP(16'h629C,4);
TASK_PP(16'h629D,4);
TASK_PP(16'h629E,4);
TASK_PP(16'h629F,4);
TASK_PP(16'h62A0,4);
TASK_PP(16'h62A1,4);
TASK_PP(16'h62A2,4);
TASK_PP(16'h62A3,4);
TASK_PP(16'h62A4,4);
TASK_PP(16'h62A5,4);
TASK_PP(16'h62A6,4);
TASK_PP(16'h62A7,4);
TASK_PP(16'h62A8,4);
TASK_PP(16'h62A9,4);
TASK_PP(16'h62AA,4);
TASK_PP(16'h62AB,4);
TASK_PP(16'h62AC,4);
TASK_PP(16'h62AD,4);
TASK_PP(16'h62AE,4);
TASK_PP(16'h62AF,4);
TASK_PP(16'h62B0,4);
TASK_PP(16'h62B1,4);
TASK_PP(16'h62B2,4);
TASK_PP(16'h62B3,4);
TASK_PP(16'h62B4,4);
TASK_PP(16'h62B5,4);
TASK_PP(16'h62B6,4);
TASK_PP(16'h62B7,4);
TASK_PP(16'h62B8,4);
TASK_PP(16'h62B9,4);
TASK_PP(16'h62BA,4);
TASK_PP(16'h62BB,4);
TASK_PP(16'h62BC,4);
TASK_PP(16'h62BD,4);
TASK_PP(16'h62BE,4);
TASK_PP(16'h62BF,4);
TASK_PP(16'h62C0,4);
TASK_PP(16'h62C1,4);
TASK_PP(16'h62C2,4);
TASK_PP(16'h62C3,4);
TASK_PP(16'h62C4,4);
TASK_PP(16'h62C5,4);
TASK_PP(16'h62C6,4);
TASK_PP(16'h62C7,4);
TASK_PP(16'h62C8,4);
TASK_PP(16'h62C9,4);
TASK_PP(16'h62CA,4);
TASK_PP(16'h62CB,4);
TASK_PP(16'h62CC,4);
TASK_PP(16'h62CD,4);
TASK_PP(16'h62CE,4);
TASK_PP(16'h62CF,4);
TASK_PP(16'h62D0,4);
TASK_PP(16'h62D1,4);
TASK_PP(16'h62D2,4);
TASK_PP(16'h62D3,4);
TASK_PP(16'h62D4,4);
TASK_PP(16'h62D5,4);
TASK_PP(16'h62D6,4);
TASK_PP(16'h62D7,4);
TASK_PP(16'h62D8,4);
TASK_PP(16'h62D9,4);
TASK_PP(16'h62DA,4);
TASK_PP(16'h62DB,4);
TASK_PP(16'h62DC,4);
TASK_PP(16'h62DD,4);
TASK_PP(16'h62DE,4);
TASK_PP(16'h62DF,4);
TASK_PP(16'h62E0,4);
TASK_PP(16'h62E1,4);
TASK_PP(16'h62E2,4);
TASK_PP(16'h62E3,4);
TASK_PP(16'h62E4,4);
TASK_PP(16'h62E5,4);
TASK_PP(16'h62E6,4);
TASK_PP(16'h62E7,4);
TASK_PP(16'h62E8,4);
TASK_PP(16'h62E9,4);
TASK_PP(16'h62EA,4);
TASK_PP(16'h62EB,4);
TASK_PP(16'h62EC,4);
TASK_PP(16'h62ED,4);
TASK_PP(16'h62EE,4);
TASK_PP(16'h62EF,4);
TASK_PP(16'h62F0,4);
TASK_PP(16'h62F1,4);
TASK_PP(16'h62F2,4);
TASK_PP(16'h62F3,4);
TASK_PP(16'h62F4,4);
TASK_PP(16'h62F5,4);
TASK_PP(16'h62F6,4);
TASK_PP(16'h62F7,4);
TASK_PP(16'h62F8,4);
TASK_PP(16'h62F9,4);
TASK_PP(16'h62FA,4);
TASK_PP(16'h62FB,4);
TASK_PP(16'h62FC,4);
TASK_PP(16'h62FD,4);
TASK_PP(16'h62FE,4);
TASK_PP(16'h62FF,4);
TASK_PP(16'h6300,4);
TASK_PP(16'h6301,4);
TASK_PP(16'h6302,4);
TASK_PP(16'h6303,4);
TASK_PP(16'h6304,4);
TASK_PP(16'h6305,4);
TASK_PP(16'h6306,4);
TASK_PP(16'h6307,4);
TASK_PP(16'h6308,4);
TASK_PP(16'h6309,4);
TASK_PP(16'h630A,4);
TASK_PP(16'h630B,4);
TASK_PP(16'h630C,4);
TASK_PP(16'h630D,4);
TASK_PP(16'h630E,4);
TASK_PP(16'h630F,4);
TASK_PP(16'h6310,4);
TASK_PP(16'h6311,4);
TASK_PP(16'h6312,4);
TASK_PP(16'h6313,4);
TASK_PP(16'h6314,4);
TASK_PP(16'h6315,4);
TASK_PP(16'h6316,4);
TASK_PP(16'h6317,4);
TASK_PP(16'h6318,4);
TASK_PP(16'h6319,4);
TASK_PP(16'h631A,4);
TASK_PP(16'h631B,4);
TASK_PP(16'h631C,4);
TASK_PP(16'h631D,4);
TASK_PP(16'h631E,4);
TASK_PP(16'h631F,4);
TASK_PP(16'h6320,4);
TASK_PP(16'h6321,4);
TASK_PP(16'h6322,4);
TASK_PP(16'h6323,4);
TASK_PP(16'h6324,4);
TASK_PP(16'h6325,4);
TASK_PP(16'h6326,4);
TASK_PP(16'h6327,4);
TASK_PP(16'h6328,4);
TASK_PP(16'h6329,4);
TASK_PP(16'h632A,4);
TASK_PP(16'h632B,4);
TASK_PP(16'h632C,4);
TASK_PP(16'h632D,4);
TASK_PP(16'h632E,4);
TASK_PP(16'h632F,4);
TASK_PP(16'h6330,4);
TASK_PP(16'h6331,4);
TASK_PP(16'h6332,4);
TASK_PP(16'h6333,4);
TASK_PP(16'h6334,4);
TASK_PP(16'h6335,4);
TASK_PP(16'h6336,4);
TASK_PP(16'h6337,4);
TASK_PP(16'h6338,4);
TASK_PP(16'h6339,4);
TASK_PP(16'h633A,4);
TASK_PP(16'h633B,4);
TASK_PP(16'h633C,4);
TASK_PP(16'h633D,4);
TASK_PP(16'h633E,4);
TASK_PP(16'h633F,4);
TASK_PP(16'h6340,4);
TASK_PP(16'h6341,4);
TASK_PP(16'h6342,4);
TASK_PP(16'h6343,4);
TASK_PP(16'h6344,4);
TASK_PP(16'h6345,4);
TASK_PP(16'h6346,4);
TASK_PP(16'h6347,4);
TASK_PP(16'h6348,4);
TASK_PP(16'h6349,4);
TASK_PP(16'h634A,4);
TASK_PP(16'h634B,4);
TASK_PP(16'h634C,4);
TASK_PP(16'h634D,4);
TASK_PP(16'h634E,4);
TASK_PP(16'h634F,4);
TASK_PP(16'h6350,4);
TASK_PP(16'h6351,4);
TASK_PP(16'h6352,4);
TASK_PP(16'h6353,4);
TASK_PP(16'h6354,4);
TASK_PP(16'h6355,4);
TASK_PP(16'h6356,4);
TASK_PP(16'h6357,4);
TASK_PP(16'h6358,4);
TASK_PP(16'h6359,4);
TASK_PP(16'h635A,4);
TASK_PP(16'h635B,4);
TASK_PP(16'h635C,4);
TASK_PP(16'h635D,4);
TASK_PP(16'h635E,4);
TASK_PP(16'h635F,4);
TASK_PP(16'h6360,4);
TASK_PP(16'h6361,4);
TASK_PP(16'h6362,4);
TASK_PP(16'h6363,4);
TASK_PP(16'h6364,4);
TASK_PP(16'h6365,4);
TASK_PP(16'h6366,4);
TASK_PP(16'h6367,4);
TASK_PP(16'h6368,4);
TASK_PP(16'h6369,4);
TASK_PP(16'h636A,4);
TASK_PP(16'h636B,4);
TASK_PP(16'h636C,4);
TASK_PP(16'h636D,4);
TASK_PP(16'h636E,4);
TASK_PP(16'h636F,4);
TASK_PP(16'h6370,4);
TASK_PP(16'h6371,4);
TASK_PP(16'h6372,4);
TASK_PP(16'h6373,4);
TASK_PP(16'h6374,4);
TASK_PP(16'h6375,4);
TASK_PP(16'h6376,4);
TASK_PP(16'h6377,4);
TASK_PP(16'h6378,4);
TASK_PP(16'h6379,4);
TASK_PP(16'h637A,4);
TASK_PP(16'h637B,4);
TASK_PP(16'h637C,4);
TASK_PP(16'h637D,4);
TASK_PP(16'h637E,4);
TASK_PP(16'h637F,4);
TASK_PP(16'h6380,4);
TASK_PP(16'h6381,4);
TASK_PP(16'h6382,4);
TASK_PP(16'h6383,4);
TASK_PP(16'h6384,4);
TASK_PP(16'h6385,4);
TASK_PP(16'h6386,4);
TASK_PP(16'h6387,4);
TASK_PP(16'h6388,4);
TASK_PP(16'h6389,4);
TASK_PP(16'h638A,4);
TASK_PP(16'h638B,4);
TASK_PP(16'h638C,4);
TASK_PP(16'h638D,4);
TASK_PP(16'h638E,4);
TASK_PP(16'h638F,4);
TASK_PP(16'h6390,4);
TASK_PP(16'h6391,4);
TASK_PP(16'h6392,4);
TASK_PP(16'h6393,4);
TASK_PP(16'h6394,4);
TASK_PP(16'h6395,4);
TASK_PP(16'h6396,4);
TASK_PP(16'h6397,4);
TASK_PP(16'h6398,4);
TASK_PP(16'h6399,4);
TASK_PP(16'h639A,4);
TASK_PP(16'h639B,4);
TASK_PP(16'h639C,4);
TASK_PP(16'h639D,4);
TASK_PP(16'h639E,4);
TASK_PP(16'h639F,4);
TASK_PP(16'h63A0,4);
TASK_PP(16'h63A1,4);
TASK_PP(16'h63A2,4);
TASK_PP(16'h63A3,4);
TASK_PP(16'h63A4,4);
TASK_PP(16'h63A5,4);
TASK_PP(16'h63A6,4);
TASK_PP(16'h63A7,4);
TASK_PP(16'h63A8,4);
TASK_PP(16'h63A9,4);
TASK_PP(16'h63AA,4);
TASK_PP(16'h63AB,4);
TASK_PP(16'h63AC,4);
TASK_PP(16'h63AD,4);
TASK_PP(16'h63AE,4);
TASK_PP(16'h63AF,4);
TASK_PP(16'h63B0,4);
TASK_PP(16'h63B1,4);
TASK_PP(16'h63B2,4);
TASK_PP(16'h63B3,4);
TASK_PP(16'h63B4,4);
TASK_PP(16'h63B5,4);
TASK_PP(16'h63B6,4);
TASK_PP(16'h63B7,4);
TASK_PP(16'h63B8,4);
TASK_PP(16'h63B9,4);
TASK_PP(16'h63BA,4);
TASK_PP(16'h63BB,4);
TASK_PP(16'h63BC,4);
TASK_PP(16'h63BD,4);
TASK_PP(16'h63BE,4);
TASK_PP(16'h63BF,4);
TASK_PP(16'h63C0,4);
TASK_PP(16'h63C1,4);
TASK_PP(16'h63C2,4);
TASK_PP(16'h63C3,4);
TASK_PP(16'h63C4,4);
TASK_PP(16'h63C5,4);
TASK_PP(16'h63C6,4);
TASK_PP(16'h63C7,4);
TASK_PP(16'h63C8,4);
TASK_PP(16'h63C9,4);
TASK_PP(16'h63CA,4);
TASK_PP(16'h63CB,4);
TASK_PP(16'h63CC,4);
TASK_PP(16'h63CD,4);
TASK_PP(16'h63CE,4);
TASK_PP(16'h63CF,4);
TASK_PP(16'h63D0,4);
TASK_PP(16'h63D1,4);
TASK_PP(16'h63D2,4);
TASK_PP(16'h63D3,4);
TASK_PP(16'h63D4,4);
TASK_PP(16'h63D5,4);
TASK_PP(16'h63D6,4);
TASK_PP(16'h63D7,4);
TASK_PP(16'h63D8,4);
TASK_PP(16'h63D9,4);
TASK_PP(16'h63DA,4);
TASK_PP(16'h63DB,4);
TASK_PP(16'h63DC,4);
TASK_PP(16'h63DD,4);
TASK_PP(16'h63DE,4);
TASK_PP(16'h63DF,4);
TASK_PP(16'h63E0,4);
TASK_PP(16'h63E1,4);
TASK_PP(16'h63E2,4);
TASK_PP(16'h63E3,4);
TASK_PP(16'h63E4,4);
TASK_PP(16'h63E5,4);
TASK_PP(16'h63E6,4);
TASK_PP(16'h63E7,4);
TASK_PP(16'h63E8,4);
TASK_PP(16'h63E9,4);
TASK_PP(16'h63EA,4);
TASK_PP(16'h63EB,4);
TASK_PP(16'h63EC,4);
TASK_PP(16'h63ED,4);
TASK_PP(16'h63EE,4);
TASK_PP(16'h63EF,4);
TASK_PP(16'h63F0,4);
TASK_PP(16'h63F1,4);
TASK_PP(16'h63F2,4);
TASK_PP(16'h63F3,4);
TASK_PP(16'h63F4,4);
TASK_PP(16'h63F5,4);
TASK_PP(16'h63F6,4);
TASK_PP(16'h63F7,4);
TASK_PP(16'h63F8,4);
TASK_PP(16'h63F9,4);
TASK_PP(16'h63FA,4);
TASK_PP(16'h63FB,4);
TASK_PP(16'h63FC,4);
TASK_PP(16'h63FD,4);
TASK_PP(16'h63FE,4);
TASK_PP(16'h63FF,4);
TASK_PP(16'h6400,4);
TASK_PP(16'h6401,4);
TASK_PP(16'h6402,4);
TASK_PP(16'h6403,4);
TASK_PP(16'h6404,4);
TASK_PP(16'h6405,4);
TASK_PP(16'h6406,4);
TASK_PP(16'h6407,4);
TASK_PP(16'h6408,4);
TASK_PP(16'h6409,4);
TASK_PP(16'h640A,4);
TASK_PP(16'h640B,4);
TASK_PP(16'h640C,4);
TASK_PP(16'h640D,4);
TASK_PP(16'h640E,4);
TASK_PP(16'h640F,4);
TASK_PP(16'h6410,4);
TASK_PP(16'h6411,4);
TASK_PP(16'h6412,4);
TASK_PP(16'h6413,4);
TASK_PP(16'h6414,4);
TASK_PP(16'h6415,4);
TASK_PP(16'h6416,4);
TASK_PP(16'h6417,4);
TASK_PP(16'h6418,4);
TASK_PP(16'h6419,4);
TASK_PP(16'h641A,4);
TASK_PP(16'h641B,4);
TASK_PP(16'h641C,4);
TASK_PP(16'h641D,4);
TASK_PP(16'h641E,4);
TASK_PP(16'h641F,4);
TASK_PP(16'h6420,4);
TASK_PP(16'h6421,4);
TASK_PP(16'h6422,4);
TASK_PP(16'h6423,4);
TASK_PP(16'h6424,4);
TASK_PP(16'h6425,4);
TASK_PP(16'h6426,4);
TASK_PP(16'h6427,4);
TASK_PP(16'h6428,4);
TASK_PP(16'h6429,4);
TASK_PP(16'h642A,4);
TASK_PP(16'h642B,4);
TASK_PP(16'h642C,4);
TASK_PP(16'h642D,4);
TASK_PP(16'h642E,4);
TASK_PP(16'h642F,4);
TASK_PP(16'h6430,4);
TASK_PP(16'h6431,4);
TASK_PP(16'h6432,4);
TASK_PP(16'h6433,4);
TASK_PP(16'h6434,4);
TASK_PP(16'h6435,4);
TASK_PP(16'h6436,4);
TASK_PP(16'h6437,4);
TASK_PP(16'h6438,4);
TASK_PP(16'h6439,4);
TASK_PP(16'h643A,4);
TASK_PP(16'h643B,4);
TASK_PP(16'h643C,4);
TASK_PP(16'h643D,4);
TASK_PP(16'h643E,4);
TASK_PP(16'h643F,4);
TASK_PP(16'h6440,4);
TASK_PP(16'h6441,4);
TASK_PP(16'h6442,4);
TASK_PP(16'h6443,4);
TASK_PP(16'h6444,4);
TASK_PP(16'h6445,4);
TASK_PP(16'h6446,4);
TASK_PP(16'h6447,4);
TASK_PP(16'h6448,4);
TASK_PP(16'h6449,4);
TASK_PP(16'h644A,4);
TASK_PP(16'h644B,4);
TASK_PP(16'h644C,4);
TASK_PP(16'h644D,4);
TASK_PP(16'h644E,4);
TASK_PP(16'h644F,4);
TASK_PP(16'h6450,4);
TASK_PP(16'h6451,4);
TASK_PP(16'h6452,4);
TASK_PP(16'h6453,4);
TASK_PP(16'h6454,4);
TASK_PP(16'h6455,4);
TASK_PP(16'h6456,4);
TASK_PP(16'h6457,4);
TASK_PP(16'h6458,4);
TASK_PP(16'h6459,4);
TASK_PP(16'h645A,4);
TASK_PP(16'h645B,4);
TASK_PP(16'h645C,4);
TASK_PP(16'h645D,4);
TASK_PP(16'h645E,4);
TASK_PP(16'h645F,4);
TASK_PP(16'h6460,4);
TASK_PP(16'h6461,4);
TASK_PP(16'h6462,4);
TASK_PP(16'h6463,4);
TASK_PP(16'h6464,4);
TASK_PP(16'h6465,4);
TASK_PP(16'h6466,4);
TASK_PP(16'h6467,4);
TASK_PP(16'h6468,4);
TASK_PP(16'h6469,4);
TASK_PP(16'h646A,4);
TASK_PP(16'h646B,4);
TASK_PP(16'h646C,4);
TASK_PP(16'h646D,4);
TASK_PP(16'h646E,4);
TASK_PP(16'h646F,4);
TASK_PP(16'h6470,4);
TASK_PP(16'h6471,4);
TASK_PP(16'h6472,4);
TASK_PP(16'h6473,4);
TASK_PP(16'h6474,4);
TASK_PP(16'h6475,4);
TASK_PP(16'h6476,4);
TASK_PP(16'h6477,4);
TASK_PP(16'h6478,4);
TASK_PP(16'h6479,4);
TASK_PP(16'h647A,4);
TASK_PP(16'h647B,4);
TASK_PP(16'h647C,4);
TASK_PP(16'h647D,4);
TASK_PP(16'h647E,4);
TASK_PP(16'h647F,4);
TASK_PP(16'h6480,4);
TASK_PP(16'h6481,4);
TASK_PP(16'h6482,4);
TASK_PP(16'h6483,4);
TASK_PP(16'h6484,4);
TASK_PP(16'h6485,4);
TASK_PP(16'h6486,4);
TASK_PP(16'h6487,4);
TASK_PP(16'h6488,4);
TASK_PP(16'h6489,4);
TASK_PP(16'h648A,4);
TASK_PP(16'h648B,4);
TASK_PP(16'h648C,4);
TASK_PP(16'h648D,4);
TASK_PP(16'h648E,4);
TASK_PP(16'h648F,4);
TASK_PP(16'h6490,4);
TASK_PP(16'h6491,4);
TASK_PP(16'h6492,4);
TASK_PP(16'h6493,4);
TASK_PP(16'h6494,4);
TASK_PP(16'h6495,4);
TASK_PP(16'h6496,4);
TASK_PP(16'h6497,4);
TASK_PP(16'h6498,4);
TASK_PP(16'h6499,4);
TASK_PP(16'h649A,4);
TASK_PP(16'h649B,4);
TASK_PP(16'h649C,4);
TASK_PP(16'h649D,4);
TASK_PP(16'h649E,4);
TASK_PP(16'h649F,4);
TASK_PP(16'h64A0,4);
TASK_PP(16'h64A1,4);
TASK_PP(16'h64A2,4);
TASK_PP(16'h64A3,4);
TASK_PP(16'h64A4,4);
TASK_PP(16'h64A5,4);
TASK_PP(16'h64A6,4);
TASK_PP(16'h64A7,4);
TASK_PP(16'h64A8,4);
TASK_PP(16'h64A9,4);
TASK_PP(16'h64AA,4);
TASK_PP(16'h64AB,4);
TASK_PP(16'h64AC,4);
TASK_PP(16'h64AD,4);
TASK_PP(16'h64AE,4);
TASK_PP(16'h64AF,4);
TASK_PP(16'h64B0,4);
TASK_PP(16'h64B1,4);
TASK_PP(16'h64B2,4);
TASK_PP(16'h64B3,4);
TASK_PP(16'h64B4,4);
TASK_PP(16'h64B5,4);
TASK_PP(16'h64B6,4);
TASK_PP(16'h64B7,4);
TASK_PP(16'h64B8,4);
TASK_PP(16'h64B9,4);
TASK_PP(16'h64BA,4);
TASK_PP(16'h64BB,4);
TASK_PP(16'h64BC,4);
TASK_PP(16'h64BD,4);
TASK_PP(16'h64BE,4);
TASK_PP(16'h64BF,4);
TASK_PP(16'h64C0,4);
TASK_PP(16'h64C1,4);
TASK_PP(16'h64C2,4);
TASK_PP(16'h64C3,4);
TASK_PP(16'h64C4,4);
TASK_PP(16'h64C5,4);
TASK_PP(16'h64C6,4);
TASK_PP(16'h64C7,4);
TASK_PP(16'h64C8,4);
TASK_PP(16'h64C9,4);
TASK_PP(16'h64CA,4);
TASK_PP(16'h64CB,4);
TASK_PP(16'h64CC,4);
TASK_PP(16'h64CD,4);
TASK_PP(16'h64CE,4);
TASK_PP(16'h64CF,4);
TASK_PP(16'h64D0,4);
TASK_PP(16'h64D1,4);
TASK_PP(16'h64D2,4);
TASK_PP(16'h64D3,4);
TASK_PP(16'h64D4,4);
TASK_PP(16'h64D5,4);
TASK_PP(16'h64D6,4);
TASK_PP(16'h64D7,4);
TASK_PP(16'h64D8,4);
TASK_PP(16'h64D9,4);
TASK_PP(16'h64DA,4);
TASK_PP(16'h64DB,4);
TASK_PP(16'h64DC,4);
TASK_PP(16'h64DD,4);
TASK_PP(16'h64DE,4);
TASK_PP(16'h64DF,4);
TASK_PP(16'h64E0,4);
TASK_PP(16'h64E1,4);
TASK_PP(16'h64E2,4);
TASK_PP(16'h64E3,4);
TASK_PP(16'h64E4,4);
TASK_PP(16'h64E5,4);
TASK_PP(16'h64E6,4);
TASK_PP(16'h64E7,4);
TASK_PP(16'h64E8,4);
TASK_PP(16'h64E9,4);
TASK_PP(16'h64EA,4);
TASK_PP(16'h64EB,4);
TASK_PP(16'h64EC,4);
TASK_PP(16'h64ED,4);
TASK_PP(16'h64EE,4);
TASK_PP(16'h64EF,4);
TASK_PP(16'h64F0,4);
TASK_PP(16'h64F1,4);
TASK_PP(16'h64F2,4);
TASK_PP(16'h64F3,4);
TASK_PP(16'h64F4,4);
TASK_PP(16'h64F5,4);
TASK_PP(16'h64F6,4);
TASK_PP(16'h64F7,4);
TASK_PP(16'h64F8,4);
TASK_PP(16'h64F9,4);
TASK_PP(16'h64FA,4);
TASK_PP(16'h64FB,4);
TASK_PP(16'h64FC,4);
TASK_PP(16'h64FD,4);
TASK_PP(16'h64FE,4);
TASK_PP(16'h64FF,4);
TASK_PP(16'h6500,4);
TASK_PP(16'h6501,4);
TASK_PP(16'h6502,4);
TASK_PP(16'h6503,4);
TASK_PP(16'h6504,4);
TASK_PP(16'h6505,4);
TASK_PP(16'h6506,4);
TASK_PP(16'h6507,4);
TASK_PP(16'h6508,4);
TASK_PP(16'h6509,4);
TASK_PP(16'h650A,4);
TASK_PP(16'h650B,4);
TASK_PP(16'h650C,4);
TASK_PP(16'h650D,4);
TASK_PP(16'h650E,4);
TASK_PP(16'h650F,4);
TASK_PP(16'h6510,4);
TASK_PP(16'h6511,4);
TASK_PP(16'h6512,4);
TASK_PP(16'h6513,4);
TASK_PP(16'h6514,4);
TASK_PP(16'h6515,4);
TASK_PP(16'h6516,4);
TASK_PP(16'h6517,4);
TASK_PP(16'h6518,4);
TASK_PP(16'h6519,4);
TASK_PP(16'h651A,4);
TASK_PP(16'h651B,4);
TASK_PP(16'h651C,4);
TASK_PP(16'h651D,4);
TASK_PP(16'h651E,4);
TASK_PP(16'h651F,4);
TASK_PP(16'h6520,4);
TASK_PP(16'h6521,4);
TASK_PP(16'h6522,4);
TASK_PP(16'h6523,4);
TASK_PP(16'h6524,4);
TASK_PP(16'h6525,4);
TASK_PP(16'h6526,4);
TASK_PP(16'h6527,4);
TASK_PP(16'h6528,4);
TASK_PP(16'h6529,4);
TASK_PP(16'h652A,4);
TASK_PP(16'h652B,4);
TASK_PP(16'h652C,4);
TASK_PP(16'h652D,4);
TASK_PP(16'h652E,4);
TASK_PP(16'h652F,4);
TASK_PP(16'h6530,4);
TASK_PP(16'h6531,4);
TASK_PP(16'h6532,4);
TASK_PP(16'h6533,4);
TASK_PP(16'h6534,4);
TASK_PP(16'h6535,4);
TASK_PP(16'h6536,4);
TASK_PP(16'h6537,4);
TASK_PP(16'h6538,4);
TASK_PP(16'h6539,4);
TASK_PP(16'h653A,4);
TASK_PP(16'h653B,4);
TASK_PP(16'h653C,4);
TASK_PP(16'h653D,4);
TASK_PP(16'h653E,4);
TASK_PP(16'h653F,4);
TASK_PP(16'h6540,4);
TASK_PP(16'h6541,4);
TASK_PP(16'h6542,4);
TASK_PP(16'h6543,4);
TASK_PP(16'h6544,4);
TASK_PP(16'h6545,4);
TASK_PP(16'h6546,4);
TASK_PP(16'h6547,4);
TASK_PP(16'h6548,4);
TASK_PP(16'h6549,4);
TASK_PP(16'h654A,4);
TASK_PP(16'h654B,4);
TASK_PP(16'h654C,4);
TASK_PP(16'h654D,4);
TASK_PP(16'h654E,4);
TASK_PP(16'h654F,4);
TASK_PP(16'h6550,4);
TASK_PP(16'h6551,4);
TASK_PP(16'h6552,4);
TASK_PP(16'h6553,4);
TASK_PP(16'h6554,4);
TASK_PP(16'h6555,4);
TASK_PP(16'h6556,4);
TASK_PP(16'h6557,4);
TASK_PP(16'h6558,4);
TASK_PP(16'h6559,4);
TASK_PP(16'h655A,4);
TASK_PP(16'h655B,4);
TASK_PP(16'h655C,4);
TASK_PP(16'h655D,4);
TASK_PP(16'h655E,4);
TASK_PP(16'h655F,4);
TASK_PP(16'h6560,4);
TASK_PP(16'h6561,4);
TASK_PP(16'h6562,4);
TASK_PP(16'h6563,4);
TASK_PP(16'h6564,4);
TASK_PP(16'h6565,4);
TASK_PP(16'h6566,4);
TASK_PP(16'h6567,4);
TASK_PP(16'h6568,4);
TASK_PP(16'h6569,4);
TASK_PP(16'h656A,4);
TASK_PP(16'h656B,4);
TASK_PP(16'h656C,4);
TASK_PP(16'h656D,4);
TASK_PP(16'h656E,4);
TASK_PP(16'h656F,4);
TASK_PP(16'h6570,4);
TASK_PP(16'h6571,4);
TASK_PP(16'h6572,4);
TASK_PP(16'h6573,4);
TASK_PP(16'h6574,4);
TASK_PP(16'h6575,4);
TASK_PP(16'h6576,4);
TASK_PP(16'h6577,4);
TASK_PP(16'h6578,4);
TASK_PP(16'h6579,4);
TASK_PP(16'h657A,4);
TASK_PP(16'h657B,4);
TASK_PP(16'h657C,4);
TASK_PP(16'h657D,4);
TASK_PP(16'h657E,4);
TASK_PP(16'h657F,4);
TASK_PP(16'h6580,4);
TASK_PP(16'h6581,4);
TASK_PP(16'h6582,4);
TASK_PP(16'h6583,4);
TASK_PP(16'h6584,4);
TASK_PP(16'h6585,4);
TASK_PP(16'h6586,4);
TASK_PP(16'h6587,4);
TASK_PP(16'h6588,4);
TASK_PP(16'h6589,4);
TASK_PP(16'h658A,4);
TASK_PP(16'h658B,4);
TASK_PP(16'h658C,4);
TASK_PP(16'h658D,4);
TASK_PP(16'h658E,4);
TASK_PP(16'h658F,4);
TASK_PP(16'h6590,4);
TASK_PP(16'h6591,4);
TASK_PP(16'h6592,4);
TASK_PP(16'h6593,4);
TASK_PP(16'h6594,4);
TASK_PP(16'h6595,4);
TASK_PP(16'h6596,4);
TASK_PP(16'h6597,4);
TASK_PP(16'h6598,4);
TASK_PP(16'h6599,4);
TASK_PP(16'h659A,4);
TASK_PP(16'h659B,4);
TASK_PP(16'h659C,4);
TASK_PP(16'h659D,4);
TASK_PP(16'h659E,4);
TASK_PP(16'h659F,4);
TASK_PP(16'h65A0,4);
TASK_PP(16'h65A1,4);
TASK_PP(16'h65A2,4);
TASK_PP(16'h65A3,4);
TASK_PP(16'h65A4,4);
TASK_PP(16'h65A5,4);
TASK_PP(16'h65A6,4);
TASK_PP(16'h65A7,4);
TASK_PP(16'h65A8,4);
TASK_PP(16'h65A9,4);
TASK_PP(16'h65AA,4);
TASK_PP(16'h65AB,4);
TASK_PP(16'h65AC,4);
TASK_PP(16'h65AD,4);
TASK_PP(16'h65AE,4);
TASK_PP(16'h65AF,4);
TASK_PP(16'h65B0,4);
TASK_PP(16'h65B1,4);
TASK_PP(16'h65B2,4);
TASK_PP(16'h65B3,4);
TASK_PP(16'h65B4,4);
TASK_PP(16'h65B5,4);
TASK_PP(16'h65B6,4);
TASK_PP(16'h65B7,4);
TASK_PP(16'h65B8,4);
TASK_PP(16'h65B9,4);
TASK_PP(16'h65BA,4);
TASK_PP(16'h65BB,4);
TASK_PP(16'h65BC,4);
TASK_PP(16'h65BD,4);
TASK_PP(16'h65BE,4);
TASK_PP(16'h65BF,4);
TASK_PP(16'h65C0,4);
TASK_PP(16'h65C1,4);
TASK_PP(16'h65C2,4);
TASK_PP(16'h65C3,4);
TASK_PP(16'h65C4,4);
TASK_PP(16'h65C5,4);
TASK_PP(16'h65C6,4);
TASK_PP(16'h65C7,4);
TASK_PP(16'h65C8,4);
TASK_PP(16'h65C9,4);
TASK_PP(16'h65CA,4);
TASK_PP(16'h65CB,4);
TASK_PP(16'h65CC,4);
TASK_PP(16'h65CD,4);
TASK_PP(16'h65CE,4);
TASK_PP(16'h65CF,4);
TASK_PP(16'h65D0,4);
TASK_PP(16'h65D1,4);
TASK_PP(16'h65D2,4);
TASK_PP(16'h65D3,4);
TASK_PP(16'h65D4,4);
TASK_PP(16'h65D5,4);
TASK_PP(16'h65D6,4);
TASK_PP(16'h65D7,4);
TASK_PP(16'h65D8,4);
TASK_PP(16'h65D9,4);
TASK_PP(16'h65DA,4);
TASK_PP(16'h65DB,4);
TASK_PP(16'h65DC,4);
TASK_PP(16'h65DD,4);
TASK_PP(16'h65DE,4);
TASK_PP(16'h65DF,4);
TASK_PP(16'h65E0,4);
TASK_PP(16'h65E1,4);
TASK_PP(16'h65E2,4);
TASK_PP(16'h65E3,4);
TASK_PP(16'h65E4,4);
TASK_PP(16'h65E5,4);
TASK_PP(16'h65E6,4);
TASK_PP(16'h65E7,4);
TASK_PP(16'h65E8,4);
TASK_PP(16'h65E9,4);
TASK_PP(16'h65EA,4);
TASK_PP(16'h65EB,4);
TASK_PP(16'h65EC,4);
TASK_PP(16'h65ED,4);
TASK_PP(16'h65EE,4);
TASK_PP(16'h65EF,4);
TASK_PP(16'h65F0,4);
TASK_PP(16'h65F1,4);
TASK_PP(16'h65F2,4);
TASK_PP(16'h65F3,4);
TASK_PP(16'h65F4,4);
TASK_PP(16'h65F5,4);
TASK_PP(16'h65F6,4);
TASK_PP(16'h65F7,4);
TASK_PP(16'h65F8,4);
TASK_PP(16'h65F9,4);
TASK_PP(16'h65FA,4);
TASK_PP(16'h65FB,4);
TASK_PP(16'h65FC,4);
TASK_PP(16'h65FD,4);
TASK_PP(16'h65FE,4);
TASK_PP(16'h65FF,4);
TASK_PP(16'h6600,4);
TASK_PP(16'h6601,4);
TASK_PP(16'h6602,4);
TASK_PP(16'h6603,4);
TASK_PP(16'h6604,4);
TASK_PP(16'h6605,4);
TASK_PP(16'h6606,4);
TASK_PP(16'h6607,4);
TASK_PP(16'h6608,4);
TASK_PP(16'h6609,4);
TASK_PP(16'h660A,4);
TASK_PP(16'h660B,4);
TASK_PP(16'h660C,4);
TASK_PP(16'h660D,4);
TASK_PP(16'h660E,4);
TASK_PP(16'h660F,4);
TASK_PP(16'h6610,4);
TASK_PP(16'h6611,4);
TASK_PP(16'h6612,4);
TASK_PP(16'h6613,4);
TASK_PP(16'h6614,4);
TASK_PP(16'h6615,4);
TASK_PP(16'h6616,4);
TASK_PP(16'h6617,4);
TASK_PP(16'h6618,4);
TASK_PP(16'h6619,4);
TASK_PP(16'h661A,4);
TASK_PP(16'h661B,4);
TASK_PP(16'h661C,4);
TASK_PP(16'h661D,4);
TASK_PP(16'h661E,4);
TASK_PP(16'h661F,4);
TASK_PP(16'h6620,4);
TASK_PP(16'h6621,4);
TASK_PP(16'h6622,4);
TASK_PP(16'h6623,4);
TASK_PP(16'h6624,4);
TASK_PP(16'h6625,4);
TASK_PP(16'h6626,4);
TASK_PP(16'h6627,4);
TASK_PP(16'h6628,4);
TASK_PP(16'h6629,4);
TASK_PP(16'h662A,4);
TASK_PP(16'h662B,4);
TASK_PP(16'h662C,4);
TASK_PP(16'h662D,4);
TASK_PP(16'h662E,4);
TASK_PP(16'h662F,4);
TASK_PP(16'h6630,4);
TASK_PP(16'h6631,4);
TASK_PP(16'h6632,4);
TASK_PP(16'h6633,4);
TASK_PP(16'h6634,4);
TASK_PP(16'h6635,4);
TASK_PP(16'h6636,4);
TASK_PP(16'h6637,4);
TASK_PP(16'h6638,4);
TASK_PP(16'h6639,4);
TASK_PP(16'h663A,4);
TASK_PP(16'h663B,4);
TASK_PP(16'h663C,4);
TASK_PP(16'h663D,4);
TASK_PP(16'h663E,4);
TASK_PP(16'h663F,4);
TASK_PP(16'h6640,4);
TASK_PP(16'h6641,4);
TASK_PP(16'h6642,4);
TASK_PP(16'h6643,4);
TASK_PP(16'h6644,4);
TASK_PP(16'h6645,4);
TASK_PP(16'h6646,4);
TASK_PP(16'h6647,4);
TASK_PP(16'h6648,4);
TASK_PP(16'h6649,4);
TASK_PP(16'h664A,4);
TASK_PP(16'h664B,4);
TASK_PP(16'h664C,4);
TASK_PP(16'h664D,4);
TASK_PP(16'h664E,4);
TASK_PP(16'h664F,4);
TASK_PP(16'h6650,4);
TASK_PP(16'h6651,4);
TASK_PP(16'h6652,4);
TASK_PP(16'h6653,4);
TASK_PP(16'h6654,4);
TASK_PP(16'h6655,4);
TASK_PP(16'h6656,4);
TASK_PP(16'h6657,4);
TASK_PP(16'h6658,4);
TASK_PP(16'h6659,4);
TASK_PP(16'h665A,4);
TASK_PP(16'h665B,4);
TASK_PP(16'h665C,4);
TASK_PP(16'h665D,4);
TASK_PP(16'h665E,4);
TASK_PP(16'h665F,4);
TASK_PP(16'h6660,4);
TASK_PP(16'h6661,4);
TASK_PP(16'h6662,4);
TASK_PP(16'h6663,4);
TASK_PP(16'h6664,4);
TASK_PP(16'h6665,4);
TASK_PP(16'h6666,4);
TASK_PP(16'h6667,4);
TASK_PP(16'h6668,4);
TASK_PP(16'h6669,4);
TASK_PP(16'h666A,4);
TASK_PP(16'h666B,4);
TASK_PP(16'h666C,4);
TASK_PP(16'h666D,4);
TASK_PP(16'h666E,4);
TASK_PP(16'h666F,4);
TASK_PP(16'h6670,4);
TASK_PP(16'h6671,4);
TASK_PP(16'h6672,4);
TASK_PP(16'h6673,4);
TASK_PP(16'h6674,4);
TASK_PP(16'h6675,4);
TASK_PP(16'h6676,4);
TASK_PP(16'h6677,4);
TASK_PP(16'h6678,4);
TASK_PP(16'h6679,4);
TASK_PP(16'h667A,4);
TASK_PP(16'h667B,4);
TASK_PP(16'h667C,4);
TASK_PP(16'h667D,4);
TASK_PP(16'h667E,4);
TASK_PP(16'h667F,4);
TASK_PP(16'h6680,4);
TASK_PP(16'h6681,4);
TASK_PP(16'h6682,4);
TASK_PP(16'h6683,4);
TASK_PP(16'h6684,4);
TASK_PP(16'h6685,4);
TASK_PP(16'h6686,4);
TASK_PP(16'h6687,4);
TASK_PP(16'h6688,4);
TASK_PP(16'h6689,4);
TASK_PP(16'h668A,4);
TASK_PP(16'h668B,4);
TASK_PP(16'h668C,4);
TASK_PP(16'h668D,4);
TASK_PP(16'h668E,4);
TASK_PP(16'h668F,4);
TASK_PP(16'h6690,4);
TASK_PP(16'h6691,4);
TASK_PP(16'h6692,4);
TASK_PP(16'h6693,4);
TASK_PP(16'h6694,4);
TASK_PP(16'h6695,4);
TASK_PP(16'h6696,4);
TASK_PP(16'h6697,4);
TASK_PP(16'h6698,4);
TASK_PP(16'h6699,4);
TASK_PP(16'h669A,4);
TASK_PP(16'h669B,4);
TASK_PP(16'h669C,4);
TASK_PP(16'h669D,4);
TASK_PP(16'h669E,4);
TASK_PP(16'h669F,4);
TASK_PP(16'h66A0,4);
TASK_PP(16'h66A1,4);
TASK_PP(16'h66A2,4);
TASK_PP(16'h66A3,4);
TASK_PP(16'h66A4,4);
TASK_PP(16'h66A5,4);
TASK_PP(16'h66A6,4);
TASK_PP(16'h66A7,4);
TASK_PP(16'h66A8,4);
TASK_PP(16'h66A9,4);
TASK_PP(16'h66AA,4);
TASK_PP(16'h66AB,4);
TASK_PP(16'h66AC,4);
TASK_PP(16'h66AD,4);
TASK_PP(16'h66AE,4);
TASK_PP(16'h66AF,4);
TASK_PP(16'h66B0,4);
TASK_PP(16'h66B1,4);
TASK_PP(16'h66B2,4);
TASK_PP(16'h66B3,4);
TASK_PP(16'h66B4,4);
TASK_PP(16'h66B5,4);
TASK_PP(16'h66B6,4);
TASK_PP(16'h66B7,4);
TASK_PP(16'h66B8,4);
TASK_PP(16'h66B9,4);
TASK_PP(16'h66BA,4);
TASK_PP(16'h66BB,4);
TASK_PP(16'h66BC,4);
TASK_PP(16'h66BD,4);
TASK_PP(16'h66BE,4);
TASK_PP(16'h66BF,4);
TASK_PP(16'h66C0,4);
TASK_PP(16'h66C1,4);
TASK_PP(16'h66C2,4);
TASK_PP(16'h66C3,4);
TASK_PP(16'h66C4,4);
TASK_PP(16'h66C5,4);
TASK_PP(16'h66C6,4);
TASK_PP(16'h66C7,4);
TASK_PP(16'h66C8,4);
TASK_PP(16'h66C9,4);
TASK_PP(16'h66CA,4);
TASK_PP(16'h66CB,4);
TASK_PP(16'h66CC,4);
TASK_PP(16'h66CD,4);
TASK_PP(16'h66CE,4);
TASK_PP(16'h66CF,4);
TASK_PP(16'h66D0,4);
TASK_PP(16'h66D1,4);
TASK_PP(16'h66D2,4);
TASK_PP(16'h66D3,4);
TASK_PP(16'h66D4,4);
TASK_PP(16'h66D5,4);
TASK_PP(16'h66D6,4);
TASK_PP(16'h66D7,4);
TASK_PP(16'h66D8,4);
TASK_PP(16'h66D9,4);
TASK_PP(16'h66DA,4);
TASK_PP(16'h66DB,4);
TASK_PP(16'h66DC,4);
TASK_PP(16'h66DD,4);
TASK_PP(16'h66DE,4);
TASK_PP(16'h66DF,4);
TASK_PP(16'h66E0,4);
TASK_PP(16'h66E1,4);
TASK_PP(16'h66E2,4);
TASK_PP(16'h66E3,4);
TASK_PP(16'h66E4,4);
TASK_PP(16'h66E5,4);
TASK_PP(16'h66E6,4);
TASK_PP(16'h66E7,4);
TASK_PP(16'h66E8,4);
TASK_PP(16'h66E9,4);
TASK_PP(16'h66EA,4);
TASK_PP(16'h66EB,4);
TASK_PP(16'h66EC,4);
TASK_PP(16'h66ED,4);
TASK_PP(16'h66EE,4);
TASK_PP(16'h66EF,4);
TASK_PP(16'h66F0,4);
TASK_PP(16'h66F1,4);
TASK_PP(16'h66F2,4);
TASK_PP(16'h66F3,4);
TASK_PP(16'h66F4,4);
TASK_PP(16'h66F5,4);
TASK_PP(16'h66F6,4);
TASK_PP(16'h66F7,4);
TASK_PP(16'h66F8,4);
TASK_PP(16'h66F9,4);
TASK_PP(16'h66FA,4);
TASK_PP(16'h66FB,4);
TASK_PP(16'h66FC,4);
TASK_PP(16'h66FD,4);
TASK_PP(16'h66FE,4);
TASK_PP(16'h66FF,4);
TASK_PP(16'h6700,4);
TASK_PP(16'h6701,4);
TASK_PP(16'h6702,4);
TASK_PP(16'h6703,4);
TASK_PP(16'h6704,4);
TASK_PP(16'h6705,4);
TASK_PP(16'h6706,4);
TASK_PP(16'h6707,4);
TASK_PP(16'h6708,4);
TASK_PP(16'h6709,4);
TASK_PP(16'h670A,4);
TASK_PP(16'h670B,4);
TASK_PP(16'h670C,4);
TASK_PP(16'h670D,4);
TASK_PP(16'h670E,4);
TASK_PP(16'h670F,4);
TASK_PP(16'h6710,4);
TASK_PP(16'h6711,4);
TASK_PP(16'h6712,4);
TASK_PP(16'h6713,4);
TASK_PP(16'h6714,4);
TASK_PP(16'h6715,4);
TASK_PP(16'h6716,4);
TASK_PP(16'h6717,4);
TASK_PP(16'h6718,4);
TASK_PP(16'h6719,4);
TASK_PP(16'h671A,4);
TASK_PP(16'h671B,4);
TASK_PP(16'h671C,4);
TASK_PP(16'h671D,4);
TASK_PP(16'h671E,4);
TASK_PP(16'h671F,4);
TASK_PP(16'h6720,4);
TASK_PP(16'h6721,4);
TASK_PP(16'h6722,4);
TASK_PP(16'h6723,4);
TASK_PP(16'h6724,4);
TASK_PP(16'h6725,4);
TASK_PP(16'h6726,4);
TASK_PP(16'h6727,4);
TASK_PP(16'h6728,4);
TASK_PP(16'h6729,4);
TASK_PP(16'h672A,4);
TASK_PP(16'h672B,4);
TASK_PP(16'h672C,4);
TASK_PP(16'h672D,4);
TASK_PP(16'h672E,4);
TASK_PP(16'h672F,4);
TASK_PP(16'h6730,4);
TASK_PP(16'h6731,4);
TASK_PP(16'h6732,4);
TASK_PP(16'h6733,4);
TASK_PP(16'h6734,4);
TASK_PP(16'h6735,4);
TASK_PP(16'h6736,4);
TASK_PP(16'h6737,4);
TASK_PP(16'h6738,4);
TASK_PP(16'h6739,4);
TASK_PP(16'h673A,4);
TASK_PP(16'h673B,4);
TASK_PP(16'h673C,4);
TASK_PP(16'h673D,4);
TASK_PP(16'h673E,4);
TASK_PP(16'h673F,4);
TASK_PP(16'h6740,4);
TASK_PP(16'h6741,4);
TASK_PP(16'h6742,4);
TASK_PP(16'h6743,4);
TASK_PP(16'h6744,4);
TASK_PP(16'h6745,4);
TASK_PP(16'h6746,4);
TASK_PP(16'h6747,4);
TASK_PP(16'h6748,4);
TASK_PP(16'h6749,4);
TASK_PP(16'h674A,4);
TASK_PP(16'h674B,4);
TASK_PP(16'h674C,4);
TASK_PP(16'h674D,4);
TASK_PP(16'h674E,4);
TASK_PP(16'h674F,4);
TASK_PP(16'h6750,4);
TASK_PP(16'h6751,4);
TASK_PP(16'h6752,4);
TASK_PP(16'h6753,4);
TASK_PP(16'h6754,4);
TASK_PP(16'h6755,4);
TASK_PP(16'h6756,4);
TASK_PP(16'h6757,4);
TASK_PP(16'h6758,4);
TASK_PP(16'h6759,4);
TASK_PP(16'h675A,4);
TASK_PP(16'h675B,4);
TASK_PP(16'h675C,4);
TASK_PP(16'h675D,4);
TASK_PP(16'h675E,4);
TASK_PP(16'h675F,4);
TASK_PP(16'h6760,4);
TASK_PP(16'h6761,4);
TASK_PP(16'h6762,4);
TASK_PP(16'h6763,4);
TASK_PP(16'h6764,4);
TASK_PP(16'h6765,4);
TASK_PP(16'h6766,4);
TASK_PP(16'h6767,4);
TASK_PP(16'h6768,4);
TASK_PP(16'h6769,4);
TASK_PP(16'h676A,4);
TASK_PP(16'h676B,4);
TASK_PP(16'h676C,4);
TASK_PP(16'h676D,4);
TASK_PP(16'h676E,4);
TASK_PP(16'h676F,4);
TASK_PP(16'h6770,4);
TASK_PP(16'h6771,4);
TASK_PP(16'h6772,4);
TASK_PP(16'h6773,4);
TASK_PP(16'h6774,4);
TASK_PP(16'h6775,4);
TASK_PP(16'h6776,4);
TASK_PP(16'h6777,4);
TASK_PP(16'h6778,4);
TASK_PP(16'h6779,4);
TASK_PP(16'h677A,4);
TASK_PP(16'h677B,4);
TASK_PP(16'h677C,4);
TASK_PP(16'h677D,4);
TASK_PP(16'h677E,4);
TASK_PP(16'h677F,4);
TASK_PP(16'h6780,4);
TASK_PP(16'h6781,4);
TASK_PP(16'h6782,4);
TASK_PP(16'h6783,4);
TASK_PP(16'h6784,4);
TASK_PP(16'h6785,4);
TASK_PP(16'h6786,4);
TASK_PP(16'h6787,4);
TASK_PP(16'h6788,4);
TASK_PP(16'h6789,4);
TASK_PP(16'h678A,4);
TASK_PP(16'h678B,4);
TASK_PP(16'h678C,4);
TASK_PP(16'h678D,4);
TASK_PP(16'h678E,4);
TASK_PP(16'h678F,4);
TASK_PP(16'h6790,4);
TASK_PP(16'h6791,4);
TASK_PP(16'h6792,4);
TASK_PP(16'h6793,4);
TASK_PP(16'h6794,4);
TASK_PP(16'h6795,4);
TASK_PP(16'h6796,4);
TASK_PP(16'h6797,4);
TASK_PP(16'h6798,4);
TASK_PP(16'h6799,4);
TASK_PP(16'h679A,4);
TASK_PP(16'h679B,4);
TASK_PP(16'h679C,4);
TASK_PP(16'h679D,4);
TASK_PP(16'h679E,4);
TASK_PP(16'h679F,4);
TASK_PP(16'h67A0,4);
TASK_PP(16'h67A1,4);
TASK_PP(16'h67A2,4);
TASK_PP(16'h67A3,4);
TASK_PP(16'h67A4,4);
TASK_PP(16'h67A5,4);
TASK_PP(16'h67A6,4);
TASK_PP(16'h67A7,4);
TASK_PP(16'h67A8,4);
TASK_PP(16'h67A9,4);
TASK_PP(16'h67AA,4);
TASK_PP(16'h67AB,4);
TASK_PP(16'h67AC,4);
TASK_PP(16'h67AD,4);
TASK_PP(16'h67AE,4);
TASK_PP(16'h67AF,4);
TASK_PP(16'h67B0,4);
TASK_PP(16'h67B1,4);
TASK_PP(16'h67B2,4);
TASK_PP(16'h67B3,4);
TASK_PP(16'h67B4,4);
TASK_PP(16'h67B5,4);
TASK_PP(16'h67B6,4);
TASK_PP(16'h67B7,4);
TASK_PP(16'h67B8,4);
TASK_PP(16'h67B9,4);
TASK_PP(16'h67BA,4);
TASK_PP(16'h67BB,4);
TASK_PP(16'h67BC,4);
TASK_PP(16'h67BD,4);
TASK_PP(16'h67BE,4);
TASK_PP(16'h67BF,4);
TASK_PP(16'h67C0,4);
TASK_PP(16'h67C1,4);
TASK_PP(16'h67C2,4);
TASK_PP(16'h67C3,4);
TASK_PP(16'h67C4,4);
TASK_PP(16'h67C5,4);
TASK_PP(16'h67C6,4);
TASK_PP(16'h67C7,4);
TASK_PP(16'h67C8,4);
TASK_PP(16'h67C9,4);
TASK_PP(16'h67CA,4);
TASK_PP(16'h67CB,4);
TASK_PP(16'h67CC,4);
TASK_PP(16'h67CD,4);
TASK_PP(16'h67CE,4);
TASK_PP(16'h67CF,4);
TASK_PP(16'h67D0,4);
TASK_PP(16'h67D1,4);
TASK_PP(16'h67D2,4);
TASK_PP(16'h67D3,4);
TASK_PP(16'h67D4,4);
TASK_PP(16'h67D5,4);
TASK_PP(16'h67D6,4);
TASK_PP(16'h67D7,4);
TASK_PP(16'h67D8,4);
TASK_PP(16'h67D9,4);
TASK_PP(16'h67DA,4);
TASK_PP(16'h67DB,4);
TASK_PP(16'h67DC,4);
TASK_PP(16'h67DD,4);
TASK_PP(16'h67DE,4);
TASK_PP(16'h67DF,4);
TASK_PP(16'h67E0,4);
TASK_PP(16'h67E1,4);
TASK_PP(16'h67E2,4);
TASK_PP(16'h67E3,4);
TASK_PP(16'h67E4,4);
TASK_PP(16'h67E5,4);
TASK_PP(16'h67E6,4);
TASK_PP(16'h67E7,4);
TASK_PP(16'h67E8,4);
TASK_PP(16'h67E9,4);
TASK_PP(16'h67EA,4);
TASK_PP(16'h67EB,4);
TASK_PP(16'h67EC,4);
TASK_PP(16'h67ED,4);
TASK_PP(16'h67EE,4);
TASK_PP(16'h67EF,4);
TASK_PP(16'h67F0,4);
TASK_PP(16'h67F1,4);
TASK_PP(16'h67F2,4);
TASK_PP(16'h67F3,4);
TASK_PP(16'h67F4,4);
TASK_PP(16'h67F5,4);
TASK_PP(16'h67F6,4);
TASK_PP(16'h67F7,4);
TASK_PP(16'h67F8,4);
TASK_PP(16'h67F9,4);
TASK_PP(16'h67FA,4);
TASK_PP(16'h67FB,4);
TASK_PP(16'h67FC,4);
TASK_PP(16'h67FD,4);
TASK_PP(16'h67FE,4);
TASK_PP(16'h67FF,4);
TASK_PP(16'h6800,4);
TASK_PP(16'h6801,4);
TASK_PP(16'h6802,4);
TASK_PP(16'h6803,4);
TASK_PP(16'h6804,4);
TASK_PP(16'h6805,4);
TASK_PP(16'h6806,4);
TASK_PP(16'h6807,4);
TASK_PP(16'h6808,4);
TASK_PP(16'h6809,4);
TASK_PP(16'h680A,4);
TASK_PP(16'h680B,4);
TASK_PP(16'h680C,4);
TASK_PP(16'h680D,4);
TASK_PP(16'h680E,4);
TASK_PP(16'h680F,4);
TASK_PP(16'h6810,4);
TASK_PP(16'h6811,4);
TASK_PP(16'h6812,4);
TASK_PP(16'h6813,4);
TASK_PP(16'h6814,4);
TASK_PP(16'h6815,4);
TASK_PP(16'h6816,4);
TASK_PP(16'h6817,4);
TASK_PP(16'h6818,4);
TASK_PP(16'h6819,4);
TASK_PP(16'h681A,4);
TASK_PP(16'h681B,4);
TASK_PP(16'h681C,4);
TASK_PP(16'h681D,4);
TASK_PP(16'h681E,4);
TASK_PP(16'h681F,4);
TASK_PP(16'h6820,4);
TASK_PP(16'h6821,4);
TASK_PP(16'h6822,4);
TASK_PP(16'h6823,4);
TASK_PP(16'h6824,4);
TASK_PP(16'h6825,4);
TASK_PP(16'h6826,4);
TASK_PP(16'h6827,4);
TASK_PP(16'h6828,4);
TASK_PP(16'h6829,4);
TASK_PP(16'h682A,4);
TASK_PP(16'h682B,4);
TASK_PP(16'h682C,4);
TASK_PP(16'h682D,4);
TASK_PP(16'h682E,4);
TASK_PP(16'h682F,4);
TASK_PP(16'h6830,4);
TASK_PP(16'h6831,4);
TASK_PP(16'h6832,4);
TASK_PP(16'h6833,4);
TASK_PP(16'h6834,4);
TASK_PP(16'h6835,4);
TASK_PP(16'h6836,4);
TASK_PP(16'h6837,4);
TASK_PP(16'h6838,4);
TASK_PP(16'h6839,4);
TASK_PP(16'h683A,4);
TASK_PP(16'h683B,4);
TASK_PP(16'h683C,4);
TASK_PP(16'h683D,4);
TASK_PP(16'h683E,4);
TASK_PP(16'h683F,4);
TASK_PP(16'h6840,4);
TASK_PP(16'h6841,4);
TASK_PP(16'h6842,4);
TASK_PP(16'h6843,4);
TASK_PP(16'h6844,4);
TASK_PP(16'h6845,4);
TASK_PP(16'h6846,4);
TASK_PP(16'h6847,4);
TASK_PP(16'h6848,4);
TASK_PP(16'h6849,4);
TASK_PP(16'h684A,4);
TASK_PP(16'h684B,4);
TASK_PP(16'h684C,4);
TASK_PP(16'h684D,4);
TASK_PP(16'h684E,4);
TASK_PP(16'h684F,4);
TASK_PP(16'h6850,4);
TASK_PP(16'h6851,4);
TASK_PP(16'h6852,4);
TASK_PP(16'h6853,4);
TASK_PP(16'h6854,4);
TASK_PP(16'h6855,4);
TASK_PP(16'h6856,4);
TASK_PP(16'h6857,4);
TASK_PP(16'h6858,4);
TASK_PP(16'h6859,4);
TASK_PP(16'h685A,4);
TASK_PP(16'h685B,4);
TASK_PP(16'h685C,4);
TASK_PP(16'h685D,4);
TASK_PP(16'h685E,4);
TASK_PP(16'h685F,4);
TASK_PP(16'h6860,4);
TASK_PP(16'h6861,4);
TASK_PP(16'h6862,4);
TASK_PP(16'h6863,4);
TASK_PP(16'h6864,4);
TASK_PP(16'h6865,4);
TASK_PP(16'h6866,4);
TASK_PP(16'h6867,4);
TASK_PP(16'h6868,4);
TASK_PP(16'h6869,4);
TASK_PP(16'h686A,4);
TASK_PP(16'h686B,4);
TASK_PP(16'h686C,4);
TASK_PP(16'h686D,4);
TASK_PP(16'h686E,4);
TASK_PP(16'h686F,4);
TASK_PP(16'h6870,4);
TASK_PP(16'h6871,4);
TASK_PP(16'h6872,4);
TASK_PP(16'h6873,4);
TASK_PP(16'h6874,4);
TASK_PP(16'h6875,4);
TASK_PP(16'h6876,4);
TASK_PP(16'h6877,4);
TASK_PP(16'h6878,4);
TASK_PP(16'h6879,4);
TASK_PP(16'h687A,4);
TASK_PP(16'h687B,4);
TASK_PP(16'h687C,4);
TASK_PP(16'h687D,4);
TASK_PP(16'h687E,4);
TASK_PP(16'h687F,4);
TASK_PP(16'h6880,4);
TASK_PP(16'h6881,4);
TASK_PP(16'h6882,4);
TASK_PP(16'h6883,4);
TASK_PP(16'h6884,4);
TASK_PP(16'h6885,4);
TASK_PP(16'h6886,4);
TASK_PP(16'h6887,4);
TASK_PP(16'h6888,4);
TASK_PP(16'h6889,4);
TASK_PP(16'h688A,4);
TASK_PP(16'h688B,4);
TASK_PP(16'h688C,4);
TASK_PP(16'h688D,4);
TASK_PP(16'h688E,4);
TASK_PP(16'h688F,4);
TASK_PP(16'h6890,4);
TASK_PP(16'h6891,4);
TASK_PP(16'h6892,4);
TASK_PP(16'h6893,4);
TASK_PP(16'h6894,4);
TASK_PP(16'h6895,4);
TASK_PP(16'h6896,4);
TASK_PP(16'h6897,4);
TASK_PP(16'h6898,4);
TASK_PP(16'h6899,4);
TASK_PP(16'h689A,4);
TASK_PP(16'h689B,4);
TASK_PP(16'h689C,4);
TASK_PP(16'h689D,4);
TASK_PP(16'h689E,4);
TASK_PP(16'h689F,4);
TASK_PP(16'h68A0,4);
TASK_PP(16'h68A1,4);
TASK_PP(16'h68A2,4);
TASK_PP(16'h68A3,4);
TASK_PP(16'h68A4,4);
TASK_PP(16'h68A5,4);
TASK_PP(16'h68A6,4);
TASK_PP(16'h68A7,4);
TASK_PP(16'h68A8,4);
TASK_PP(16'h68A9,4);
TASK_PP(16'h68AA,4);
TASK_PP(16'h68AB,4);
TASK_PP(16'h68AC,4);
TASK_PP(16'h68AD,4);
TASK_PP(16'h68AE,4);
TASK_PP(16'h68AF,4);
TASK_PP(16'h68B0,4);
TASK_PP(16'h68B1,4);
TASK_PP(16'h68B2,4);
TASK_PP(16'h68B3,4);
TASK_PP(16'h68B4,4);
TASK_PP(16'h68B5,4);
TASK_PP(16'h68B6,4);
TASK_PP(16'h68B7,4);
TASK_PP(16'h68B8,4);
TASK_PP(16'h68B9,4);
TASK_PP(16'h68BA,4);
TASK_PP(16'h68BB,4);
TASK_PP(16'h68BC,4);
TASK_PP(16'h68BD,4);
TASK_PP(16'h68BE,4);
TASK_PP(16'h68BF,4);
TASK_PP(16'h68C0,4);
TASK_PP(16'h68C1,4);
TASK_PP(16'h68C2,4);
TASK_PP(16'h68C3,4);
TASK_PP(16'h68C4,4);
TASK_PP(16'h68C5,4);
TASK_PP(16'h68C6,4);
TASK_PP(16'h68C7,4);
TASK_PP(16'h68C8,4);
TASK_PP(16'h68C9,4);
TASK_PP(16'h68CA,4);
TASK_PP(16'h68CB,4);
TASK_PP(16'h68CC,4);
TASK_PP(16'h68CD,4);
TASK_PP(16'h68CE,4);
TASK_PP(16'h68CF,4);
TASK_PP(16'h68D0,4);
TASK_PP(16'h68D1,4);
TASK_PP(16'h68D2,4);
TASK_PP(16'h68D3,4);
TASK_PP(16'h68D4,4);
TASK_PP(16'h68D5,4);
TASK_PP(16'h68D6,4);
TASK_PP(16'h68D7,4);
TASK_PP(16'h68D8,4);
TASK_PP(16'h68D9,4);
TASK_PP(16'h68DA,4);
TASK_PP(16'h68DB,4);
TASK_PP(16'h68DC,4);
TASK_PP(16'h68DD,4);
TASK_PP(16'h68DE,4);
TASK_PP(16'h68DF,4);
TASK_PP(16'h68E0,4);
TASK_PP(16'h68E1,4);
TASK_PP(16'h68E2,4);
TASK_PP(16'h68E3,4);
TASK_PP(16'h68E4,4);
TASK_PP(16'h68E5,4);
TASK_PP(16'h68E6,4);
TASK_PP(16'h68E7,4);
TASK_PP(16'h68E8,4);
TASK_PP(16'h68E9,4);
TASK_PP(16'h68EA,4);
TASK_PP(16'h68EB,4);
TASK_PP(16'h68EC,4);
TASK_PP(16'h68ED,4);
TASK_PP(16'h68EE,4);
TASK_PP(16'h68EF,4);
TASK_PP(16'h68F0,4);
TASK_PP(16'h68F1,4);
TASK_PP(16'h68F2,4);
TASK_PP(16'h68F3,4);
TASK_PP(16'h68F4,4);
TASK_PP(16'h68F5,4);
TASK_PP(16'h68F6,4);
TASK_PP(16'h68F7,4);
TASK_PP(16'h68F8,4);
TASK_PP(16'h68F9,4);
TASK_PP(16'h68FA,4);
TASK_PP(16'h68FB,4);
TASK_PP(16'h68FC,4);
TASK_PP(16'h68FD,4);
TASK_PP(16'h68FE,4);
TASK_PP(16'h68FF,4);
TASK_PP(16'h6900,4);
TASK_PP(16'h6901,4);
TASK_PP(16'h6902,4);
TASK_PP(16'h6903,4);
TASK_PP(16'h6904,4);
TASK_PP(16'h6905,4);
TASK_PP(16'h6906,4);
TASK_PP(16'h6907,4);
TASK_PP(16'h6908,4);
TASK_PP(16'h6909,4);
TASK_PP(16'h690A,4);
TASK_PP(16'h690B,4);
TASK_PP(16'h690C,4);
TASK_PP(16'h690D,4);
TASK_PP(16'h690E,4);
TASK_PP(16'h690F,4);
TASK_PP(16'h6910,4);
TASK_PP(16'h6911,4);
TASK_PP(16'h6912,4);
TASK_PP(16'h6913,4);
TASK_PP(16'h6914,4);
TASK_PP(16'h6915,4);
TASK_PP(16'h6916,4);
TASK_PP(16'h6917,4);
TASK_PP(16'h6918,4);
TASK_PP(16'h6919,4);
TASK_PP(16'h691A,4);
TASK_PP(16'h691B,4);
TASK_PP(16'h691C,4);
TASK_PP(16'h691D,4);
TASK_PP(16'h691E,4);
TASK_PP(16'h691F,4);
TASK_PP(16'h6920,4);
TASK_PP(16'h6921,4);
TASK_PP(16'h6922,4);
TASK_PP(16'h6923,4);
TASK_PP(16'h6924,4);
TASK_PP(16'h6925,4);
TASK_PP(16'h6926,4);
TASK_PP(16'h6927,4);
TASK_PP(16'h6928,4);
TASK_PP(16'h6929,4);
TASK_PP(16'h692A,4);
TASK_PP(16'h692B,4);
TASK_PP(16'h692C,4);
TASK_PP(16'h692D,4);
TASK_PP(16'h692E,4);
TASK_PP(16'h692F,4);
TASK_PP(16'h6930,4);
TASK_PP(16'h6931,4);
TASK_PP(16'h6932,4);
TASK_PP(16'h6933,4);
TASK_PP(16'h6934,4);
TASK_PP(16'h6935,4);
TASK_PP(16'h6936,4);
TASK_PP(16'h6937,4);
TASK_PP(16'h6938,4);
TASK_PP(16'h6939,4);
TASK_PP(16'h693A,4);
TASK_PP(16'h693B,4);
TASK_PP(16'h693C,4);
TASK_PP(16'h693D,4);
TASK_PP(16'h693E,4);
TASK_PP(16'h693F,4);
TASK_PP(16'h6940,4);
TASK_PP(16'h6941,4);
TASK_PP(16'h6942,4);
TASK_PP(16'h6943,4);
TASK_PP(16'h6944,4);
TASK_PP(16'h6945,4);
TASK_PP(16'h6946,4);
TASK_PP(16'h6947,4);
TASK_PP(16'h6948,4);
TASK_PP(16'h6949,4);
TASK_PP(16'h694A,4);
TASK_PP(16'h694B,4);
TASK_PP(16'h694C,4);
TASK_PP(16'h694D,4);
TASK_PP(16'h694E,4);
TASK_PP(16'h694F,4);
TASK_PP(16'h6950,4);
TASK_PP(16'h6951,4);
TASK_PP(16'h6952,4);
TASK_PP(16'h6953,4);
TASK_PP(16'h6954,4);
TASK_PP(16'h6955,4);
TASK_PP(16'h6956,4);
TASK_PP(16'h6957,4);
TASK_PP(16'h6958,4);
TASK_PP(16'h6959,4);
TASK_PP(16'h695A,4);
TASK_PP(16'h695B,4);
TASK_PP(16'h695C,4);
TASK_PP(16'h695D,4);
TASK_PP(16'h695E,4);
TASK_PP(16'h695F,4);
TASK_PP(16'h6960,4);
TASK_PP(16'h6961,4);
TASK_PP(16'h6962,4);
TASK_PP(16'h6963,4);
TASK_PP(16'h6964,4);
TASK_PP(16'h6965,4);
TASK_PP(16'h6966,4);
TASK_PP(16'h6967,4);
TASK_PP(16'h6968,4);
TASK_PP(16'h6969,4);
TASK_PP(16'h696A,4);
TASK_PP(16'h696B,4);
TASK_PP(16'h696C,4);
TASK_PP(16'h696D,4);
TASK_PP(16'h696E,4);
TASK_PP(16'h696F,4);
TASK_PP(16'h6970,4);
TASK_PP(16'h6971,4);
TASK_PP(16'h6972,4);
TASK_PP(16'h6973,4);
TASK_PP(16'h6974,4);
TASK_PP(16'h6975,4);
TASK_PP(16'h6976,4);
TASK_PP(16'h6977,4);
TASK_PP(16'h6978,4);
TASK_PP(16'h6979,4);
TASK_PP(16'h697A,4);
TASK_PP(16'h697B,4);
TASK_PP(16'h697C,4);
TASK_PP(16'h697D,4);
TASK_PP(16'h697E,4);
TASK_PP(16'h697F,4);
TASK_PP(16'h6980,4);
TASK_PP(16'h6981,4);
TASK_PP(16'h6982,4);
TASK_PP(16'h6983,4);
TASK_PP(16'h6984,4);
TASK_PP(16'h6985,4);
TASK_PP(16'h6986,4);
TASK_PP(16'h6987,4);
TASK_PP(16'h6988,4);
TASK_PP(16'h6989,4);
TASK_PP(16'h698A,4);
TASK_PP(16'h698B,4);
TASK_PP(16'h698C,4);
TASK_PP(16'h698D,4);
TASK_PP(16'h698E,4);
TASK_PP(16'h698F,4);
TASK_PP(16'h6990,4);
TASK_PP(16'h6991,4);
TASK_PP(16'h6992,4);
TASK_PP(16'h6993,4);
TASK_PP(16'h6994,4);
TASK_PP(16'h6995,4);
TASK_PP(16'h6996,4);
TASK_PP(16'h6997,4);
TASK_PP(16'h6998,4);
TASK_PP(16'h6999,4);
TASK_PP(16'h699A,4);
TASK_PP(16'h699B,4);
TASK_PP(16'h699C,4);
TASK_PP(16'h699D,4);
TASK_PP(16'h699E,4);
TASK_PP(16'h699F,4);
TASK_PP(16'h69A0,4);
TASK_PP(16'h69A1,4);
TASK_PP(16'h69A2,4);
TASK_PP(16'h69A3,4);
TASK_PP(16'h69A4,4);
TASK_PP(16'h69A5,4);
TASK_PP(16'h69A6,4);
TASK_PP(16'h69A7,4);
TASK_PP(16'h69A8,4);
TASK_PP(16'h69A9,4);
TASK_PP(16'h69AA,4);
TASK_PP(16'h69AB,4);
TASK_PP(16'h69AC,4);
TASK_PP(16'h69AD,4);
TASK_PP(16'h69AE,4);
TASK_PP(16'h69AF,4);
TASK_PP(16'h69B0,4);
TASK_PP(16'h69B1,4);
TASK_PP(16'h69B2,4);
TASK_PP(16'h69B3,4);
TASK_PP(16'h69B4,4);
TASK_PP(16'h69B5,4);
TASK_PP(16'h69B6,4);
TASK_PP(16'h69B7,4);
TASK_PP(16'h69B8,4);
TASK_PP(16'h69B9,4);
TASK_PP(16'h69BA,4);
TASK_PP(16'h69BB,4);
TASK_PP(16'h69BC,4);
TASK_PP(16'h69BD,4);
TASK_PP(16'h69BE,4);
TASK_PP(16'h69BF,4);
TASK_PP(16'h69C0,4);
TASK_PP(16'h69C1,4);
TASK_PP(16'h69C2,4);
TASK_PP(16'h69C3,4);
TASK_PP(16'h69C4,4);
TASK_PP(16'h69C5,4);
TASK_PP(16'h69C6,4);
TASK_PP(16'h69C7,4);
TASK_PP(16'h69C8,4);
TASK_PP(16'h69C9,4);
TASK_PP(16'h69CA,4);
TASK_PP(16'h69CB,4);
TASK_PP(16'h69CC,4);
TASK_PP(16'h69CD,4);
TASK_PP(16'h69CE,4);
TASK_PP(16'h69CF,4);
TASK_PP(16'h69D0,4);
TASK_PP(16'h69D1,4);
TASK_PP(16'h69D2,4);
TASK_PP(16'h69D3,4);
TASK_PP(16'h69D4,4);
TASK_PP(16'h69D5,4);
TASK_PP(16'h69D6,4);
TASK_PP(16'h69D7,4);
TASK_PP(16'h69D8,4);
TASK_PP(16'h69D9,4);
TASK_PP(16'h69DA,4);
TASK_PP(16'h69DB,4);
TASK_PP(16'h69DC,4);
TASK_PP(16'h69DD,4);
TASK_PP(16'h69DE,4);
TASK_PP(16'h69DF,4);
TASK_PP(16'h69E0,4);
TASK_PP(16'h69E1,4);
TASK_PP(16'h69E2,4);
TASK_PP(16'h69E3,4);
TASK_PP(16'h69E4,4);
TASK_PP(16'h69E5,4);
TASK_PP(16'h69E6,4);
TASK_PP(16'h69E7,4);
TASK_PP(16'h69E8,4);
TASK_PP(16'h69E9,4);
TASK_PP(16'h69EA,4);
TASK_PP(16'h69EB,4);
TASK_PP(16'h69EC,4);
TASK_PP(16'h69ED,4);
TASK_PP(16'h69EE,4);
TASK_PP(16'h69EF,4);
TASK_PP(16'h69F0,4);
TASK_PP(16'h69F1,4);
TASK_PP(16'h69F2,4);
TASK_PP(16'h69F3,4);
TASK_PP(16'h69F4,4);
TASK_PP(16'h69F5,4);
TASK_PP(16'h69F6,4);
TASK_PP(16'h69F7,4);
TASK_PP(16'h69F8,4);
TASK_PP(16'h69F9,4);
TASK_PP(16'h69FA,4);
TASK_PP(16'h69FB,4);
TASK_PP(16'h69FC,4);
TASK_PP(16'h69FD,4);
TASK_PP(16'h69FE,4);
TASK_PP(16'h69FF,4);
TASK_PP(16'h6A00,4);
TASK_PP(16'h6A01,4);
TASK_PP(16'h6A02,4);
TASK_PP(16'h6A03,4);
TASK_PP(16'h6A04,4);
TASK_PP(16'h6A05,4);
TASK_PP(16'h6A06,4);
TASK_PP(16'h6A07,4);
TASK_PP(16'h6A08,4);
TASK_PP(16'h6A09,4);
TASK_PP(16'h6A0A,4);
TASK_PP(16'h6A0B,4);
TASK_PP(16'h6A0C,4);
TASK_PP(16'h6A0D,4);
TASK_PP(16'h6A0E,4);
TASK_PP(16'h6A0F,4);
TASK_PP(16'h6A10,4);
TASK_PP(16'h6A11,4);
TASK_PP(16'h6A12,4);
TASK_PP(16'h6A13,4);
TASK_PP(16'h6A14,4);
TASK_PP(16'h6A15,4);
TASK_PP(16'h6A16,4);
TASK_PP(16'h6A17,4);
TASK_PP(16'h6A18,4);
TASK_PP(16'h6A19,4);
TASK_PP(16'h6A1A,4);
TASK_PP(16'h6A1B,4);
TASK_PP(16'h6A1C,4);
TASK_PP(16'h6A1D,4);
TASK_PP(16'h6A1E,4);
TASK_PP(16'h6A1F,4);
TASK_PP(16'h6A20,4);
TASK_PP(16'h6A21,4);
TASK_PP(16'h6A22,4);
TASK_PP(16'h6A23,4);
TASK_PP(16'h6A24,4);
TASK_PP(16'h6A25,4);
TASK_PP(16'h6A26,4);
TASK_PP(16'h6A27,4);
TASK_PP(16'h6A28,4);
TASK_PP(16'h6A29,4);
TASK_PP(16'h6A2A,4);
TASK_PP(16'h6A2B,4);
TASK_PP(16'h6A2C,4);
TASK_PP(16'h6A2D,4);
TASK_PP(16'h6A2E,4);
TASK_PP(16'h6A2F,4);
TASK_PP(16'h6A30,4);
TASK_PP(16'h6A31,4);
TASK_PP(16'h6A32,4);
TASK_PP(16'h6A33,4);
TASK_PP(16'h6A34,4);
TASK_PP(16'h6A35,4);
TASK_PP(16'h6A36,4);
TASK_PP(16'h6A37,4);
TASK_PP(16'h6A38,4);
TASK_PP(16'h6A39,4);
TASK_PP(16'h6A3A,4);
TASK_PP(16'h6A3B,4);
TASK_PP(16'h6A3C,4);
TASK_PP(16'h6A3D,4);
TASK_PP(16'h6A3E,4);
TASK_PP(16'h6A3F,4);
TASK_PP(16'h6A40,4);
TASK_PP(16'h6A41,4);
TASK_PP(16'h6A42,4);
TASK_PP(16'h6A43,4);
TASK_PP(16'h6A44,4);
TASK_PP(16'h6A45,4);
TASK_PP(16'h6A46,4);
TASK_PP(16'h6A47,4);
TASK_PP(16'h6A48,4);
TASK_PP(16'h6A49,4);
TASK_PP(16'h6A4A,4);
TASK_PP(16'h6A4B,4);
TASK_PP(16'h6A4C,4);
TASK_PP(16'h6A4D,4);
TASK_PP(16'h6A4E,4);
TASK_PP(16'h6A4F,4);
TASK_PP(16'h6A50,4);
TASK_PP(16'h6A51,4);
TASK_PP(16'h6A52,4);
TASK_PP(16'h6A53,4);
TASK_PP(16'h6A54,4);
TASK_PP(16'h6A55,4);
TASK_PP(16'h6A56,4);
TASK_PP(16'h6A57,4);
TASK_PP(16'h6A58,4);
TASK_PP(16'h6A59,4);
TASK_PP(16'h6A5A,4);
TASK_PP(16'h6A5B,4);
TASK_PP(16'h6A5C,4);
TASK_PP(16'h6A5D,4);
TASK_PP(16'h6A5E,4);
TASK_PP(16'h6A5F,4);
TASK_PP(16'h6A60,4);
TASK_PP(16'h6A61,4);
TASK_PP(16'h6A62,4);
TASK_PP(16'h6A63,4);
TASK_PP(16'h6A64,4);
TASK_PP(16'h6A65,4);
TASK_PP(16'h6A66,4);
TASK_PP(16'h6A67,4);
TASK_PP(16'h6A68,4);
TASK_PP(16'h6A69,4);
TASK_PP(16'h6A6A,4);
TASK_PP(16'h6A6B,4);
TASK_PP(16'h6A6C,4);
TASK_PP(16'h6A6D,4);
TASK_PP(16'h6A6E,4);
TASK_PP(16'h6A6F,4);
TASK_PP(16'h6A70,4);
TASK_PP(16'h6A71,4);
TASK_PP(16'h6A72,4);
TASK_PP(16'h6A73,4);
TASK_PP(16'h6A74,4);
TASK_PP(16'h6A75,4);
TASK_PP(16'h6A76,4);
TASK_PP(16'h6A77,4);
TASK_PP(16'h6A78,4);
TASK_PP(16'h6A79,4);
TASK_PP(16'h6A7A,4);
TASK_PP(16'h6A7B,4);
TASK_PP(16'h6A7C,4);
TASK_PP(16'h6A7D,4);
TASK_PP(16'h6A7E,4);
TASK_PP(16'h6A7F,4);
TASK_PP(16'h6A80,4);
TASK_PP(16'h6A81,4);
TASK_PP(16'h6A82,4);
TASK_PP(16'h6A83,4);
TASK_PP(16'h6A84,4);
TASK_PP(16'h6A85,4);
TASK_PP(16'h6A86,4);
TASK_PP(16'h6A87,4);
TASK_PP(16'h6A88,4);
TASK_PP(16'h6A89,4);
TASK_PP(16'h6A8A,4);
TASK_PP(16'h6A8B,4);
TASK_PP(16'h6A8C,4);
TASK_PP(16'h6A8D,4);
TASK_PP(16'h6A8E,4);
TASK_PP(16'h6A8F,4);
TASK_PP(16'h6A90,4);
TASK_PP(16'h6A91,4);
TASK_PP(16'h6A92,4);
TASK_PP(16'h6A93,4);
TASK_PP(16'h6A94,4);
TASK_PP(16'h6A95,4);
TASK_PP(16'h6A96,4);
TASK_PP(16'h6A97,4);
TASK_PP(16'h6A98,4);
TASK_PP(16'h6A99,4);
TASK_PP(16'h6A9A,4);
TASK_PP(16'h6A9B,4);
TASK_PP(16'h6A9C,4);
TASK_PP(16'h6A9D,4);
TASK_PP(16'h6A9E,4);
TASK_PP(16'h6A9F,4);
TASK_PP(16'h6AA0,4);
TASK_PP(16'h6AA1,4);
TASK_PP(16'h6AA2,4);
TASK_PP(16'h6AA3,4);
TASK_PP(16'h6AA4,4);
TASK_PP(16'h6AA5,4);
TASK_PP(16'h6AA6,4);
TASK_PP(16'h6AA7,4);
TASK_PP(16'h6AA8,4);
TASK_PP(16'h6AA9,4);
TASK_PP(16'h6AAA,4);
TASK_PP(16'h6AAB,4);
TASK_PP(16'h6AAC,4);
TASK_PP(16'h6AAD,4);
TASK_PP(16'h6AAE,4);
TASK_PP(16'h6AAF,4);
TASK_PP(16'h6AB0,4);
TASK_PP(16'h6AB1,4);
TASK_PP(16'h6AB2,4);
TASK_PP(16'h6AB3,4);
TASK_PP(16'h6AB4,4);
TASK_PP(16'h6AB5,4);
TASK_PP(16'h6AB6,4);
TASK_PP(16'h6AB7,4);
TASK_PP(16'h6AB8,4);
TASK_PP(16'h6AB9,4);
TASK_PP(16'h6ABA,4);
TASK_PP(16'h6ABB,4);
TASK_PP(16'h6ABC,4);
TASK_PP(16'h6ABD,4);
TASK_PP(16'h6ABE,4);
TASK_PP(16'h6ABF,4);
TASK_PP(16'h6AC0,4);
TASK_PP(16'h6AC1,4);
TASK_PP(16'h6AC2,4);
TASK_PP(16'h6AC3,4);
TASK_PP(16'h6AC4,4);
TASK_PP(16'h6AC5,4);
TASK_PP(16'h6AC6,4);
TASK_PP(16'h6AC7,4);
TASK_PP(16'h6AC8,4);
TASK_PP(16'h6AC9,4);
TASK_PP(16'h6ACA,4);
TASK_PP(16'h6ACB,4);
TASK_PP(16'h6ACC,4);
TASK_PP(16'h6ACD,4);
TASK_PP(16'h6ACE,4);
TASK_PP(16'h6ACF,4);
TASK_PP(16'h6AD0,4);
TASK_PP(16'h6AD1,4);
TASK_PP(16'h6AD2,4);
TASK_PP(16'h6AD3,4);
TASK_PP(16'h6AD4,4);
TASK_PP(16'h6AD5,4);
TASK_PP(16'h6AD6,4);
TASK_PP(16'h6AD7,4);
TASK_PP(16'h6AD8,4);
TASK_PP(16'h6AD9,4);
TASK_PP(16'h6ADA,4);
TASK_PP(16'h6ADB,4);
TASK_PP(16'h6ADC,4);
TASK_PP(16'h6ADD,4);
TASK_PP(16'h6ADE,4);
TASK_PP(16'h6ADF,4);
TASK_PP(16'h6AE0,4);
TASK_PP(16'h6AE1,4);
TASK_PP(16'h6AE2,4);
TASK_PP(16'h6AE3,4);
TASK_PP(16'h6AE4,4);
TASK_PP(16'h6AE5,4);
TASK_PP(16'h6AE6,4);
TASK_PP(16'h6AE7,4);
TASK_PP(16'h6AE8,4);
TASK_PP(16'h6AE9,4);
TASK_PP(16'h6AEA,4);
TASK_PP(16'h6AEB,4);
TASK_PP(16'h6AEC,4);
TASK_PP(16'h6AED,4);
TASK_PP(16'h6AEE,4);
TASK_PP(16'h6AEF,4);
TASK_PP(16'h6AF0,4);
TASK_PP(16'h6AF1,4);
TASK_PP(16'h6AF2,4);
TASK_PP(16'h6AF3,4);
TASK_PP(16'h6AF4,4);
TASK_PP(16'h6AF5,4);
TASK_PP(16'h6AF6,4);
TASK_PP(16'h6AF7,4);
TASK_PP(16'h6AF8,4);
TASK_PP(16'h6AF9,4);
TASK_PP(16'h6AFA,4);
TASK_PP(16'h6AFB,4);
TASK_PP(16'h6AFC,4);
TASK_PP(16'h6AFD,4);
TASK_PP(16'h6AFE,4);
TASK_PP(16'h6AFF,4);
TASK_PP(16'h6B00,4);
TASK_PP(16'h6B01,4);
TASK_PP(16'h6B02,4);
TASK_PP(16'h6B03,4);
TASK_PP(16'h6B04,4);
TASK_PP(16'h6B05,4);
TASK_PP(16'h6B06,4);
TASK_PP(16'h6B07,4);
TASK_PP(16'h6B08,4);
TASK_PP(16'h6B09,4);
TASK_PP(16'h6B0A,4);
TASK_PP(16'h6B0B,4);
TASK_PP(16'h6B0C,4);
TASK_PP(16'h6B0D,4);
TASK_PP(16'h6B0E,4);
TASK_PP(16'h6B0F,4);
TASK_PP(16'h6B10,4);
TASK_PP(16'h6B11,4);
TASK_PP(16'h6B12,4);
TASK_PP(16'h6B13,4);
TASK_PP(16'h6B14,4);
TASK_PP(16'h6B15,4);
TASK_PP(16'h6B16,4);
TASK_PP(16'h6B17,4);
TASK_PP(16'h6B18,4);
TASK_PP(16'h6B19,4);
TASK_PP(16'h6B1A,4);
TASK_PP(16'h6B1B,4);
TASK_PP(16'h6B1C,4);
TASK_PP(16'h6B1D,4);
TASK_PP(16'h6B1E,4);
TASK_PP(16'h6B1F,4);
TASK_PP(16'h6B20,4);
TASK_PP(16'h6B21,4);
TASK_PP(16'h6B22,4);
TASK_PP(16'h6B23,4);
TASK_PP(16'h6B24,4);
TASK_PP(16'h6B25,4);
TASK_PP(16'h6B26,4);
TASK_PP(16'h6B27,4);
TASK_PP(16'h6B28,4);
TASK_PP(16'h6B29,4);
TASK_PP(16'h6B2A,4);
TASK_PP(16'h6B2B,4);
TASK_PP(16'h6B2C,4);
TASK_PP(16'h6B2D,4);
TASK_PP(16'h6B2E,4);
TASK_PP(16'h6B2F,4);
TASK_PP(16'h6B30,4);
TASK_PP(16'h6B31,4);
TASK_PP(16'h6B32,4);
TASK_PP(16'h6B33,4);
TASK_PP(16'h6B34,4);
TASK_PP(16'h6B35,4);
TASK_PP(16'h6B36,4);
TASK_PP(16'h6B37,4);
TASK_PP(16'h6B38,4);
TASK_PP(16'h6B39,4);
TASK_PP(16'h6B3A,4);
TASK_PP(16'h6B3B,4);
TASK_PP(16'h6B3C,4);
TASK_PP(16'h6B3D,4);
TASK_PP(16'h6B3E,4);
TASK_PP(16'h6B3F,4);
TASK_PP(16'h6B40,4);
TASK_PP(16'h6B41,4);
TASK_PP(16'h6B42,4);
TASK_PP(16'h6B43,4);
TASK_PP(16'h6B44,4);
TASK_PP(16'h6B45,4);
TASK_PP(16'h6B46,4);
TASK_PP(16'h6B47,4);
TASK_PP(16'h6B48,4);
TASK_PP(16'h6B49,4);
TASK_PP(16'h6B4A,4);
TASK_PP(16'h6B4B,4);
TASK_PP(16'h6B4C,4);
TASK_PP(16'h6B4D,4);
TASK_PP(16'h6B4E,4);
TASK_PP(16'h6B4F,4);
TASK_PP(16'h6B50,4);
TASK_PP(16'h6B51,4);
TASK_PP(16'h6B52,4);
TASK_PP(16'h6B53,4);
TASK_PP(16'h6B54,4);
TASK_PP(16'h6B55,4);
TASK_PP(16'h6B56,4);
TASK_PP(16'h6B57,4);
TASK_PP(16'h6B58,4);
TASK_PP(16'h6B59,4);
TASK_PP(16'h6B5A,4);
TASK_PP(16'h6B5B,4);
TASK_PP(16'h6B5C,4);
TASK_PP(16'h6B5D,4);
TASK_PP(16'h6B5E,4);
TASK_PP(16'h6B5F,4);
TASK_PP(16'h6B60,4);
TASK_PP(16'h6B61,4);
TASK_PP(16'h6B62,4);
TASK_PP(16'h6B63,4);
TASK_PP(16'h6B64,4);
TASK_PP(16'h6B65,4);
TASK_PP(16'h6B66,4);
TASK_PP(16'h6B67,4);
TASK_PP(16'h6B68,4);
TASK_PP(16'h6B69,4);
TASK_PP(16'h6B6A,4);
TASK_PP(16'h6B6B,4);
TASK_PP(16'h6B6C,4);
TASK_PP(16'h6B6D,4);
TASK_PP(16'h6B6E,4);
TASK_PP(16'h6B6F,4);
TASK_PP(16'h6B70,4);
TASK_PP(16'h6B71,4);
TASK_PP(16'h6B72,4);
TASK_PP(16'h6B73,4);
TASK_PP(16'h6B74,4);
TASK_PP(16'h6B75,4);
TASK_PP(16'h6B76,4);
TASK_PP(16'h6B77,4);
TASK_PP(16'h6B78,4);
TASK_PP(16'h6B79,4);
TASK_PP(16'h6B7A,4);
TASK_PP(16'h6B7B,4);
TASK_PP(16'h6B7C,4);
TASK_PP(16'h6B7D,4);
TASK_PP(16'h6B7E,4);
TASK_PP(16'h6B7F,4);
TASK_PP(16'h6B80,4);
TASK_PP(16'h6B81,4);
TASK_PP(16'h6B82,4);
TASK_PP(16'h6B83,4);
TASK_PP(16'h6B84,4);
TASK_PP(16'h6B85,4);
TASK_PP(16'h6B86,4);
TASK_PP(16'h6B87,4);
TASK_PP(16'h6B88,4);
TASK_PP(16'h6B89,4);
TASK_PP(16'h6B8A,4);
TASK_PP(16'h6B8B,4);
TASK_PP(16'h6B8C,4);
TASK_PP(16'h6B8D,4);
TASK_PP(16'h6B8E,4);
TASK_PP(16'h6B8F,4);
TASK_PP(16'h6B90,4);
TASK_PP(16'h6B91,4);
TASK_PP(16'h6B92,4);
TASK_PP(16'h6B93,4);
TASK_PP(16'h6B94,4);
TASK_PP(16'h6B95,4);
TASK_PP(16'h6B96,4);
TASK_PP(16'h6B97,4);
TASK_PP(16'h6B98,4);
TASK_PP(16'h6B99,4);
TASK_PP(16'h6B9A,4);
TASK_PP(16'h6B9B,4);
TASK_PP(16'h6B9C,4);
TASK_PP(16'h6B9D,4);
TASK_PP(16'h6B9E,4);
TASK_PP(16'h6B9F,4);
TASK_PP(16'h6BA0,4);
TASK_PP(16'h6BA1,4);
TASK_PP(16'h6BA2,4);
TASK_PP(16'h6BA3,4);
TASK_PP(16'h6BA4,4);
TASK_PP(16'h6BA5,4);
TASK_PP(16'h6BA6,4);
TASK_PP(16'h6BA7,4);
TASK_PP(16'h6BA8,4);
TASK_PP(16'h6BA9,4);
TASK_PP(16'h6BAA,4);
TASK_PP(16'h6BAB,4);
TASK_PP(16'h6BAC,4);
TASK_PP(16'h6BAD,4);
TASK_PP(16'h6BAE,4);
TASK_PP(16'h6BAF,4);
TASK_PP(16'h6BB0,4);
TASK_PP(16'h6BB1,4);
TASK_PP(16'h6BB2,4);
TASK_PP(16'h6BB3,4);
TASK_PP(16'h6BB4,4);
TASK_PP(16'h6BB5,4);
TASK_PP(16'h6BB6,4);
TASK_PP(16'h6BB7,4);
TASK_PP(16'h6BB8,4);
TASK_PP(16'h6BB9,4);
TASK_PP(16'h6BBA,4);
TASK_PP(16'h6BBB,4);
TASK_PP(16'h6BBC,4);
TASK_PP(16'h6BBD,4);
TASK_PP(16'h6BBE,4);
TASK_PP(16'h6BBF,4);
TASK_PP(16'h6BC0,4);
TASK_PP(16'h6BC1,4);
TASK_PP(16'h6BC2,4);
TASK_PP(16'h6BC3,4);
TASK_PP(16'h6BC4,4);
TASK_PP(16'h6BC5,4);
TASK_PP(16'h6BC6,4);
TASK_PP(16'h6BC7,4);
TASK_PP(16'h6BC8,4);
TASK_PP(16'h6BC9,4);
TASK_PP(16'h6BCA,4);
TASK_PP(16'h6BCB,4);
TASK_PP(16'h6BCC,4);
TASK_PP(16'h6BCD,4);
TASK_PP(16'h6BCE,4);
TASK_PP(16'h6BCF,4);
TASK_PP(16'h6BD0,4);
TASK_PP(16'h6BD1,4);
TASK_PP(16'h6BD2,4);
TASK_PP(16'h6BD3,4);
TASK_PP(16'h6BD4,4);
TASK_PP(16'h6BD5,4);
TASK_PP(16'h6BD6,4);
TASK_PP(16'h6BD7,4);
TASK_PP(16'h6BD8,4);
TASK_PP(16'h6BD9,4);
TASK_PP(16'h6BDA,4);
TASK_PP(16'h6BDB,4);
TASK_PP(16'h6BDC,4);
TASK_PP(16'h6BDD,4);
TASK_PP(16'h6BDE,4);
TASK_PP(16'h6BDF,4);
TASK_PP(16'h6BE0,4);
TASK_PP(16'h6BE1,4);
TASK_PP(16'h6BE2,4);
TASK_PP(16'h6BE3,4);
TASK_PP(16'h6BE4,4);
TASK_PP(16'h6BE5,4);
TASK_PP(16'h6BE6,4);
TASK_PP(16'h6BE7,4);
TASK_PP(16'h6BE8,4);
TASK_PP(16'h6BE9,4);
TASK_PP(16'h6BEA,4);
TASK_PP(16'h6BEB,4);
TASK_PP(16'h6BEC,4);
TASK_PP(16'h6BED,4);
TASK_PP(16'h6BEE,4);
TASK_PP(16'h6BEF,4);
TASK_PP(16'h6BF0,4);
TASK_PP(16'h6BF1,4);
TASK_PP(16'h6BF2,4);
TASK_PP(16'h6BF3,4);
TASK_PP(16'h6BF4,4);
TASK_PP(16'h6BF5,4);
TASK_PP(16'h6BF6,4);
TASK_PP(16'h6BF7,4);
TASK_PP(16'h6BF8,4);
TASK_PP(16'h6BF9,4);
TASK_PP(16'h6BFA,4);
TASK_PP(16'h6BFB,4);
TASK_PP(16'h6BFC,4);
TASK_PP(16'h6BFD,4);
TASK_PP(16'h6BFE,4);
TASK_PP(16'h6BFF,4);
TASK_PP(16'h6C00,4);
TASK_PP(16'h6C01,4);
TASK_PP(16'h6C02,4);
TASK_PP(16'h6C03,4);
TASK_PP(16'h6C04,4);
TASK_PP(16'h6C05,4);
TASK_PP(16'h6C06,4);
TASK_PP(16'h6C07,4);
TASK_PP(16'h6C08,4);
TASK_PP(16'h6C09,4);
TASK_PP(16'h6C0A,4);
TASK_PP(16'h6C0B,4);
TASK_PP(16'h6C0C,4);
TASK_PP(16'h6C0D,4);
TASK_PP(16'h6C0E,4);
TASK_PP(16'h6C0F,4);
TASK_PP(16'h6C10,4);
TASK_PP(16'h6C11,4);
TASK_PP(16'h6C12,4);
TASK_PP(16'h6C13,4);
TASK_PP(16'h6C14,4);
TASK_PP(16'h6C15,4);
TASK_PP(16'h6C16,4);
TASK_PP(16'h6C17,4);
TASK_PP(16'h6C18,4);
TASK_PP(16'h6C19,4);
TASK_PP(16'h6C1A,4);
TASK_PP(16'h6C1B,4);
TASK_PP(16'h6C1C,4);
TASK_PP(16'h6C1D,4);
TASK_PP(16'h6C1E,4);
TASK_PP(16'h6C1F,4);
TASK_PP(16'h6C20,4);
TASK_PP(16'h6C21,4);
TASK_PP(16'h6C22,4);
TASK_PP(16'h6C23,4);
TASK_PP(16'h6C24,4);
TASK_PP(16'h6C25,4);
TASK_PP(16'h6C26,4);
TASK_PP(16'h6C27,4);
TASK_PP(16'h6C28,4);
TASK_PP(16'h6C29,4);
TASK_PP(16'h6C2A,4);
TASK_PP(16'h6C2B,4);
TASK_PP(16'h6C2C,4);
TASK_PP(16'h6C2D,4);
TASK_PP(16'h6C2E,4);
TASK_PP(16'h6C2F,4);
TASK_PP(16'h6C30,4);
TASK_PP(16'h6C31,4);
TASK_PP(16'h6C32,4);
TASK_PP(16'h6C33,4);
TASK_PP(16'h6C34,4);
TASK_PP(16'h6C35,4);
TASK_PP(16'h6C36,4);
TASK_PP(16'h6C37,4);
TASK_PP(16'h6C38,4);
TASK_PP(16'h6C39,4);
TASK_PP(16'h6C3A,4);
TASK_PP(16'h6C3B,4);
TASK_PP(16'h6C3C,4);
TASK_PP(16'h6C3D,4);
TASK_PP(16'h6C3E,4);
TASK_PP(16'h6C3F,4);
TASK_PP(16'h6C40,4);
TASK_PP(16'h6C41,4);
TASK_PP(16'h6C42,4);
TASK_PP(16'h6C43,4);
TASK_PP(16'h6C44,4);
TASK_PP(16'h6C45,4);
TASK_PP(16'h6C46,4);
TASK_PP(16'h6C47,4);
TASK_PP(16'h6C48,4);
TASK_PP(16'h6C49,4);
TASK_PP(16'h6C4A,4);
TASK_PP(16'h6C4B,4);
TASK_PP(16'h6C4C,4);
TASK_PP(16'h6C4D,4);
TASK_PP(16'h6C4E,4);
TASK_PP(16'h6C4F,4);
TASK_PP(16'h6C50,4);
TASK_PP(16'h6C51,4);
TASK_PP(16'h6C52,4);
TASK_PP(16'h6C53,4);
TASK_PP(16'h6C54,4);
TASK_PP(16'h6C55,4);
TASK_PP(16'h6C56,4);
TASK_PP(16'h6C57,4);
TASK_PP(16'h6C58,4);
TASK_PP(16'h6C59,4);
TASK_PP(16'h6C5A,4);
TASK_PP(16'h6C5B,4);
TASK_PP(16'h6C5C,4);
TASK_PP(16'h6C5D,4);
TASK_PP(16'h6C5E,4);
TASK_PP(16'h6C5F,4);
TASK_PP(16'h6C60,4);
TASK_PP(16'h6C61,4);
TASK_PP(16'h6C62,4);
TASK_PP(16'h6C63,4);
TASK_PP(16'h6C64,4);
TASK_PP(16'h6C65,4);
TASK_PP(16'h6C66,4);
TASK_PP(16'h6C67,4);
TASK_PP(16'h6C68,4);
TASK_PP(16'h6C69,4);
TASK_PP(16'h6C6A,4);
TASK_PP(16'h6C6B,4);
TASK_PP(16'h6C6C,4);
TASK_PP(16'h6C6D,4);
TASK_PP(16'h6C6E,4);
TASK_PP(16'h6C6F,4);
TASK_PP(16'h6C70,4);
TASK_PP(16'h6C71,4);
TASK_PP(16'h6C72,4);
TASK_PP(16'h6C73,4);
TASK_PP(16'h6C74,4);
TASK_PP(16'h6C75,4);
TASK_PP(16'h6C76,4);
TASK_PP(16'h6C77,4);
TASK_PP(16'h6C78,4);
TASK_PP(16'h6C79,4);
TASK_PP(16'h6C7A,4);
TASK_PP(16'h6C7B,4);
TASK_PP(16'h6C7C,4);
TASK_PP(16'h6C7D,4);
TASK_PP(16'h6C7E,4);
TASK_PP(16'h6C7F,4);
TASK_PP(16'h6C80,4);
TASK_PP(16'h6C81,4);
TASK_PP(16'h6C82,4);
TASK_PP(16'h6C83,4);
TASK_PP(16'h6C84,4);
TASK_PP(16'h6C85,4);
TASK_PP(16'h6C86,4);
TASK_PP(16'h6C87,4);
TASK_PP(16'h6C88,4);
TASK_PP(16'h6C89,4);
TASK_PP(16'h6C8A,4);
TASK_PP(16'h6C8B,4);
TASK_PP(16'h6C8C,4);
TASK_PP(16'h6C8D,4);
TASK_PP(16'h6C8E,4);
TASK_PP(16'h6C8F,4);
TASK_PP(16'h6C90,4);
TASK_PP(16'h6C91,4);
TASK_PP(16'h6C92,4);
TASK_PP(16'h6C93,4);
TASK_PP(16'h6C94,4);
TASK_PP(16'h6C95,4);
TASK_PP(16'h6C96,4);
TASK_PP(16'h6C97,4);
TASK_PP(16'h6C98,4);
TASK_PP(16'h6C99,4);
TASK_PP(16'h6C9A,4);
TASK_PP(16'h6C9B,4);
TASK_PP(16'h6C9C,4);
TASK_PP(16'h6C9D,4);
TASK_PP(16'h6C9E,4);
TASK_PP(16'h6C9F,4);
TASK_PP(16'h6CA0,4);
TASK_PP(16'h6CA1,4);
TASK_PP(16'h6CA2,4);
TASK_PP(16'h6CA3,4);
TASK_PP(16'h6CA4,4);
TASK_PP(16'h6CA5,4);
TASK_PP(16'h6CA6,4);
TASK_PP(16'h6CA7,4);
TASK_PP(16'h6CA8,4);
TASK_PP(16'h6CA9,4);
TASK_PP(16'h6CAA,4);
TASK_PP(16'h6CAB,4);
TASK_PP(16'h6CAC,4);
TASK_PP(16'h6CAD,4);
TASK_PP(16'h6CAE,4);
TASK_PP(16'h6CAF,4);
TASK_PP(16'h6CB0,4);
TASK_PP(16'h6CB1,4);
TASK_PP(16'h6CB2,4);
TASK_PP(16'h6CB3,4);
TASK_PP(16'h6CB4,4);
TASK_PP(16'h6CB5,4);
TASK_PP(16'h6CB6,4);
TASK_PP(16'h6CB7,4);
TASK_PP(16'h6CB8,4);
TASK_PP(16'h6CB9,4);
TASK_PP(16'h6CBA,4);
TASK_PP(16'h6CBB,4);
TASK_PP(16'h6CBC,4);
TASK_PP(16'h6CBD,4);
TASK_PP(16'h6CBE,4);
TASK_PP(16'h6CBF,4);
TASK_PP(16'h6CC0,4);
TASK_PP(16'h6CC1,4);
TASK_PP(16'h6CC2,4);
TASK_PP(16'h6CC3,4);
TASK_PP(16'h6CC4,4);
TASK_PP(16'h6CC5,4);
TASK_PP(16'h6CC6,4);
TASK_PP(16'h6CC7,4);
TASK_PP(16'h6CC8,4);
TASK_PP(16'h6CC9,4);
TASK_PP(16'h6CCA,4);
TASK_PP(16'h6CCB,4);
TASK_PP(16'h6CCC,4);
TASK_PP(16'h6CCD,4);
TASK_PP(16'h6CCE,4);
TASK_PP(16'h6CCF,4);
TASK_PP(16'h6CD0,4);
TASK_PP(16'h6CD1,4);
TASK_PP(16'h6CD2,4);
TASK_PP(16'h6CD3,4);
TASK_PP(16'h6CD4,4);
TASK_PP(16'h6CD5,4);
TASK_PP(16'h6CD6,4);
TASK_PP(16'h6CD7,4);
TASK_PP(16'h6CD8,4);
TASK_PP(16'h6CD9,4);
TASK_PP(16'h6CDA,4);
TASK_PP(16'h6CDB,4);
TASK_PP(16'h6CDC,4);
TASK_PP(16'h6CDD,4);
TASK_PP(16'h6CDE,4);
TASK_PP(16'h6CDF,4);
TASK_PP(16'h6CE0,4);
TASK_PP(16'h6CE1,4);
TASK_PP(16'h6CE2,4);
TASK_PP(16'h6CE3,4);
TASK_PP(16'h6CE4,4);
TASK_PP(16'h6CE5,4);
TASK_PP(16'h6CE6,4);
TASK_PP(16'h6CE7,4);
TASK_PP(16'h6CE8,4);
TASK_PP(16'h6CE9,4);
TASK_PP(16'h6CEA,4);
TASK_PP(16'h6CEB,4);
TASK_PP(16'h6CEC,4);
TASK_PP(16'h6CED,4);
TASK_PP(16'h6CEE,4);
TASK_PP(16'h6CEF,4);
TASK_PP(16'h6CF0,4);
TASK_PP(16'h6CF1,4);
TASK_PP(16'h6CF2,4);
TASK_PP(16'h6CF3,4);
TASK_PP(16'h6CF4,4);
TASK_PP(16'h6CF5,4);
TASK_PP(16'h6CF6,4);
TASK_PP(16'h6CF7,4);
TASK_PP(16'h6CF8,4);
TASK_PP(16'h6CF9,4);
TASK_PP(16'h6CFA,4);
TASK_PP(16'h6CFB,4);
TASK_PP(16'h6CFC,4);
TASK_PP(16'h6CFD,4);
TASK_PP(16'h6CFE,4);
TASK_PP(16'h6CFF,4);
TASK_PP(16'h6D00,4);
TASK_PP(16'h6D01,4);
TASK_PP(16'h6D02,4);
TASK_PP(16'h6D03,4);
TASK_PP(16'h6D04,4);
TASK_PP(16'h6D05,4);
TASK_PP(16'h6D06,4);
TASK_PP(16'h6D07,4);
TASK_PP(16'h6D08,4);
TASK_PP(16'h6D09,4);
TASK_PP(16'h6D0A,4);
TASK_PP(16'h6D0B,4);
TASK_PP(16'h6D0C,4);
TASK_PP(16'h6D0D,4);
TASK_PP(16'h6D0E,4);
TASK_PP(16'h6D0F,4);
TASK_PP(16'h6D10,4);
TASK_PP(16'h6D11,4);
TASK_PP(16'h6D12,4);
TASK_PP(16'h6D13,4);
TASK_PP(16'h6D14,4);
TASK_PP(16'h6D15,4);
TASK_PP(16'h6D16,4);
TASK_PP(16'h6D17,4);
TASK_PP(16'h6D18,4);
TASK_PP(16'h6D19,4);
TASK_PP(16'h6D1A,4);
TASK_PP(16'h6D1B,4);
TASK_PP(16'h6D1C,4);
TASK_PP(16'h6D1D,4);
TASK_PP(16'h6D1E,4);
TASK_PP(16'h6D1F,4);
TASK_PP(16'h6D20,4);
TASK_PP(16'h6D21,4);
TASK_PP(16'h6D22,4);
TASK_PP(16'h6D23,4);
TASK_PP(16'h6D24,4);
TASK_PP(16'h6D25,4);
TASK_PP(16'h6D26,4);
TASK_PP(16'h6D27,4);
TASK_PP(16'h6D28,4);
TASK_PP(16'h6D29,4);
TASK_PP(16'h6D2A,4);
TASK_PP(16'h6D2B,4);
TASK_PP(16'h6D2C,4);
TASK_PP(16'h6D2D,4);
TASK_PP(16'h6D2E,4);
TASK_PP(16'h6D2F,4);
TASK_PP(16'h6D30,4);
TASK_PP(16'h6D31,4);
TASK_PP(16'h6D32,4);
TASK_PP(16'h6D33,4);
TASK_PP(16'h6D34,4);
TASK_PP(16'h6D35,4);
TASK_PP(16'h6D36,4);
TASK_PP(16'h6D37,4);
TASK_PP(16'h6D38,4);
TASK_PP(16'h6D39,4);
TASK_PP(16'h6D3A,4);
TASK_PP(16'h6D3B,4);
TASK_PP(16'h6D3C,4);
TASK_PP(16'h6D3D,4);
TASK_PP(16'h6D3E,4);
TASK_PP(16'h6D3F,4);
TASK_PP(16'h6D40,4);
TASK_PP(16'h6D41,4);
TASK_PP(16'h6D42,4);
TASK_PP(16'h6D43,4);
TASK_PP(16'h6D44,4);
TASK_PP(16'h6D45,4);
TASK_PP(16'h6D46,4);
TASK_PP(16'h6D47,4);
TASK_PP(16'h6D48,4);
TASK_PP(16'h6D49,4);
TASK_PP(16'h6D4A,4);
TASK_PP(16'h6D4B,4);
TASK_PP(16'h6D4C,4);
TASK_PP(16'h6D4D,4);
TASK_PP(16'h6D4E,4);
TASK_PP(16'h6D4F,4);
TASK_PP(16'h6D50,4);
TASK_PP(16'h6D51,4);
TASK_PP(16'h6D52,4);
TASK_PP(16'h6D53,4);
TASK_PP(16'h6D54,4);
TASK_PP(16'h6D55,4);
TASK_PP(16'h6D56,4);
TASK_PP(16'h6D57,4);
TASK_PP(16'h6D58,4);
TASK_PP(16'h6D59,4);
TASK_PP(16'h6D5A,4);
TASK_PP(16'h6D5B,4);
TASK_PP(16'h6D5C,4);
TASK_PP(16'h6D5D,4);
TASK_PP(16'h6D5E,4);
TASK_PP(16'h6D5F,4);
TASK_PP(16'h6D60,4);
TASK_PP(16'h6D61,4);
TASK_PP(16'h6D62,4);
TASK_PP(16'h6D63,4);
TASK_PP(16'h6D64,4);
TASK_PP(16'h6D65,4);
TASK_PP(16'h6D66,4);
TASK_PP(16'h6D67,4);
TASK_PP(16'h6D68,4);
TASK_PP(16'h6D69,4);
TASK_PP(16'h6D6A,4);
TASK_PP(16'h6D6B,4);
TASK_PP(16'h6D6C,4);
TASK_PP(16'h6D6D,4);
TASK_PP(16'h6D6E,4);
TASK_PP(16'h6D6F,4);
TASK_PP(16'h6D70,4);
TASK_PP(16'h6D71,4);
TASK_PP(16'h6D72,4);
TASK_PP(16'h6D73,4);
TASK_PP(16'h6D74,4);
TASK_PP(16'h6D75,4);
TASK_PP(16'h6D76,4);
TASK_PP(16'h6D77,4);
TASK_PP(16'h6D78,4);
TASK_PP(16'h6D79,4);
TASK_PP(16'h6D7A,4);
TASK_PP(16'h6D7B,4);
TASK_PP(16'h6D7C,4);
TASK_PP(16'h6D7D,4);
TASK_PP(16'h6D7E,4);
TASK_PP(16'h6D7F,4);
TASK_PP(16'h6D80,4);
TASK_PP(16'h6D81,4);
TASK_PP(16'h6D82,4);
TASK_PP(16'h6D83,4);
TASK_PP(16'h6D84,4);
TASK_PP(16'h6D85,4);
TASK_PP(16'h6D86,4);
TASK_PP(16'h6D87,4);
TASK_PP(16'h6D88,4);
TASK_PP(16'h6D89,4);
TASK_PP(16'h6D8A,4);
TASK_PP(16'h6D8B,4);
TASK_PP(16'h6D8C,4);
TASK_PP(16'h6D8D,4);
TASK_PP(16'h6D8E,4);
TASK_PP(16'h6D8F,4);
TASK_PP(16'h6D90,4);
TASK_PP(16'h6D91,4);
TASK_PP(16'h6D92,4);
TASK_PP(16'h6D93,4);
TASK_PP(16'h6D94,4);
TASK_PP(16'h6D95,4);
TASK_PP(16'h6D96,4);
TASK_PP(16'h6D97,4);
TASK_PP(16'h6D98,4);
TASK_PP(16'h6D99,4);
TASK_PP(16'h6D9A,4);
TASK_PP(16'h6D9B,4);
TASK_PP(16'h6D9C,4);
TASK_PP(16'h6D9D,4);
TASK_PP(16'h6D9E,4);
TASK_PP(16'h6D9F,4);
TASK_PP(16'h6DA0,4);
TASK_PP(16'h6DA1,4);
TASK_PP(16'h6DA2,4);
TASK_PP(16'h6DA3,4);
TASK_PP(16'h6DA4,4);
TASK_PP(16'h6DA5,4);
TASK_PP(16'h6DA6,4);
TASK_PP(16'h6DA7,4);
TASK_PP(16'h6DA8,4);
TASK_PP(16'h6DA9,4);
TASK_PP(16'h6DAA,4);
TASK_PP(16'h6DAB,4);
TASK_PP(16'h6DAC,4);
TASK_PP(16'h6DAD,4);
TASK_PP(16'h6DAE,4);
TASK_PP(16'h6DAF,4);
TASK_PP(16'h6DB0,4);
TASK_PP(16'h6DB1,4);
TASK_PP(16'h6DB2,4);
TASK_PP(16'h6DB3,4);
TASK_PP(16'h6DB4,4);
TASK_PP(16'h6DB5,4);
TASK_PP(16'h6DB6,4);
TASK_PP(16'h6DB7,4);
TASK_PP(16'h6DB8,4);
TASK_PP(16'h6DB9,4);
TASK_PP(16'h6DBA,4);
TASK_PP(16'h6DBB,4);
TASK_PP(16'h6DBC,4);
TASK_PP(16'h6DBD,4);
TASK_PP(16'h6DBE,4);
TASK_PP(16'h6DBF,4);
TASK_PP(16'h6DC0,4);
TASK_PP(16'h6DC1,4);
TASK_PP(16'h6DC2,4);
TASK_PP(16'h6DC3,4);
TASK_PP(16'h6DC4,4);
TASK_PP(16'h6DC5,4);
TASK_PP(16'h6DC6,4);
TASK_PP(16'h6DC7,4);
TASK_PP(16'h6DC8,4);
TASK_PP(16'h6DC9,4);
TASK_PP(16'h6DCA,4);
TASK_PP(16'h6DCB,4);
TASK_PP(16'h6DCC,4);
TASK_PP(16'h6DCD,4);
TASK_PP(16'h6DCE,4);
TASK_PP(16'h6DCF,4);
TASK_PP(16'h6DD0,4);
TASK_PP(16'h6DD1,4);
TASK_PP(16'h6DD2,4);
TASK_PP(16'h6DD3,4);
TASK_PP(16'h6DD4,4);
TASK_PP(16'h6DD5,4);
TASK_PP(16'h6DD6,4);
TASK_PP(16'h6DD7,4);
TASK_PP(16'h6DD8,4);
TASK_PP(16'h6DD9,4);
TASK_PP(16'h6DDA,4);
TASK_PP(16'h6DDB,4);
TASK_PP(16'h6DDC,4);
TASK_PP(16'h6DDD,4);
TASK_PP(16'h6DDE,4);
TASK_PP(16'h6DDF,4);
TASK_PP(16'h6DE0,4);
TASK_PP(16'h6DE1,4);
TASK_PP(16'h6DE2,4);
TASK_PP(16'h6DE3,4);
TASK_PP(16'h6DE4,4);
TASK_PP(16'h6DE5,4);
TASK_PP(16'h6DE6,4);
TASK_PP(16'h6DE7,4);
TASK_PP(16'h6DE8,4);
TASK_PP(16'h6DE9,4);
TASK_PP(16'h6DEA,4);
TASK_PP(16'h6DEB,4);
TASK_PP(16'h6DEC,4);
TASK_PP(16'h6DED,4);
TASK_PP(16'h6DEE,4);
TASK_PP(16'h6DEF,4);
TASK_PP(16'h6DF0,4);
TASK_PP(16'h6DF1,4);
TASK_PP(16'h6DF2,4);
TASK_PP(16'h6DF3,4);
TASK_PP(16'h6DF4,4);
TASK_PP(16'h6DF5,4);
TASK_PP(16'h6DF6,4);
TASK_PP(16'h6DF7,4);
TASK_PP(16'h6DF8,4);
TASK_PP(16'h6DF9,4);
TASK_PP(16'h6DFA,4);
TASK_PP(16'h6DFB,4);
TASK_PP(16'h6DFC,4);
TASK_PP(16'h6DFD,4);
TASK_PP(16'h6DFE,4);
TASK_PP(16'h6DFF,4);
TASK_PP(16'h6E00,4);
TASK_PP(16'h6E01,4);
TASK_PP(16'h6E02,4);
TASK_PP(16'h6E03,4);
TASK_PP(16'h6E04,4);
TASK_PP(16'h6E05,4);
TASK_PP(16'h6E06,4);
TASK_PP(16'h6E07,4);
TASK_PP(16'h6E08,4);
TASK_PP(16'h6E09,4);
TASK_PP(16'h6E0A,4);
TASK_PP(16'h6E0B,4);
TASK_PP(16'h6E0C,4);
TASK_PP(16'h6E0D,4);
TASK_PP(16'h6E0E,4);
TASK_PP(16'h6E0F,4);
TASK_PP(16'h6E10,4);
TASK_PP(16'h6E11,4);
TASK_PP(16'h6E12,4);
TASK_PP(16'h6E13,4);
TASK_PP(16'h6E14,4);
TASK_PP(16'h6E15,4);
TASK_PP(16'h6E16,4);
TASK_PP(16'h6E17,4);
TASK_PP(16'h6E18,4);
TASK_PP(16'h6E19,4);
TASK_PP(16'h6E1A,4);
TASK_PP(16'h6E1B,4);
TASK_PP(16'h6E1C,4);
TASK_PP(16'h6E1D,4);
TASK_PP(16'h6E1E,4);
TASK_PP(16'h6E1F,4);
TASK_PP(16'h6E20,4);
TASK_PP(16'h6E21,4);
TASK_PP(16'h6E22,4);
TASK_PP(16'h6E23,4);
TASK_PP(16'h6E24,4);
TASK_PP(16'h6E25,4);
TASK_PP(16'h6E26,4);
TASK_PP(16'h6E27,4);
TASK_PP(16'h6E28,4);
TASK_PP(16'h6E29,4);
TASK_PP(16'h6E2A,4);
TASK_PP(16'h6E2B,4);
TASK_PP(16'h6E2C,4);
TASK_PP(16'h6E2D,4);
TASK_PP(16'h6E2E,4);
TASK_PP(16'h6E2F,4);
TASK_PP(16'h6E30,4);
TASK_PP(16'h6E31,4);
TASK_PP(16'h6E32,4);
TASK_PP(16'h6E33,4);
TASK_PP(16'h6E34,4);
TASK_PP(16'h6E35,4);
TASK_PP(16'h6E36,4);
TASK_PP(16'h6E37,4);
TASK_PP(16'h6E38,4);
TASK_PP(16'h6E39,4);
TASK_PP(16'h6E3A,4);
TASK_PP(16'h6E3B,4);
TASK_PP(16'h6E3C,4);
TASK_PP(16'h6E3D,4);
TASK_PP(16'h6E3E,4);
TASK_PP(16'h6E3F,4);
TASK_PP(16'h6E40,4);
TASK_PP(16'h6E41,4);
TASK_PP(16'h6E42,4);
TASK_PP(16'h6E43,4);
TASK_PP(16'h6E44,4);
TASK_PP(16'h6E45,4);
TASK_PP(16'h6E46,4);
TASK_PP(16'h6E47,4);
TASK_PP(16'h6E48,4);
TASK_PP(16'h6E49,4);
TASK_PP(16'h6E4A,4);
TASK_PP(16'h6E4B,4);
TASK_PP(16'h6E4C,4);
TASK_PP(16'h6E4D,4);
TASK_PP(16'h6E4E,4);
TASK_PP(16'h6E4F,4);
TASK_PP(16'h6E50,4);
TASK_PP(16'h6E51,4);
TASK_PP(16'h6E52,4);
TASK_PP(16'h6E53,4);
TASK_PP(16'h6E54,4);
TASK_PP(16'h6E55,4);
TASK_PP(16'h6E56,4);
TASK_PP(16'h6E57,4);
TASK_PP(16'h6E58,4);
TASK_PP(16'h6E59,4);
TASK_PP(16'h6E5A,4);
TASK_PP(16'h6E5B,4);
TASK_PP(16'h6E5C,4);
TASK_PP(16'h6E5D,4);
TASK_PP(16'h6E5E,4);
TASK_PP(16'h6E5F,4);
TASK_PP(16'h6E60,4);
TASK_PP(16'h6E61,4);
TASK_PP(16'h6E62,4);
TASK_PP(16'h6E63,4);
TASK_PP(16'h6E64,4);
TASK_PP(16'h6E65,4);
TASK_PP(16'h6E66,4);
TASK_PP(16'h6E67,4);
TASK_PP(16'h6E68,4);
TASK_PP(16'h6E69,4);
TASK_PP(16'h6E6A,4);
TASK_PP(16'h6E6B,4);
TASK_PP(16'h6E6C,4);
TASK_PP(16'h6E6D,4);
TASK_PP(16'h6E6E,4);
TASK_PP(16'h6E6F,4);
TASK_PP(16'h6E70,4);
TASK_PP(16'h6E71,4);
TASK_PP(16'h6E72,4);
TASK_PP(16'h6E73,4);
TASK_PP(16'h6E74,4);
TASK_PP(16'h6E75,4);
TASK_PP(16'h6E76,4);
TASK_PP(16'h6E77,4);
TASK_PP(16'h6E78,4);
TASK_PP(16'h6E79,4);
TASK_PP(16'h6E7A,4);
TASK_PP(16'h6E7B,4);
TASK_PP(16'h6E7C,4);
TASK_PP(16'h6E7D,4);
TASK_PP(16'h6E7E,4);
TASK_PP(16'h6E7F,4);
TASK_PP(16'h6E80,4);
TASK_PP(16'h6E81,4);
TASK_PP(16'h6E82,4);
TASK_PP(16'h6E83,4);
TASK_PP(16'h6E84,4);
TASK_PP(16'h6E85,4);
TASK_PP(16'h6E86,4);
TASK_PP(16'h6E87,4);
TASK_PP(16'h6E88,4);
TASK_PP(16'h6E89,4);
TASK_PP(16'h6E8A,4);
TASK_PP(16'h6E8B,4);
TASK_PP(16'h6E8C,4);
TASK_PP(16'h6E8D,4);
TASK_PP(16'h6E8E,4);
TASK_PP(16'h6E8F,4);
TASK_PP(16'h6E90,4);
TASK_PP(16'h6E91,4);
TASK_PP(16'h6E92,4);
TASK_PP(16'h6E93,4);
TASK_PP(16'h6E94,4);
TASK_PP(16'h6E95,4);
TASK_PP(16'h6E96,4);
TASK_PP(16'h6E97,4);
TASK_PP(16'h6E98,4);
TASK_PP(16'h6E99,4);
TASK_PP(16'h6E9A,4);
TASK_PP(16'h6E9B,4);
TASK_PP(16'h6E9C,4);
TASK_PP(16'h6E9D,4);
TASK_PP(16'h6E9E,4);
TASK_PP(16'h6E9F,4);
TASK_PP(16'h6EA0,4);
TASK_PP(16'h6EA1,4);
TASK_PP(16'h6EA2,4);
TASK_PP(16'h6EA3,4);
TASK_PP(16'h6EA4,4);
TASK_PP(16'h6EA5,4);
TASK_PP(16'h6EA6,4);
TASK_PP(16'h6EA7,4);
TASK_PP(16'h6EA8,4);
TASK_PP(16'h6EA9,4);
TASK_PP(16'h6EAA,4);
TASK_PP(16'h6EAB,4);
TASK_PP(16'h6EAC,4);
TASK_PP(16'h6EAD,4);
TASK_PP(16'h6EAE,4);
TASK_PP(16'h6EAF,4);
TASK_PP(16'h6EB0,4);
TASK_PP(16'h6EB1,4);
TASK_PP(16'h6EB2,4);
TASK_PP(16'h6EB3,4);
TASK_PP(16'h6EB4,4);
TASK_PP(16'h6EB5,4);
TASK_PP(16'h6EB6,4);
TASK_PP(16'h6EB7,4);
TASK_PP(16'h6EB8,4);
TASK_PP(16'h6EB9,4);
TASK_PP(16'h6EBA,4);
TASK_PP(16'h6EBB,4);
TASK_PP(16'h6EBC,4);
TASK_PP(16'h6EBD,4);
TASK_PP(16'h6EBE,4);
TASK_PP(16'h6EBF,4);
TASK_PP(16'h6EC0,4);
TASK_PP(16'h6EC1,4);
TASK_PP(16'h6EC2,4);
TASK_PP(16'h6EC3,4);
TASK_PP(16'h6EC4,4);
TASK_PP(16'h6EC5,4);
TASK_PP(16'h6EC6,4);
TASK_PP(16'h6EC7,4);
TASK_PP(16'h6EC8,4);
TASK_PP(16'h6EC9,4);
TASK_PP(16'h6ECA,4);
TASK_PP(16'h6ECB,4);
TASK_PP(16'h6ECC,4);
TASK_PP(16'h6ECD,4);
TASK_PP(16'h6ECE,4);
TASK_PP(16'h6ECF,4);
TASK_PP(16'h6ED0,4);
TASK_PP(16'h6ED1,4);
TASK_PP(16'h6ED2,4);
TASK_PP(16'h6ED3,4);
TASK_PP(16'h6ED4,4);
TASK_PP(16'h6ED5,4);
TASK_PP(16'h6ED6,4);
TASK_PP(16'h6ED7,4);
TASK_PP(16'h6ED8,4);
TASK_PP(16'h6ED9,4);
TASK_PP(16'h6EDA,4);
TASK_PP(16'h6EDB,4);
TASK_PP(16'h6EDC,4);
TASK_PP(16'h6EDD,4);
TASK_PP(16'h6EDE,4);
TASK_PP(16'h6EDF,4);
TASK_PP(16'h6EE0,4);
TASK_PP(16'h6EE1,4);
TASK_PP(16'h6EE2,4);
TASK_PP(16'h6EE3,4);
TASK_PP(16'h6EE4,4);
TASK_PP(16'h6EE5,4);
TASK_PP(16'h6EE6,4);
TASK_PP(16'h6EE7,4);
TASK_PP(16'h6EE8,4);
TASK_PP(16'h6EE9,4);
TASK_PP(16'h6EEA,4);
TASK_PP(16'h6EEB,4);
TASK_PP(16'h6EEC,4);
TASK_PP(16'h6EED,4);
TASK_PP(16'h6EEE,4);
TASK_PP(16'h6EEF,4);
TASK_PP(16'h6EF0,4);
TASK_PP(16'h6EF1,4);
TASK_PP(16'h6EF2,4);
TASK_PP(16'h6EF3,4);
TASK_PP(16'h6EF4,4);
TASK_PP(16'h6EF5,4);
TASK_PP(16'h6EF6,4);
TASK_PP(16'h6EF7,4);
TASK_PP(16'h6EF8,4);
TASK_PP(16'h6EF9,4);
TASK_PP(16'h6EFA,4);
TASK_PP(16'h6EFB,4);
TASK_PP(16'h6EFC,4);
TASK_PP(16'h6EFD,4);
TASK_PP(16'h6EFE,4);
TASK_PP(16'h6EFF,4);
TASK_PP(16'h6F00,4);
TASK_PP(16'h6F01,4);
TASK_PP(16'h6F02,4);
TASK_PP(16'h6F03,4);
TASK_PP(16'h6F04,4);
TASK_PP(16'h6F05,4);
TASK_PP(16'h6F06,4);
TASK_PP(16'h6F07,4);
TASK_PP(16'h6F08,4);
TASK_PP(16'h6F09,4);
TASK_PP(16'h6F0A,4);
TASK_PP(16'h6F0B,4);
TASK_PP(16'h6F0C,4);
TASK_PP(16'h6F0D,4);
TASK_PP(16'h6F0E,4);
TASK_PP(16'h6F0F,4);
TASK_PP(16'h6F10,4);
TASK_PP(16'h6F11,4);
TASK_PP(16'h6F12,4);
TASK_PP(16'h6F13,4);
TASK_PP(16'h6F14,4);
TASK_PP(16'h6F15,4);
TASK_PP(16'h6F16,4);
TASK_PP(16'h6F17,4);
TASK_PP(16'h6F18,4);
TASK_PP(16'h6F19,4);
TASK_PP(16'h6F1A,4);
TASK_PP(16'h6F1B,4);
TASK_PP(16'h6F1C,4);
TASK_PP(16'h6F1D,4);
TASK_PP(16'h6F1E,4);
TASK_PP(16'h6F1F,4);
TASK_PP(16'h6F20,4);
TASK_PP(16'h6F21,4);
TASK_PP(16'h6F22,4);
TASK_PP(16'h6F23,4);
TASK_PP(16'h6F24,4);
TASK_PP(16'h6F25,4);
TASK_PP(16'h6F26,4);
TASK_PP(16'h6F27,4);
TASK_PP(16'h6F28,4);
TASK_PP(16'h6F29,4);
TASK_PP(16'h6F2A,4);
TASK_PP(16'h6F2B,4);
TASK_PP(16'h6F2C,4);
TASK_PP(16'h6F2D,4);
TASK_PP(16'h6F2E,4);
TASK_PP(16'h6F2F,4);
TASK_PP(16'h6F30,4);
TASK_PP(16'h6F31,4);
TASK_PP(16'h6F32,4);
TASK_PP(16'h6F33,4);
TASK_PP(16'h6F34,4);
TASK_PP(16'h6F35,4);
TASK_PP(16'h6F36,4);
TASK_PP(16'h6F37,4);
TASK_PP(16'h6F38,4);
TASK_PP(16'h6F39,4);
TASK_PP(16'h6F3A,4);
TASK_PP(16'h6F3B,4);
TASK_PP(16'h6F3C,4);
TASK_PP(16'h6F3D,4);
TASK_PP(16'h6F3E,4);
TASK_PP(16'h6F3F,4);
TASK_PP(16'h6F40,4);
TASK_PP(16'h6F41,4);
TASK_PP(16'h6F42,4);
TASK_PP(16'h6F43,4);
TASK_PP(16'h6F44,4);
TASK_PP(16'h6F45,4);
TASK_PP(16'h6F46,4);
TASK_PP(16'h6F47,4);
TASK_PP(16'h6F48,4);
TASK_PP(16'h6F49,4);
TASK_PP(16'h6F4A,4);
TASK_PP(16'h6F4B,4);
TASK_PP(16'h6F4C,4);
TASK_PP(16'h6F4D,4);
TASK_PP(16'h6F4E,4);
TASK_PP(16'h6F4F,4);
TASK_PP(16'h6F50,4);
TASK_PP(16'h6F51,4);
TASK_PP(16'h6F52,4);
TASK_PP(16'h6F53,4);
TASK_PP(16'h6F54,4);
TASK_PP(16'h6F55,4);
TASK_PP(16'h6F56,4);
TASK_PP(16'h6F57,4);
TASK_PP(16'h6F58,4);
TASK_PP(16'h6F59,4);
TASK_PP(16'h6F5A,4);
TASK_PP(16'h6F5B,4);
TASK_PP(16'h6F5C,4);
TASK_PP(16'h6F5D,4);
TASK_PP(16'h6F5E,4);
TASK_PP(16'h6F5F,4);
TASK_PP(16'h6F60,4);
TASK_PP(16'h6F61,4);
TASK_PP(16'h6F62,4);
TASK_PP(16'h6F63,4);
TASK_PP(16'h6F64,4);
TASK_PP(16'h6F65,4);
TASK_PP(16'h6F66,4);
TASK_PP(16'h6F67,4);
TASK_PP(16'h6F68,4);
TASK_PP(16'h6F69,4);
TASK_PP(16'h6F6A,4);
TASK_PP(16'h6F6B,4);
TASK_PP(16'h6F6C,4);
TASK_PP(16'h6F6D,4);
TASK_PP(16'h6F6E,4);
TASK_PP(16'h6F6F,4);
TASK_PP(16'h6F70,4);
TASK_PP(16'h6F71,4);
TASK_PP(16'h6F72,4);
TASK_PP(16'h6F73,4);
TASK_PP(16'h6F74,4);
TASK_PP(16'h6F75,4);
TASK_PP(16'h6F76,4);
TASK_PP(16'h6F77,4);
TASK_PP(16'h6F78,4);
TASK_PP(16'h6F79,4);
TASK_PP(16'h6F7A,4);
TASK_PP(16'h6F7B,4);
TASK_PP(16'h6F7C,4);
TASK_PP(16'h6F7D,4);
TASK_PP(16'h6F7E,4);
TASK_PP(16'h6F7F,4);
TASK_PP(16'h6F80,4);
TASK_PP(16'h6F81,4);
TASK_PP(16'h6F82,4);
TASK_PP(16'h6F83,4);
TASK_PP(16'h6F84,4);
TASK_PP(16'h6F85,4);
TASK_PP(16'h6F86,4);
TASK_PP(16'h6F87,4);
TASK_PP(16'h6F88,4);
TASK_PP(16'h6F89,4);
TASK_PP(16'h6F8A,4);
TASK_PP(16'h6F8B,4);
TASK_PP(16'h6F8C,4);
TASK_PP(16'h6F8D,4);
TASK_PP(16'h6F8E,4);
TASK_PP(16'h6F8F,4);
TASK_PP(16'h6F90,4);
TASK_PP(16'h6F91,4);
TASK_PP(16'h6F92,4);
TASK_PP(16'h6F93,4);
TASK_PP(16'h6F94,4);
TASK_PP(16'h6F95,4);
TASK_PP(16'h6F96,4);
TASK_PP(16'h6F97,4);
TASK_PP(16'h6F98,4);
TASK_PP(16'h6F99,4);
TASK_PP(16'h6F9A,4);
TASK_PP(16'h6F9B,4);
TASK_PP(16'h6F9C,4);
TASK_PP(16'h6F9D,4);
TASK_PP(16'h6F9E,4);
TASK_PP(16'h6F9F,4);
TASK_PP(16'h6FA0,4);
TASK_PP(16'h6FA1,4);
TASK_PP(16'h6FA2,4);
TASK_PP(16'h6FA3,4);
TASK_PP(16'h6FA4,4);
TASK_PP(16'h6FA5,4);
TASK_PP(16'h6FA6,4);
TASK_PP(16'h6FA7,4);
TASK_PP(16'h6FA8,4);
TASK_PP(16'h6FA9,4);
TASK_PP(16'h6FAA,4);
TASK_PP(16'h6FAB,4);
TASK_PP(16'h6FAC,4);
TASK_PP(16'h6FAD,4);
TASK_PP(16'h6FAE,4);
TASK_PP(16'h6FAF,4);
TASK_PP(16'h6FB0,4);
TASK_PP(16'h6FB1,4);
TASK_PP(16'h6FB2,4);
TASK_PP(16'h6FB3,4);
TASK_PP(16'h6FB4,4);
TASK_PP(16'h6FB5,4);
TASK_PP(16'h6FB6,4);
TASK_PP(16'h6FB7,4);
TASK_PP(16'h6FB8,4);
TASK_PP(16'h6FB9,4);
TASK_PP(16'h6FBA,4);
TASK_PP(16'h6FBB,4);
TASK_PP(16'h6FBC,4);
TASK_PP(16'h6FBD,4);
TASK_PP(16'h6FBE,4);
TASK_PP(16'h6FBF,4);
TASK_PP(16'h6FC0,4);
TASK_PP(16'h6FC1,4);
TASK_PP(16'h6FC2,4);
TASK_PP(16'h6FC3,4);
TASK_PP(16'h6FC4,4);
TASK_PP(16'h6FC5,4);
TASK_PP(16'h6FC6,4);
TASK_PP(16'h6FC7,4);
TASK_PP(16'h6FC8,4);
TASK_PP(16'h6FC9,4);
TASK_PP(16'h6FCA,4);
TASK_PP(16'h6FCB,4);
TASK_PP(16'h6FCC,4);
TASK_PP(16'h6FCD,4);
TASK_PP(16'h6FCE,4);
TASK_PP(16'h6FCF,4);
TASK_PP(16'h6FD0,4);
TASK_PP(16'h6FD1,4);
TASK_PP(16'h6FD2,4);
TASK_PP(16'h6FD3,4);
TASK_PP(16'h6FD4,4);
TASK_PP(16'h6FD5,4);
TASK_PP(16'h6FD6,4);
TASK_PP(16'h6FD7,4);
TASK_PP(16'h6FD8,4);
TASK_PP(16'h6FD9,4);
TASK_PP(16'h6FDA,4);
TASK_PP(16'h6FDB,4);
TASK_PP(16'h6FDC,4);
TASK_PP(16'h6FDD,4);
TASK_PP(16'h6FDE,4);
TASK_PP(16'h6FDF,4);
TASK_PP(16'h6FE0,4);
TASK_PP(16'h6FE1,4);
TASK_PP(16'h6FE2,4);
TASK_PP(16'h6FE3,4);
TASK_PP(16'h6FE4,4);
TASK_PP(16'h6FE5,4);
TASK_PP(16'h6FE6,4);
TASK_PP(16'h6FE7,4);
TASK_PP(16'h6FE8,4);
TASK_PP(16'h6FE9,4);
TASK_PP(16'h6FEA,4);
TASK_PP(16'h6FEB,4);
TASK_PP(16'h6FEC,4);
TASK_PP(16'h6FED,4);
TASK_PP(16'h6FEE,4);
TASK_PP(16'h6FEF,4);
TASK_PP(16'h6FF0,4);
TASK_PP(16'h6FF1,4);
TASK_PP(16'h6FF2,4);
TASK_PP(16'h6FF3,4);
TASK_PP(16'h6FF4,4);
TASK_PP(16'h6FF5,4);
TASK_PP(16'h6FF6,4);
TASK_PP(16'h6FF7,4);
TASK_PP(16'h6FF8,4);
TASK_PP(16'h6FF9,4);
TASK_PP(16'h6FFA,4);
TASK_PP(16'h6FFB,4);
TASK_PP(16'h6FFC,4);
TASK_PP(16'h6FFD,4);
TASK_PP(16'h6FFE,4);
TASK_PP(16'h6FFF,4);
TASK_PP(16'h7000,4);
TASK_PP(16'h7001,4);
TASK_PP(16'h7002,4);
TASK_PP(16'h7003,4);
TASK_PP(16'h7004,4);
TASK_PP(16'h7005,4);
TASK_PP(16'h7006,4);
TASK_PP(16'h7007,4);
TASK_PP(16'h7008,4);
TASK_PP(16'h7009,4);
TASK_PP(16'h700A,4);
TASK_PP(16'h700B,4);
TASK_PP(16'h700C,4);
TASK_PP(16'h700D,4);
TASK_PP(16'h700E,4);
TASK_PP(16'h700F,4);
TASK_PP(16'h7010,4);
TASK_PP(16'h7011,4);
TASK_PP(16'h7012,4);
TASK_PP(16'h7013,4);
TASK_PP(16'h7014,4);
TASK_PP(16'h7015,4);
TASK_PP(16'h7016,4);
TASK_PP(16'h7017,4);
TASK_PP(16'h7018,4);
TASK_PP(16'h7019,4);
TASK_PP(16'h701A,4);
TASK_PP(16'h701B,4);
TASK_PP(16'h701C,4);
TASK_PP(16'h701D,4);
TASK_PP(16'h701E,4);
TASK_PP(16'h701F,4);
TASK_PP(16'h7020,4);
TASK_PP(16'h7021,4);
TASK_PP(16'h7022,4);
TASK_PP(16'h7023,4);
TASK_PP(16'h7024,4);
TASK_PP(16'h7025,4);
TASK_PP(16'h7026,4);
TASK_PP(16'h7027,4);
TASK_PP(16'h7028,4);
TASK_PP(16'h7029,4);
TASK_PP(16'h702A,4);
TASK_PP(16'h702B,4);
TASK_PP(16'h702C,4);
TASK_PP(16'h702D,4);
TASK_PP(16'h702E,4);
TASK_PP(16'h702F,4);
TASK_PP(16'h7030,4);
TASK_PP(16'h7031,4);
TASK_PP(16'h7032,4);
TASK_PP(16'h7033,4);
TASK_PP(16'h7034,4);
TASK_PP(16'h7035,4);
TASK_PP(16'h7036,4);
TASK_PP(16'h7037,4);
TASK_PP(16'h7038,4);
TASK_PP(16'h7039,4);
TASK_PP(16'h703A,4);
TASK_PP(16'h703B,4);
TASK_PP(16'h703C,4);
TASK_PP(16'h703D,4);
TASK_PP(16'h703E,4);
TASK_PP(16'h703F,4);
TASK_PP(16'h7040,4);
TASK_PP(16'h7041,4);
TASK_PP(16'h7042,4);
TASK_PP(16'h7043,4);
TASK_PP(16'h7044,4);
TASK_PP(16'h7045,4);
TASK_PP(16'h7046,4);
TASK_PP(16'h7047,4);
TASK_PP(16'h7048,4);
TASK_PP(16'h7049,4);
TASK_PP(16'h704A,4);
TASK_PP(16'h704B,4);
TASK_PP(16'h704C,4);
TASK_PP(16'h704D,4);
TASK_PP(16'h704E,4);
TASK_PP(16'h704F,4);
TASK_PP(16'h7050,4);
TASK_PP(16'h7051,4);
TASK_PP(16'h7052,4);
TASK_PP(16'h7053,4);
TASK_PP(16'h7054,4);
TASK_PP(16'h7055,4);
TASK_PP(16'h7056,4);
TASK_PP(16'h7057,4);
TASK_PP(16'h7058,4);
TASK_PP(16'h7059,4);
TASK_PP(16'h705A,4);
TASK_PP(16'h705B,4);
TASK_PP(16'h705C,4);
TASK_PP(16'h705D,4);
TASK_PP(16'h705E,4);
TASK_PP(16'h705F,4);
TASK_PP(16'h7060,4);
TASK_PP(16'h7061,4);
TASK_PP(16'h7062,4);
TASK_PP(16'h7063,4);
TASK_PP(16'h7064,4);
TASK_PP(16'h7065,4);
TASK_PP(16'h7066,4);
TASK_PP(16'h7067,4);
TASK_PP(16'h7068,4);
TASK_PP(16'h7069,4);
TASK_PP(16'h706A,4);
TASK_PP(16'h706B,4);
TASK_PP(16'h706C,4);
TASK_PP(16'h706D,4);
TASK_PP(16'h706E,4);
TASK_PP(16'h706F,4);
TASK_PP(16'h7070,4);
TASK_PP(16'h7071,4);
TASK_PP(16'h7072,4);
TASK_PP(16'h7073,4);
TASK_PP(16'h7074,4);
TASK_PP(16'h7075,4);
TASK_PP(16'h7076,4);
TASK_PP(16'h7077,4);
TASK_PP(16'h7078,4);
TASK_PP(16'h7079,4);
TASK_PP(16'h707A,4);
TASK_PP(16'h707B,4);
TASK_PP(16'h707C,4);
TASK_PP(16'h707D,4);
TASK_PP(16'h707E,4);
TASK_PP(16'h707F,4);
TASK_PP(16'h7080,4);
TASK_PP(16'h7081,4);
TASK_PP(16'h7082,4);
TASK_PP(16'h7083,4);
TASK_PP(16'h7084,4);
TASK_PP(16'h7085,4);
TASK_PP(16'h7086,4);
TASK_PP(16'h7087,4);
TASK_PP(16'h7088,4);
TASK_PP(16'h7089,4);
TASK_PP(16'h708A,4);
TASK_PP(16'h708B,4);
TASK_PP(16'h708C,4);
TASK_PP(16'h708D,4);
TASK_PP(16'h708E,4);
TASK_PP(16'h708F,4);
TASK_PP(16'h7090,4);
TASK_PP(16'h7091,4);
TASK_PP(16'h7092,4);
TASK_PP(16'h7093,4);
TASK_PP(16'h7094,4);
TASK_PP(16'h7095,4);
TASK_PP(16'h7096,4);
TASK_PP(16'h7097,4);
TASK_PP(16'h7098,4);
TASK_PP(16'h7099,4);
TASK_PP(16'h709A,4);
TASK_PP(16'h709B,4);
TASK_PP(16'h709C,4);
TASK_PP(16'h709D,4);
TASK_PP(16'h709E,4);
TASK_PP(16'h709F,4);
TASK_PP(16'h70A0,4);
TASK_PP(16'h70A1,4);
TASK_PP(16'h70A2,4);
TASK_PP(16'h70A3,4);
TASK_PP(16'h70A4,4);
TASK_PP(16'h70A5,4);
TASK_PP(16'h70A6,4);
TASK_PP(16'h70A7,4);
TASK_PP(16'h70A8,4);
TASK_PP(16'h70A9,4);
TASK_PP(16'h70AA,4);
TASK_PP(16'h70AB,4);
TASK_PP(16'h70AC,4);
TASK_PP(16'h70AD,4);
TASK_PP(16'h70AE,4);
TASK_PP(16'h70AF,4);
TASK_PP(16'h70B0,4);
TASK_PP(16'h70B1,4);
TASK_PP(16'h70B2,4);
TASK_PP(16'h70B3,4);
TASK_PP(16'h70B4,4);
TASK_PP(16'h70B5,4);
TASK_PP(16'h70B6,4);
TASK_PP(16'h70B7,4);
TASK_PP(16'h70B8,4);
TASK_PP(16'h70B9,4);
TASK_PP(16'h70BA,4);
TASK_PP(16'h70BB,4);
TASK_PP(16'h70BC,4);
TASK_PP(16'h70BD,4);
TASK_PP(16'h70BE,4);
TASK_PP(16'h70BF,4);
TASK_PP(16'h70C0,4);
TASK_PP(16'h70C1,4);
TASK_PP(16'h70C2,4);
TASK_PP(16'h70C3,4);
TASK_PP(16'h70C4,4);
TASK_PP(16'h70C5,4);
TASK_PP(16'h70C6,4);
TASK_PP(16'h70C7,4);
TASK_PP(16'h70C8,4);
TASK_PP(16'h70C9,4);
TASK_PP(16'h70CA,4);
TASK_PP(16'h70CB,4);
TASK_PP(16'h70CC,4);
TASK_PP(16'h70CD,4);
TASK_PP(16'h70CE,4);
TASK_PP(16'h70CF,4);
TASK_PP(16'h70D0,4);
TASK_PP(16'h70D1,4);
TASK_PP(16'h70D2,4);
TASK_PP(16'h70D3,4);
TASK_PP(16'h70D4,4);
TASK_PP(16'h70D5,4);
TASK_PP(16'h70D6,4);
TASK_PP(16'h70D7,4);
TASK_PP(16'h70D8,4);
TASK_PP(16'h70D9,4);
TASK_PP(16'h70DA,4);
TASK_PP(16'h70DB,4);
TASK_PP(16'h70DC,4);
TASK_PP(16'h70DD,4);
TASK_PP(16'h70DE,4);
TASK_PP(16'h70DF,4);
TASK_PP(16'h70E0,4);
TASK_PP(16'h70E1,4);
TASK_PP(16'h70E2,4);
TASK_PP(16'h70E3,4);
TASK_PP(16'h70E4,4);
TASK_PP(16'h70E5,4);
TASK_PP(16'h70E6,4);
TASK_PP(16'h70E7,4);
TASK_PP(16'h70E8,4);
TASK_PP(16'h70E9,4);
TASK_PP(16'h70EA,4);
TASK_PP(16'h70EB,4);
TASK_PP(16'h70EC,4);
TASK_PP(16'h70ED,4);
TASK_PP(16'h70EE,4);
TASK_PP(16'h70EF,4);
TASK_PP(16'h70F0,4);
TASK_PP(16'h70F1,4);
TASK_PP(16'h70F2,4);
TASK_PP(16'h70F3,4);
TASK_PP(16'h70F4,4);
TASK_PP(16'h70F5,4);
TASK_PP(16'h70F6,4);
TASK_PP(16'h70F7,4);
TASK_PP(16'h70F8,4);
TASK_PP(16'h70F9,4);
TASK_PP(16'h70FA,4);
TASK_PP(16'h70FB,4);
TASK_PP(16'h70FC,4);
TASK_PP(16'h70FD,4);
TASK_PP(16'h70FE,4);
TASK_PP(16'h70FF,4);
TASK_PP(16'h7100,4);
TASK_PP(16'h7101,4);
TASK_PP(16'h7102,4);
TASK_PP(16'h7103,4);
TASK_PP(16'h7104,4);
TASK_PP(16'h7105,4);
TASK_PP(16'h7106,4);
TASK_PP(16'h7107,4);
TASK_PP(16'h7108,4);
TASK_PP(16'h7109,4);
TASK_PP(16'h710A,4);
TASK_PP(16'h710B,4);
TASK_PP(16'h710C,4);
TASK_PP(16'h710D,4);
TASK_PP(16'h710E,4);
TASK_PP(16'h710F,4);
TASK_PP(16'h7110,4);
TASK_PP(16'h7111,4);
TASK_PP(16'h7112,4);
TASK_PP(16'h7113,4);
TASK_PP(16'h7114,4);
TASK_PP(16'h7115,4);
TASK_PP(16'h7116,4);
TASK_PP(16'h7117,4);
TASK_PP(16'h7118,4);
TASK_PP(16'h7119,4);
TASK_PP(16'h711A,4);
TASK_PP(16'h711B,4);
TASK_PP(16'h711C,4);
TASK_PP(16'h711D,4);
TASK_PP(16'h711E,4);
TASK_PP(16'h711F,4);
TASK_PP(16'h7120,4);
TASK_PP(16'h7121,4);
TASK_PP(16'h7122,4);
TASK_PP(16'h7123,4);
TASK_PP(16'h7124,4);
TASK_PP(16'h7125,4);
TASK_PP(16'h7126,4);
TASK_PP(16'h7127,4);
TASK_PP(16'h7128,4);
TASK_PP(16'h7129,4);
TASK_PP(16'h712A,4);
TASK_PP(16'h712B,4);
TASK_PP(16'h712C,4);
TASK_PP(16'h712D,4);
TASK_PP(16'h712E,4);
TASK_PP(16'h712F,4);
TASK_PP(16'h7130,4);
TASK_PP(16'h7131,4);
TASK_PP(16'h7132,4);
TASK_PP(16'h7133,4);
TASK_PP(16'h7134,4);
TASK_PP(16'h7135,4);
TASK_PP(16'h7136,4);
TASK_PP(16'h7137,4);
TASK_PP(16'h7138,4);
TASK_PP(16'h7139,4);
TASK_PP(16'h713A,4);
TASK_PP(16'h713B,4);
TASK_PP(16'h713C,4);
TASK_PP(16'h713D,4);
TASK_PP(16'h713E,4);
TASK_PP(16'h713F,4);
TASK_PP(16'h7140,4);
TASK_PP(16'h7141,4);
TASK_PP(16'h7142,4);
TASK_PP(16'h7143,4);
TASK_PP(16'h7144,4);
TASK_PP(16'h7145,4);
TASK_PP(16'h7146,4);
TASK_PP(16'h7147,4);
TASK_PP(16'h7148,4);
TASK_PP(16'h7149,4);
TASK_PP(16'h714A,4);
TASK_PP(16'h714B,4);
TASK_PP(16'h714C,4);
TASK_PP(16'h714D,4);
TASK_PP(16'h714E,4);
TASK_PP(16'h714F,4);
TASK_PP(16'h7150,4);
TASK_PP(16'h7151,4);
TASK_PP(16'h7152,4);
TASK_PP(16'h7153,4);
TASK_PP(16'h7154,4);
TASK_PP(16'h7155,4);
TASK_PP(16'h7156,4);
TASK_PP(16'h7157,4);
TASK_PP(16'h7158,4);
TASK_PP(16'h7159,4);
TASK_PP(16'h715A,4);
TASK_PP(16'h715B,4);
TASK_PP(16'h715C,4);
TASK_PP(16'h715D,4);
TASK_PP(16'h715E,4);
TASK_PP(16'h715F,4);
TASK_PP(16'h7160,4);
TASK_PP(16'h7161,4);
TASK_PP(16'h7162,4);
TASK_PP(16'h7163,4);
TASK_PP(16'h7164,4);
TASK_PP(16'h7165,4);
TASK_PP(16'h7166,4);
TASK_PP(16'h7167,4);
TASK_PP(16'h7168,4);
TASK_PP(16'h7169,4);
TASK_PP(16'h716A,4);
TASK_PP(16'h716B,4);
TASK_PP(16'h716C,4);
TASK_PP(16'h716D,4);
TASK_PP(16'h716E,4);
TASK_PP(16'h716F,4);
TASK_PP(16'h7170,4);
TASK_PP(16'h7171,4);
TASK_PP(16'h7172,4);
TASK_PP(16'h7173,4);
TASK_PP(16'h7174,4);
TASK_PP(16'h7175,4);
TASK_PP(16'h7176,4);
TASK_PP(16'h7177,4);
TASK_PP(16'h7178,4);
TASK_PP(16'h7179,4);
TASK_PP(16'h717A,4);
TASK_PP(16'h717B,4);
TASK_PP(16'h717C,4);
TASK_PP(16'h717D,4);
TASK_PP(16'h717E,4);
TASK_PP(16'h717F,4);
TASK_PP(16'h7180,4);
TASK_PP(16'h7181,4);
TASK_PP(16'h7182,4);
TASK_PP(16'h7183,4);
TASK_PP(16'h7184,4);
TASK_PP(16'h7185,4);
TASK_PP(16'h7186,4);
TASK_PP(16'h7187,4);
TASK_PP(16'h7188,4);
TASK_PP(16'h7189,4);
TASK_PP(16'h718A,4);
TASK_PP(16'h718B,4);
TASK_PP(16'h718C,4);
TASK_PP(16'h718D,4);
TASK_PP(16'h718E,4);
TASK_PP(16'h718F,4);
TASK_PP(16'h7190,4);
TASK_PP(16'h7191,4);
TASK_PP(16'h7192,4);
TASK_PP(16'h7193,4);
TASK_PP(16'h7194,4);
TASK_PP(16'h7195,4);
TASK_PP(16'h7196,4);
TASK_PP(16'h7197,4);
TASK_PP(16'h7198,4);
TASK_PP(16'h7199,4);
TASK_PP(16'h719A,4);
TASK_PP(16'h719B,4);
TASK_PP(16'h719C,4);
TASK_PP(16'h719D,4);
TASK_PP(16'h719E,4);
TASK_PP(16'h719F,4);
TASK_PP(16'h71A0,4);
TASK_PP(16'h71A1,4);
TASK_PP(16'h71A2,4);
TASK_PP(16'h71A3,4);
TASK_PP(16'h71A4,4);
TASK_PP(16'h71A5,4);
TASK_PP(16'h71A6,4);
TASK_PP(16'h71A7,4);
TASK_PP(16'h71A8,4);
TASK_PP(16'h71A9,4);
TASK_PP(16'h71AA,4);
TASK_PP(16'h71AB,4);
TASK_PP(16'h71AC,4);
TASK_PP(16'h71AD,4);
TASK_PP(16'h71AE,4);
TASK_PP(16'h71AF,4);
TASK_PP(16'h71B0,4);
TASK_PP(16'h71B1,4);
TASK_PP(16'h71B2,4);
TASK_PP(16'h71B3,4);
TASK_PP(16'h71B4,4);
TASK_PP(16'h71B5,4);
TASK_PP(16'h71B6,4);
TASK_PP(16'h71B7,4);
TASK_PP(16'h71B8,4);
TASK_PP(16'h71B9,4);
TASK_PP(16'h71BA,4);
TASK_PP(16'h71BB,4);
TASK_PP(16'h71BC,4);
TASK_PP(16'h71BD,4);
TASK_PP(16'h71BE,4);
TASK_PP(16'h71BF,4);
TASK_PP(16'h71C0,4);
TASK_PP(16'h71C1,4);
TASK_PP(16'h71C2,4);
TASK_PP(16'h71C3,4);
TASK_PP(16'h71C4,4);
TASK_PP(16'h71C5,4);
TASK_PP(16'h71C6,4);
TASK_PP(16'h71C7,4);
TASK_PP(16'h71C8,4);
TASK_PP(16'h71C9,4);
TASK_PP(16'h71CA,4);
TASK_PP(16'h71CB,4);
TASK_PP(16'h71CC,4);
TASK_PP(16'h71CD,4);
TASK_PP(16'h71CE,4);
TASK_PP(16'h71CF,4);
TASK_PP(16'h71D0,4);
TASK_PP(16'h71D1,4);
TASK_PP(16'h71D2,4);
TASK_PP(16'h71D3,4);
TASK_PP(16'h71D4,4);
TASK_PP(16'h71D5,4);
TASK_PP(16'h71D6,4);
TASK_PP(16'h71D7,4);
TASK_PP(16'h71D8,4);
TASK_PP(16'h71D9,4);
TASK_PP(16'h71DA,4);
TASK_PP(16'h71DB,4);
TASK_PP(16'h71DC,4);
TASK_PP(16'h71DD,4);
TASK_PP(16'h71DE,4);
TASK_PP(16'h71DF,4);
TASK_PP(16'h71E0,4);
TASK_PP(16'h71E1,4);
TASK_PP(16'h71E2,4);
TASK_PP(16'h71E3,4);
TASK_PP(16'h71E4,4);
TASK_PP(16'h71E5,4);
TASK_PP(16'h71E6,4);
TASK_PP(16'h71E7,4);
TASK_PP(16'h71E8,4);
TASK_PP(16'h71E9,4);
TASK_PP(16'h71EA,4);
TASK_PP(16'h71EB,4);
TASK_PP(16'h71EC,4);
TASK_PP(16'h71ED,4);
TASK_PP(16'h71EE,4);
TASK_PP(16'h71EF,4);
TASK_PP(16'h71F0,4);
TASK_PP(16'h71F1,4);
TASK_PP(16'h71F2,4);
TASK_PP(16'h71F3,4);
TASK_PP(16'h71F4,4);
TASK_PP(16'h71F5,4);
TASK_PP(16'h71F6,4);
TASK_PP(16'h71F7,4);
TASK_PP(16'h71F8,4);
TASK_PP(16'h71F9,4);
TASK_PP(16'h71FA,4);
TASK_PP(16'h71FB,4);
TASK_PP(16'h71FC,4);
TASK_PP(16'h71FD,4);
TASK_PP(16'h71FE,4);
TASK_PP(16'h71FF,4);
TASK_PP(16'h7200,4);
TASK_PP(16'h7201,4);
TASK_PP(16'h7202,4);
TASK_PP(16'h7203,4);
TASK_PP(16'h7204,4);
TASK_PP(16'h7205,4);
TASK_PP(16'h7206,4);
TASK_PP(16'h7207,4);
TASK_PP(16'h7208,4);
TASK_PP(16'h7209,4);
TASK_PP(16'h720A,4);
TASK_PP(16'h720B,4);
TASK_PP(16'h720C,4);
TASK_PP(16'h720D,4);
TASK_PP(16'h720E,4);
TASK_PP(16'h720F,4);
TASK_PP(16'h7210,4);
TASK_PP(16'h7211,4);
TASK_PP(16'h7212,4);
TASK_PP(16'h7213,4);
TASK_PP(16'h7214,4);
TASK_PP(16'h7215,4);
TASK_PP(16'h7216,4);
TASK_PP(16'h7217,4);
TASK_PP(16'h7218,4);
TASK_PP(16'h7219,4);
TASK_PP(16'h721A,4);
TASK_PP(16'h721B,4);
TASK_PP(16'h721C,4);
TASK_PP(16'h721D,4);
TASK_PP(16'h721E,4);
TASK_PP(16'h721F,4);
TASK_PP(16'h7220,4);
TASK_PP(16'h7221,4);
TASK_PP(16'h7222,4);
TASK_PP(16'h7223,4);
TASK_PP(16'h7224,4);
TASK_PP(16'h7225,4);
TASK_PP(16'h7226,4);
TASK_PP(16'h7227,4);
TASK_PP(16'h7228,4);
TASK_PP(16'h7229,4);
TASK_PP(16'h722A,4);
TASK_PP(16'h722B,4);
TASK_PP(16'h722C,4);
TASK_PP(16'h722D,4);
TASK_PP(16'h722E,4);
TASK_PP(16'h722F,4);
TASK_PP(16'h7230,4);
TASK_PP(16'h7231,4);
TASK_PP(16'h7232,4);
TASK_PP(16'h7233,4);
TASK_PP(16'h7234,4);
TASK_PP(16'h7235,4);
TASK_PP(16'h7236,4);
TASK_PP(16'h7237,4);
TASK_PP(16'h7238,4);
TASK_PP(16'h7239,4);
TASK_PP(16'h723A,4);
TASK_PP(16'h723B,4);
TASK_PP(16'h723C,4);
TASK_PP(16'h723D,4);
TASK_PP(16'h723E,4);
TASK_PP(16'h723F,4);
TASK_PP(16'h7240,4);
TASK_PP(16'h7241,4);
TASK_PP(16'h7242,4);
TASK_PP(16'h7243,4);
TASK_PP(16'h7244,4);
TASK_PP(16'h7245,4);
TASK_PP(16'h7246,4);
TASK_PP(16'h7247,4);
TASK_PP(16'h7248,4);
TASK_PP(16'h7249,4);
TASK_PP(16'h724A,4);
TASK_PP(16'h724B,4);
TASK_PP(16'h724C,4);
TASK_PP(16'h724D,4);
TASK_PP(16'h724E,4);
TASK_PP(16'h724F,4);
TASK_PP(16'h7250,4);
TASK_PP(16'h7251,4);
TASK_PP(16'h7252,4);
TASK_PP(16'h7253,4);
TASK_PP(16'h7254,4);
TASK_PP(16'h7255,4);
TASK_PP(16'h7256,4);
TASK_PP(16'h7257,4);
TASK_PP(16'h7258,4);
TASK_PP(16'h7259,4);
TASK_PP(16'h725A,4);
TASK_PP(16'h725B,4);
TASK_PP(16'h725C,4);
TASK_PP(16'h725D,4);
TASK_PP(16'h725E,4);
TASK_PP(16'h725F,4);
TASK_PP(16'h7260,4);
TASK_PP(16'h7261,4);
TASK_PP(16'h7262,4);
TASK_PP(16'h7263,4);
TASK_PP(16'h7264,4);
TASK_PP(16'h7265,4);
TASK_PP(16'h7266,4);
TASK_PP(16'h7267,4);
TASK_PP(16'h7268,4);
TASK_PP(16'h7269,4);
TASK_PP(16'h726A,4);
TASK_PP(16'h726B,4);
TASK_PP(16'h726C,4);
TASK_PP(16'h726D,4);
TASK_PP(16'h726E,4);
TASK_PP(16'h726F,4);
TASK_PP(16'h7270,4);
TASK_PP(16'h7271,4);
TASK_PP(16'h7272,4);
TASK_PP(16'h7273,4);
TASK_PP(16'h7274,4);
TASK_PP(16'h7275,4);
TASK_PP(16'h7276,4);
TASK_PP(16'h7277,4);
TASK_PP(16'h7278,4);
TASK_PP(16'h7279,4);
TASK_PP(16'h727A,4);
TASK_PP(16'h727B,4);
TASK_PP(16'h727C,4);
TASK_PP(16'h727D,4);
TASK_PP(16'h727E,4);
TASK_PP(16'h727F,4);
TASK_PP(16'h7280,4);
TASK_PP(16'h7281,4);
TASK_PP(16'h7282,4);
TASK_PP(16'h7283,4);
TASK_PP(16'h7284,4);
TASK_PP(16'h7285,4);
TASK_PP(16'h7286,4);
TASK_PP(16'h7287,4);
TASK_PP(16'h7288,4);
TASK_PP(16'h7289,4);
TASK_PP(16'h728A,4);
TASK_PP(16'h728B,4);
TASK_PP(16'h728C,4);
TASK_PP(16'h728D,4);
TASK_PP(16'h728E,4);
TASK_PP(16'h728F,4);
TASK_PP(16'h7290,4);
TASK_PP(16'h7291,4);
TASK_PP(16'h7292,4);
TASK_PP(16'h7293,4);
TASK_PP(16'h7294,4);
TASK_PP(16'h7295,4);
TASK_PP(16'h7296,4);
TASK_PP(16'h7297,4);
TASK_PP(16'h7298,4);
TASK_PP(16'h7299,4);
TASK_PP(16'h729A,4);
TASK_PP(16'h729B,4);
TASK_PP(16'h729C,4);
TASK_PP(16'h729D,4);
TASK_PP(16'h729E,4);
TASK_PP(16'h729F,4);
TASK_PP(16'h72A0,4);
TASK_PP(16'h72A1,4);
TASK_PP(16'h72A2,4);
TASK_PP(16'h72A3,4);
TASK_PP(16'h72A4,4);
TASK_PP(16'h72A5,4);
TASK_PP(16'h72A6,4);
TASK_PP(16'h72A7,4);
TASK_PP(16'h72A8,4);
TASK_PP(16'h72A9,4);
TASK_PP(16'h72AA,4);
TASK_PP(16'h72AB,4);
TASK_PP(16'h72AC,4);
TASK_PP(16'h72AD,4);
TASK_PP(16'h72AE,4);
TASK_PP(16'h72AF,4);
TASK_PP(16'h72B0,4);
TASK_PP(16'h72B1,4);
TASK_PP(16'h72B2,4);
TASK_PP(16'h72B3,4);
TASK_PP(16'h72B4,4);
TASK_PP(16'h72B5,4);
TASK_PP(16'h72B6,4);
TASK_PP(16'h72B7,4);
TASK_PP(16'h72B8,4);
TASK_PP(16'h72B9,4);
TASK_PP(16'h72BA,4);
TASK_PP(16'h72BB,4);
TASK_PP(16'h72BC,4);
TASK_PP(16'h72BD,4);
TASK_PP(16'h72BE,4);
TASK_PP(16'h72BF,4);
TASK_PP(16'h72C0,4);
TASK_PP(16'h72C1,4);
TASK_PP(16'h72C2,4);
TASK_PP(16'h72C3,4);
TASK_PP(16'h72C4,4);
TASK_PP(16'h72C5,4);
TASK_PP(16'h72C6,4);
TASK_PP(16'h72C7,4);
TASK_PP(16'h72C8,4);
TASK_PP(16'h72C9,4);
TASK_PP(16'h72CA,4);
TASK_PP(16'h72CB,4);
TASK_PP(16'h72CC,4);
TASK_PP(16'h72CD,4);
TASK_PP(16'h72CE,4);
TASK_PP(16'h72CF,4);
TASK_PP(16'h72D0,4);
TASK_PP(16'h72D1,4);
TASK_PP(16'h72D2,4);
TASK_PP(16'h72D3,4);
TASK_PP(16'h72D4,4);
TASK_PP(16'h72D5,4);
TASK_PP(16'h72D6,4);
TASK_PP(16'h72D7,4);
TASK_PP(16'h72D8,4);
TASK_PP(16'h72D9,4);
TASK_PP(16'h72DA,4);
TASK_PP(16'h72DB,4);
TASK_PP(16'h72DC,4);
TASK_PP(16'h72DD,4);
TASK_PP(16'h72DE,4);
TASK_PP(16'h72DF,4);
TASK_PP(16'h72E0,4);
TASK_PP(16'h72E1,4);
TASK_PP(16'h72E2,4);
TASK_PP(16'h72E3,4);
TASK_PP(16'h72E4,4);
TASK_PP(16'h72E5,4);
TASK_PP(16'h72E6,4);
TASK_PP(16'h72E7,4);
TASK_PP(16'h72E8,4);
TASK_PP(16'h72E9,4);
TASK_PP(16'h72EA,4);
TASK_PP(16'h72EB,4);
TASK_PP(16'h72EC,4);
TASK_PP(16'h72ED,4);
TASK_PP(16'h72EE,4);
TASK_PP(16'h72EF,4);
TASK_PP(16'h72F0,4);
TASK_PP(16'h72F1,4);
TASK_PP(16'h72F2,4);
TASK_PP(16'h72F3,4);
TASK_PP(16'h72F4,4);
TASK_PP(16'h72F5,4);
TASK_PP(16'h72F6,4);
TASK_PP(16'h72F7,4);
TASK_PP(16'h72F8,4);
TASK_PP(16'h72F9,4);
TASK_PP(16'h72FA,4);
TASK_PP(16'h72FB,4);
TASK_PP(16'h72FC,4);
TASK_PP(16'h72FD,4);
TASK_PP(16'h72FE,4);
TASK_PP(16'h72FF,4);
TASK_PP(16'h7300,4);
TASK_PP(16'h7301,4);
TASK_PP(16'h7302,4);
TASK_PP(16'h7303,4);
TASK_PP(16'h7304,4);
TASK_PP(16'h7305,4);
TASK_PP(16'h7306,4);
TASK_PP(16'h7307,4);
TASK_PP(16'h7308,4);
TASK_PP(16'h7309,4);
TASK_PP(16'h730A,4);
TASK_PP(16'h730B,4);
TASK_PP(16'h730C,4);
TASK_PP(16'h730D,4);
TASK_PP(16'h730E,4);
TASK_PP(16'h730F,4);
TASK_PP(16'h7310,4);
TASK_PP(16'h7311,4);
TASK_PP(16'h7312,4);
TASK_PP(16'h7313,4);
TASK_PP(16'h7314,4);
TASK_PP(16'h7315,4);
TASK_PP(16'h7316,4);
TASK_PP(16'h7317,4);
TASK_PP(16'h7318,4);
TASK_PP(16'h7319,4);
TASK_PP(16'h731A,4);
TASK_PP(16'h731B,4);
TASK_PP(16'h731C,4);
TASK_PP(16'h731D,4);
TASK_PP(16'h731E,4);
TASK_PP(16'h731F,4);
TASK_PP(16'h7320,4);
TASK_PP(16'h7321,4);
TASK_PP(16'h7322,4);
TASK_PP(16'h7323,4);
TASK_PP(16'h7324,4);
TASK_PP(16'h7325,4);
TASK_PP(16'h7326,4);
TASK_PP(16'h7327,4);
TASK_PP(16'h7328,4);
TASK_PP(16'h7329,4);
TASK_PP(16'h732A,4);
TASK_PP(16'h732B,4);
TASK_PP(16'h732C,4);
TASK_PP(16'h732D,4);
TASK_PP(16'h732E,4);
TASK_PP(16'h732F,4);
TASK_PP(16'h7330,4);
TASK_PP(16'h7331,4);
TASK_PP(16'h7332,4);
TASK_PP(16'h7333,4);
TASK_PP(16'h7334,4);
TASK_PP(16'h7335,4);
TASK_PP(16'h7336,4);
TASK_PP(16'h7337,4);
TASK_PP(16'h7338,4);
TASK_PP(16'h7339,4);
TASK_PP(16'h733A,4);
TASK_PP(16'h733B,4);
TASK_PP(16'h733C,4);
TASK_PP(16'h733D,4);
TASK_PP(16'h733E,4);
TASK_PP(16'h733F,4);
TASK_PP(16'h7340,4);
TASK_PP(16'h7341,4);
TASK_PP(16'h7342,4);
TASK_PP(16'h7343,4);
TASK_PP(16'h7344,4);
TASK_PP(16'h7345,4);
TASK_PP(16'h7346,4);
TASK_PP(16'h7347,4);
TASK_PP(16'h7348,4);
TASK_PP(16'h7349,4);
TASK_PP(16'h734A,4);
TASK_PP(16'h734B,4);
TASK_PP(16'h734C,4);
TASK_PP(16'h734D,4);
TASK_PP(16'h734E,4);
TASK_PP(16'h734F,4);
TASK_PP(16'h7350,4);
TASK_PP(16'h7351,4);
TASK_PP(16'h7352,4);
TASK_PP(16'h7353,4);
TASK_PP(16'h7354,4);
TASK_PP(16'h7355,4);
TASK_PP(16'h7356,4);
TASK_PP(16'h7357,4);
TASK_PP(16'h7358,4);
TASK_PP(16'h7359,4);
TASK_PP(16'h735A,4);
TASK_PP(16'h735B,4);
TASK_PP(16'h735C,4);
TASK_PP(16'h735D,4);
TASK_PP(16'h735E,4);
TASK_PP(16'h735F,4);
TASK_PP(16'h7360,4);
TASK_PP(16'h7361,4);
TASK_PP(16'h7362,4);
TASK_PP(16'h7363,4);
TASK_PP(16'h7364,4);
TASK_PP(16'h7365,4);
TASK_PP(16'h7366,4);
TASK_PP(16'h7367,4);
TASK_PP(16'h7368,4);
TASK_PP(16'h7369,4);
TASK_PP(16'h736A,4);
TASK_PP(16'h736B,4);
TASK_PP(16'h736C,4);
TASK_PP(16'h736D,4);
TASK_PP(16'h736E,4);
TASK_PP(16'h736F,4);
TASK_PP(16'h7370,4);
TASK_PP(16'h7371,4);
TASK_PP(16'h7372,4);
TASK_PP(16'h7373,4);
TASK_PP(16'h7374,4);
TASK_PP(16'h7375,4);
TASK_PP(16'h7376,4);
TASK_PP(16'h7377,4);
TASK_PP(16'h7378,4);
TASK_PP(16'h7379,4);
TASK_PP(16'h737A,4);
TASK_PP(16'h737B,4);
TASK_PP(16'h737C,4);
TASK_PP(16'h737D,4);
TASK_PP(16'h737E,4);
TASK_PP(16'h737F,4);
TASK_PP(16'h7380,4);
TASK_PP(16'h7381,4);
TASK_PP(16'h7382,4);
TASK_PP(16'h7383,4);
TASK_PP(16'h7384,4);
TASK_PP(16'h7385,4);
TASK_PP(16'h7386,4);
TASK_PP(16'h7387,4);
TASK_PP(16'h7388,4);
TASK_PP(16'h7389,4);
TASK_PP(16'h738A,4);
TASK_PP(16'h738B,4);
TASK_PP(16'h738C,4);
TASK_PP(16'h738D,4);
TASK_PP(16'h738E,4);
TASK_PP(16'h738F,4);
TASK_PP(16'h7390,4);
TASK_PP(16'h7391,4);
TASK_PP(16'h7392,4);
TASK_PP(16'h7393,4);
TASK_PP(16'h7394,4);
TASK_PP(16'h7395,4);
TASK_PP(16'h7396,4);
TASK_PP(16'h7397,4);
TASK_PP(16'h7398,4);
TASK_PP(16'h7399,4);
TASK_PP(16'h739A,4);
TASK_PP(16'h739B,4);
TASK_PP(16'h739C,4);
TASK_PP(16'h739D,4);
TASK_PP(16'h739E,4);
TASK_PP(16'h739F,4);
TASK_PP(16'h73A0,4);
TASK_PP(16'h73A1,4);
TASK_PP(16'h73A2,4);
TASK_PP(16'h73A3,4);
TASK_PP(16'h73A4,4);
TASK_PP(16'h73A5,4);
TASK_PP(16'h73A6,4);
TASK_PP(16'h73A7,4);
TASK_PP(16'h73A8,4);
TASK_PP(16'h73A9,4);
TASK_PP(16'h73AA,4);
TASK_PP(16'h73AB,4);
TASK_PP(16'h73AC,4);
TASK_PP(16'h73AD,4);
TASK_PP(16'h73AE,4);
TASK_PP(16'h73AF,4);
TASK_PP(16'h73B0,4);
TASK_PP(16'h73B1,4);
TASK_PP(16'h73B2,4);
TASK_PP(16'h73B3,4);
TASK_PP(16'h73B4,4);
TASK_PP(16'h73B5,4);
TASK_PP(16'h73B6,4);
TASK_PP(16'h73B7,4);
TASK_PP(16'h73B8,4);
TASK_PP(16'h73B9,4);
TASK_PP(16'h73BA,4);
TASK_PP(16'h73BB,4);
TASK_PP(16'h73BC,4);
TASK_PP(16'h73BD,4);
TASK_PP(16'h73BE,4);
TASK_PP(16'h73BF,4);
TASK_PP(16'h73C0,4);
TASK_PP(16'h73C1,4);
TASK_PP(16'h73C2,4);
TASK_PP(16'h73C3,4);
TASK_PP(16'h73C4,4);
TASK_PP(16'h73C5,4);
TASK_PP(16'h73C6,4);
TASK_PP(16'h73C7,4);
TASK_PP(16'h73C8,4);
TASK_PP(16'h73C9,4);
TASK_PP(16'h73CA,4);
TASK_PP(16'h73CB,4);
TASK_PP(16'h73CC,4);
TASK_PP(16'h73CD,4);
TASK_PP(16'h73CE,4);
TASK_PP(16'h73CF,4);
TASK_PP(16'h73D0,4);
TASK_PP(16'h73D1,4);
TASK_PP(16'h73D2,4);
TASK_PP(16'h73D3,4);
TASK_PP(16'h73D4,4);
TASK_PP(16'h73D5,4);
TASK_PP(16'h73D6,4);
TASK_PP(16'h73D7,4);
TASK_PP(16'h73D8,4);
TASK_PP(16'h73D9,4);
TASK_PP(16'h73DA,4);
TASK_PP(16'h73DB,4);
TASK_PP(16'h73DC,4);
TASK_PP(16'h73DD,4);
TASK_PP(16'h73DE,4);
TASK_PP(16'h73DF,4);
TASK_PP(16'h73E0,4);
TASK_PP(16'h73E1,4);
TASK_PP(16'h73E2,4);
TASK_PP(16'h73E3,4);
TASK_PP(16'h73E4,4);
TASK_PP(16'h73E5,4);
TASK_PP(16'h73E6,4);
TASK_PP(16'h73E7,4);
TASK_PP(16'h73E8,4);
TASK_PP(16'h73E9,4);
TASK_PP(16'h73EA,4);
TASK_PP(16'h73EB,4);
TASK_PP(16'h73EC,4);
TASK_PP(16'h73ED,4);
TASK_PP(16'h73EE,4);
TASK_PP(16'h73EF,4);
TASK_PP(16'h73F0,4);
TASK_PP(16'h73F1,4);
TASK_PP(16'h73F2,4);
TASK_PP(16'h73F3,4);
TASK_PP(16'h73F4,4);
TASK_PP(16'h73F5,4);
TASK_PP(16'h73F6,4);
TASK_PP(16'h73F7,4);
TASK_PP(16'h73F8,4);
TASK_PP(16'h73F9,4);
TASK_PP(16'h73FA,4);
TASK_PP(16'h73FB,4);
TASK_PP(16'h73FC,4);
TASK_PP(16'h73FD,4);
TASK_PP(16'h73FE,4);
TASK_PP(16'h73FF,4);
TASK_PP(16'h7400,4);
TASK_PP(16'h7401,4);
TASK_PP(16'h7402,4);
TASK_PP(16'h7403,4);
TASK_PP(16'h7404,4);
TASK_PP(16'h7405,4);
TASK_PP(16'h7406,4);
TASK_PP(16'h7407,4);
TASK_PP(16'h7408,4);
TASK_PP(16'h7409,4);
TASK_PP(16'h740A,4);
TASK_PP(16'h740B,4);
TASK_PP(16'h740C,4);
TASK_PP(16'h740D,4);
TASK_PP(16'h740E,4);
TASK_PP(16'h740F,4);
TASK_PP(16'h7410,4);
TASK_PP(16'h7411,4);
TASK_PP(16'h7412,4);
TASK_PP(16'h7413,4);
TASK_PP(16'h7414,4);
TASK_PP(16'h7415,4);
TASK_PP(16'h7416,4);
TASK_PP(16'h7417,4);
TASK_PP(16'h7418,4);
TASK_PP(16'h7419,4);
TASK_PP(16'h741A,4);
TASK_PP(16'h741B,4);
TASK_PP(16'h741C,4);
TASK_PP(16'h741D,4);
TASK_PP(16'h741E,4);
TASK_PP(16'h741F,4);
TASK_PP(16'h7420,4);
TASK_PP(16'h7421,4);
TASK_PP(16'h7422,4);
TASK_PP(16'h7423,4);
TASK_PP(16'h7424,4);
TASK_PP(16'h7425,4);
TASK_PP(16'h7426,4);
TASK_PP(16'h7427,4);
TASK_PP(16'h7428,4);
TASK_PP(16'h7429,4);
TASK_PP(16'h742A,4);
TASK_PP(16'h742B,4);
TASK_PP(16'h742C,4);
TASK_PP(16'h742D,4);
TASK_PP(16'h742E,4);
TASK_PP(16'h742F,4);
TASK_PP(16'h7430,4);
TASK_PP(16'h7431,4);
TASK_PP(16'h7432,4);
TASK_PP(16'h7433,4);
TASK_PP(16'h7434,4);
TASK_PP(16'h7435,4);
TASK_PP(16'h7436,4);
TASK_PP(16'h7437,4);
TASK_PP(16'h7438,4);
TASK_PP(16'h7439,4);
TASK_PP(16'h743A,4);
TASK_PP(16'h743B,4);
TASK_PP(16'h743C,4);
TASK_PP(16'h743D,4);
TASK_PP(16'h743E,4);
TASK_PP(16'h743F,4);
TASK_PP(16'h7440,4);
TASK_PP(16'h7441,4);
TASK_PP(16'h7442,4);
TASK_PP(16'h7443,4);
TASK_PP(16'h7444,4);
TASK_PP(16'h7445,4);
TASK_PP(16'h7446,4);
TASK_PP(16'h7447,4);
TASK_PP(16'h7448,4);
TASK_PP(16'h7449,4);
TASK_PP(16'h744A,4);
TASK_PP(16'h744B,4);
TASK_PP(16'h744C,4);
TASK_PP(16'h744D,4);
TASK_PP(16'h744E,4);
TASK_PP(16'h744F,4);
TASK_PP(16'h7450,4);
TASK_PP(16'h7451,4);
TASK_PP(16'h7452,4);
TASK_PP(16'h7453,4);
TASK_PP(16'h7454,4);
TASK_PP(16'h7455,4);
TASK_PP(16'h7456,4);
TASK_PP(16'h7457,4);
TASK_PP(16'h7458,4);
TASK_PP(16'h7459,4);
TASK_PP(16'h745A,4);
TASK_PP(16'h745B,4);
TASK_PP(16'h745C,4);
TASK_PP(16'h745D,4);
TASK_PP(16'h745E,4);
TASK_PP(16'h745F,4);
TASK_PP(16'h7460,4);
TASK_PP(16'h7461,4);
TASK_PP(16'h7462,4);
TASK_PP(16'h7463,4);
TASK_PP(16'h7464,4);
TASK_PP(16'h7465,4);
TASK_PP(16'h7466,4);
TASK_PP(16'h7467,4);
TASK_PP(16'h7468,4);
TASK_PP(16'h7469,4);
TASK_PP(16'h746A,4);
TASK_PP(16'h746B,4);
TASK_PP(16'h746C,4);
TASK_PP(16'h746D,4);
TASK_PP(16'h746E,4);
TASK_PP(16'h746F,4);
TASK_PP(16'h7470,4);
TASK_PP(16'h7471,4);
TASK_PP(16'h7472,4);
TASK_PP(16'h7473,4);
TASK_PP(16'h7474,4);
TASK_PP(16'h7475,4);
TASK_PP(16'h7476,4);
TASK_PP(16'h7477,4);
TASK_PP(16'h7478,4);
TASK_PP(16'h7479,4);
TASK_PP(16'h747A,4);
TASK_PP(16'h747B,4);
TASK_PP(16'h747C,4);
TASK_PP(16'h747D,4);
TASK_PP(16'h747E,4);
TASK_PP(16'h747F,4);
TASK_PP(16'h7480,4);
TASK_PP(16'h7481,4);
TASK_PP(16'h7482,4);
TASK_PP(16'h7483,4);
TASK_PP(16'h7484,4);
TASK_PP(16'h7485,4);
TASK_PP(16'h7486,4);
TASK_PP(16'h7487,4);
TASK_PP(16'h7488,4);
TASK_PP(16'h7489,4);
TASK_PP(16'h748A,4);
TASK_PP(16'h748B,4);
TASK_PP(16'h748C,4);
TASK_PP(16'h748D,4);
TASK_PP(16'h748E,4);
TASK_PP(16'h748F,4);
TASK_PP(16'h7490,4);
TASK_PP(16'h7491,4);
TASK_PP(16'h7492,4);
TASK_PP(16'h7493,4);
TASK_PP(16'h7494,4);
TASK_PP(16'h7495,4);
TASK_PP(16'h7496,4);
TASK_PP(16'h7497,4);
TASK_PP(16'h7498,4);
TASK_PP(16'h7499,4);
TASK_PP(16'h749A,4);
TASK_PP(16'h749B,4);
TASK_PP(16'h749C,4);
TASK_PP(16'h749D,4);
TASK_PP(16'h749E,4);
TASK_PP(16'h749F,4);
TASK_PP(16'h74A0,4);
TASK_PP(16'h74A1,4);
TASK_PP(16'h74A2,4);
TASK_PP(16'h74A3,4);
TASK_PP(16'h74A4,4);
TASK_PP(16'h74A5,4);
TASK_PP(16'h74A6,4);
TASK_PP(16'h74A7,4);
TASK_PP(16'h74A8,4);
TASK_PP(16'h74A9,4);
TASK_PP(16'h74AA,4);
TASK_PP(16'h74AB,4);
TASK_PP(16'h74AC,4);
TASK_PP(16'h74AD,4);
TASK_PP(16'h74AE,4);
TASK_PP(16'h74AF,4);
TASK_PP(16'h74B0,4);
TASK_PP(16'h74B1,4);
TASK_PP(16'h74B2,4);
TASK_PP(16'h74B3,4);
TASK_PP(16'h74B4,4);
TASK_PP(16'h74B5,4);
TASK_PP(16'h74B6,4);
TASK_PP(16'h74B7,4);
TASK_PP(16'h74B8,4);
TASK_PP(16'h74B9,4);
TASK_PP(16'h74BA,4);
TASK_PP(16'h74BB,4);
TASK_PP(16'h74BC,4);
TASK_PP(16'h74BD,4);
TASK_PP(16'h74BE,4);
TASK_PP(16'h74BF,4);
TASK_PP(16'h74C0,4);
TASK_PP(16'h74C1,4);
TASK_PP(16'h74C2,4);
TASK_PP(16'h74C3,4);
TASK_PP(16'h74C4,4);
TASK_PP(16'h74C5,4);
TASK_PP(16'h74C6,4);
TASK_PP(16'h74C7,4);
TASK_PP(16'h74C8,4);
TASK_PP(16'h74C9,4);
TASK_PP(16'h74CA,4);
TASK_PP(16'h74CB,4);
TASK_PP(16'h74CC,4);
TASK_PP(16'h74CD,4);
TASK_PP(16'h74CE,4);
TASK_PP(16'h74CF,4);
TASK_PP(16'h74D0,4);
TASK_PP(16'h74D1,4);
TASK_PP(16'h74D2,4);
TASK_PP(16'h74D3,4);
TASK_PP(16'h74D4,4);
TASK_PP(16'h74D5,4);
TASK_PP(16'h74D6,4);
TASK_PP(16'h74D7,4);
TASK_PP(16'h74D8,4);
TASK_PP(16'h74D9,4);
TASK_PP(16'h74DA,4);
TASK_PP(16'h74DB,4);
TASK_PP(16'h74DC,4);
TASK_PP(16'h74DD,4);
TASK_PP(16'h74DE,4);
TASK_PP(16'h74DF,4);
TASK_PP(16'h74E0,4);
TASK_PP(16'h74E1,4);
TASK_PP(16'h74E2,4);
TASK_PP(16'h74E3,4);
TASK_PP(16'h74E4,4);
TASK_PP(16'h74E5,4);
TASK_PP(16'h74E6,4);
TASK_PP(16'h74E7,4);
TASK_PP(16'h74E8,4);
TASK_PP(16'h74E9,4);
TASK_PP(16'h74EA,4);
TASK_PP(16'h74EB,4);
TASK_PP(16'h74EC,4);
TASK_PP(16'h74ED,4);
TASK_PP(16'h74EE,4);
TASK_PP(16'h74EF,4);
TASK_PP(16'h74F0,4);
TASK_PP(16'h74F1,4);
TASK_PP(16'h74F2,4);
TASK_PP(16'h74F3,4);
TASK_PP(16'h74F4,4);
TASK_PP(16'h74F5,4);
TASK_PP(16'h74F6,4);
TASK_PP(16'h74F7,4);
TASK_PP(16'h74F8,4);
TASK_PP(16'h74F9,4);
TASK_PP(16'h74FA,4);
TASK_PP(16'h74FB,4);
TASK_PP(16'h74FC,4);
TASK_PP(16'h74FD,4);
TASK_PP(16'h74FE,4);
TASK_PP(16'h74FF,4);
TASK_PP(16'h7500,4);
TASK_PP(16'h7501,4);
TASK_PP(16'h7502,4);
TASK_PP(16'h7503,4);
TASK_PP(16'h7504,4);
TASK_PP(16'h7505,4);
TASK_PP(16'h7506,4);
TASK_PP(16'h7507,4);
TASK_PP(16'h7508,4);
TASK_PP(16'h7509,4);
TASK_PP(16'h750A,4);
TASK_PP(16'h750B,4);
TASK_PP(16'h750C,4);
TASK_PP(16'h750D,4);
TASK_PP(16'h750E,4);
TASK_PP(16'h750F,4);
TASK_PP(16'h7510,4);
TASK_PP(16'h7511,4);
TASK_PP(16'h7512,4);
TASK_PP(16'h7513,4);
TASK_PP(16'h7514,4);
TASK_PP(16'h7515,4);
TASK_PP(16'h7516,4);
TASK_PP(16'h7517,4);
TASK_PP(16'h7518,4);
TASK_PP(16'h7519,4);
TASK_PP(16'h751A,4);
TASK_PP(16'h751B,4);
TASK_PP(16'h751C,4);
TASK_PP(16'h751D,4);
TASK_PP(16'h751E,4);
TASK_PP(16'h751F,4);
TASK_PP(16'h7520,4);
TASK_PP(16'h7521,4);
TASK_PP(16'h7522,4);
TASK_PP(16'h7523,4);
TASK_PP(16'h7524,4);
TASK_PP(16'h7525,4);
TASK_PP(16'h7526,4);
TASK_PP(16'h7527,4);
TASK_PP(16'h7528,4);
TASK_PP(16'h7529,4);
TASK_PP(16'h752A,4);
TASK_PP(16'h752B,4);
TASK_PP(16'h752C,4);
TASK_PP(16'h752D,4);
TASK_PP(16'h752E,4);
TASK_PP(16'h752F,4);
TASK_PP(16'h7530,4);
TASK_PP(16'h7531,4);
TASK_PP(16'h7532,4);
TASK_PP(16'h7533,4);
TASK_PP(16'h7534,4);
TASK_PP(16'h7535,4);
TASK_PP(16'h7536,4);
TASK_PP(16'h7537,4);
TASK_PP(16'h7538,4);
TASK_PP(16'h7539,4);
TASK_PP(16'h753A,4);
TASK_PP(16'h753B,4);
TASK_PP(16'h753C,4);
TASK_PP(16'h753D,4);
TASK_PP(16'h753E,4);
TASK_PP(16'h753F,4);
TASK_PP(16'h7540,4);
TASK_PP(16'h7541,4);
TASK_PP(16'h7542,4);
TASK_PP(16'h7543,4);
TASK_PP(16'h7544,4);
TASK_PP(16'h7545,4);
TASK_PP(16'h7546,4);
TASK_PP(16'h7547,4);
TASK_PP(16'h7548,4);
TASK_PP(16'h7549,4);
TASK_PP(16'h754A,4);
TASK_PP(16'h754B,4);
TASK_PP(16'h754C,4);
TASK_PP(16'h754D,4);
TASK_PP(16'h754E,4);
TASK_PP(16'h754F,4);
TASK_PP(16'h7550,4);
TASK_PP(16'h7551,4);
TASK_PP(16'h7552,4);
TASK_PP(16'h7553,4);
TASK_PP(16'h7554,4);
TASK_PP(16'h7555,4);
TASK_PP(16'h7556,4);
TASK_PP(16'h7557,4);
TASK_PP(16'h7558,4);
TASK_PP(16'h7559,4);
TASK_PP(16'h755A,4);
TASK_PP(16'h755B,4);
TASK_PP(16'h755C,4);
TASK_PP(16'h755D,4);
TASK_PP(16'h755E,4);
TASK_PP(16'h755F,4);
TASK_PP(16'h7560,4);
TASK_PP(16'h7561,4);
TASK_PP(16'h7562,4);
TASK_PP(16'h7563,4);
TASK_PP(16'h7564,4);
TASK_PP(16'h7565,4);
TASK_PP(16'h7566,4);
TASK_PP(16'h7567,4);
TASK_PP(16'h7568,4);
TASK_PP(16'h7569,4);
TASK_PP(16'h756A,4);
TASK_PP(16'h756B,4);
TASK_PP(16'h756C,4);
TASK_PP(16'h756D,4);
TASK_PP(16'h756E,4);
TASK_PP(16'h756F,4);
TASK_PP(16'h7570,4);
TASK_PP(16'h7571,4);
TASK_PP(16'h7572,4);
TASK_PP(16'h7573,4);
TASK_PP(16'h7574,4);
TASK_PP(16'h7575,4);
TASK_PP(16'h7576,4);
TASK_PP(16'h7577,4);
TASK_PP(16'h7578,4);
TASK_PP(16'h7579,4);
TASK_PP(16'h757A,4);
TASK_PP(16'h757B,4);
TASK_PP(16'h757C,4);
TASK_PP(16'h757D,4);
TASK_PP(16'h757E,4);
TASK_PP(16'h757F,4);
TASK_PP(16'h7580,4);
TASK_PP(16'h7581,4);
TASK_PP(16'h7582,4);
TASK_PP(16'h7583,4);
TASK_PP(16'h7584,4);
TASK_PP(16'h7585,4);
TASK_PP(16'h7586,4);
TASK_PP(16'h7587,4);
TASK_PP(16'h7588,4);
TASK_PP(16'h7589,4);
TASK_PP(16'h758A,4);
TASK_PP(16'h758B,4);
TASK_PP(16'h758C,4);
TASK_PP(16'h758D,4);
TASK_PP(16'h758E,4);
TASK_PP(16'h758F,4);
TASK_PP(16'h7590,4);
TASK_PP(16'h7591,4);
TASK_PP(16'h7592,4);
TASK_PP(16'h7593,4);
TASK_PP(16'h7594,4);
TASK_PP(16'h7595,4);
TASK_PP(16'h7596,4);
TASK_PP(16'h7597,4);
TASK_PP(16'h7598,4);
TASK_PP(16'h7599,4);
TASK_PP(16'h759A,4);
TASK_PP(16'h759B,4);
TASK_PP(16'h759C,4);
TASK_PP(16'h759D,4);
TASK_PP(16'h759E,4);
TASK_PP(16'h759F,4);
TASK_PP(16'h75A0,4);
TASK_PP(16'h75A1,4);
TASK_PP(16'h75A2,4);
TASK_PP(16'h75A3,4);
TASK_PP(16'h75A4,4);
TASK_PP(16'h75A5,4);
TASK_PP(16'h75A6,4);
TASK_PP(16'h75A7,4);
TASK_PP(16'h75A8,4);
TASK_PP(16'h75A9,4);
TASK_PP(16'h75AA,4);
TASK_PP(16'h75AB,4);
TASK_PP(16'h75AC,4);
TASK_PP(16'h75AD,4);
TASK_PP(16'h75AE,4);
TASK_PP(16'h75AF,4);
TASK_PP(16'h75B0,4);
TASK_PP(16'h75B1,4);
TASK_PP(16'h75B2,4);
TASK_PP(16'h75B3,4);
TASK_PP(16'h75B4,4);
TASK_PP(16'h75B5,4);
TASK_PP(16'h75B6,4);
TASK_PP(16'h75B7,4);
TASK_PP(16'h75B8,4);
TASK_PP(16'h75B9,4);
TASK_PP(16'h75BA,4);
TASK_PP(16'h75BB,4);
TASK_PP(16'h75BC,4);
TASK_PP(16'h75BD,4);
TASK_PP(16'h75BE,4);
TASK_PP(16'h75BF,4);
TASK_PP(16'h75C0,4);
TASK_PP(16'h75C1,4);
TASK_PP(16'h75C2,4);
TASK_PP(16'h75C3,4);
TASK_PP(16'h75C4,4);
TASK_PP(16'h75C5,4);
TASK_PP(16'h75C6,4);
TASK_PP(16'h75C7,4);
TASK_PP(16'h75C8,4);
TASK_PP(16'h75C9,4);
TASK_PP(16'h75CA,4);
TASK_PP(16'h75CB,4);
TASK_PP(16'h75CC,4);
TASK_PP(16'h75CD,4);
TASK_PP(16'h75CE,4);
TASK_PP(16'h75CF,4);
TASK_PP(16'h75D0,4);
TASK_PP(16'h75D1,4);
TASK_PP(16'h75D2,4);
TASK_PP(16'h75D3,4);
TASK_PP(16'h75D4,4);
TASK_PP(16'h75D5,4);
TASK_PP(16'h75D6,4);
TASK_PP(16'h75D7,4);
TASK_PP(16'h75D8,4);
TASK_PP(16'h75D9,4);
TASK_PP(16'h75DA,4);
TASK_PP(16'h75DB,4);
TASK_PP(16'h75DC,4);
TASK_PP(16'h75DD,4);
TASK_PP(16'h75DE,4);
TASK_PP(16'h75DF,4);
TASK_PP(16'h75E0,4);
TASK_PP(16'h75E1,4);
TASK_PP(16'h75E2,4);
TASK_PP(16'h75E3,4);
TASK_PP(16'h75E4,4);
TASK_PP(16'h75E5,4);
TASK_PP(16'h75E6,4);
TASK_PP(16'h75E7,4);
TASK_PP(16'h75E8,4);
TASK_PP(16'h75E9,4);
TASK_PP(16'h75EA,4);
TASK_PP(16'h75EB,4);
TASK_PP(16'h75EC,4);
TASK_PP(16'h75ED,4);
TASK_PP(16'h75EE,4);
TASK_PP(16'h75EF,4);
TASK_PP(16'h75F0,4);
TASK_PP(16'h75F1,4);
TASK_PP(16'h75F2,4);
TASK_PP(16'h75F3,4);
TASK_PP(16'h75F4,4);
TASK_PP(16'h75F5,4);
TASK_PP(16'h75F6,4);
TASK_PP(16'h75F7,4);
TASK_PP(16'h75F8,4);
TASK_PP(16'h75F9,4);
TASK_PP(16'h75FA,4);
TASK_PP(16'h75FB,4);
TASK_PP(16'h75FC,4);
TASK_PP(16'h75FD,4);
TASK_PP(16'h75FE,4);
TASK_PP(16'h75FF,4);
TASK_PP(16'h7600,4);
TASK_PP(16'h7601,4);
TASK_PP(16'h7602,4);
TASK_PP(16'h7603,4);
TASK_PP(16'h7604,4);
TASK_PP(16'h7605,4);
TASK_PP(16'h7606,4);
TASK_PP(16'h7607,4);
TASK_PP(16'h7608,4);
TASK_PP(16'h7609,4);
TASK_PP(16'h760A,4);
TASK_PP(16'h760B,4);
TASK_PP(16'h760C,4);
TASK_PP(16'h760D,4);
TASK_PP(16'h760E,4);
TASK_PP(16'h760F,4);
TASK_PP(16'h7610,4);
TASK_PP(16'h7611,4);
TASK_PP(16'h7612,4);
TASK_PP(16'h7613,4);
TASK_PP(16'h7614,4);
TASK_PP(16'h7615,4);
TASK_PP(16'h7616,4);
TASK_PP(16'h7617,4);
TASK_PP(16'h7618,4);
TASK_PP(16'h7619,4);
TASK_PP(16'h761A,4);
TASK_PP(16'h761B,4);
TASK_PP(16'h761C,4);
TASK_PP(16'h761D,4);
TASK_PP(16'h761E,4);
TASK_PP(16'h761F,4);
TASK_PP(16'h7620,4);
TASK_PP(16'h7621,4);
TASK_PP(16'h7622,4);
TASK_PP(16'h7623,4);
TASK_PP(16'h7624,4);
TASK_PP(16'h7625,4);
TASK_PP(16'h7626,4);
TASK_PP(16'h7627,4);
TASK_PP(16'h7628,4);
TASK_PP(16'h7629,4);
TASK_PP(16'h762A,4);
TASK_PP(16'h762B,4);
TASK_PP(16'h762C,4);
TASK_PP(16'h762D,4);
TASK_PP(16'h762E,4);
TASK_PP(16'h762F,4);
TASK_PP(16'h7630,4);
TASK_PP(16'h7631,4);
TASK_PP(16'h7632,4);
TASK_PP(16'h7633,4);
TASK_PP(16'h7634,4);
TASK_PP(16'h7635,4);
TASK_PP(16'h7636,4);
TASK_PP(16'h7637,4);
TASK_PP(16'h7638,4);
TASK_PP(16'h7639,4);
TASK_PP(16'h763A,4);
TASK_PP(16'h763B,4);
TASK_PP(16'h763C,4);
TASK_PP(16'h763D,4);
TASK_PP(16'h763E,4);
TASK_PP(16'h763F,4);
TASK_PP(16'h7640,4);
TASK_PP(16'h7641,4);
TASK_PP(16'h7642,4);
TASK_PP(16'h7643,4);
TASK_PP(16'h7644,4);
TASK_PP(16'h7645,4);
TASK_PP(16'h7646,4);
TASK_PP(16'h7647,4);
TASK_PP(16'h7648,4);
TASK_PP(16'h7649,4);
TASK_PP(16'h764A,4);
TASK_PP(16'h764B,4);
TASK_PP(16'h764C,4);
TASK_PP(16'h764D,4);
TASK_PP(16'h764E,4);
TASK_PP(16'h764F,4);
TASK_PP(16'h7650,4);
TASK_PP(16'h7651,4);
TASK_PP(16'h7652,4);
TASK_PP(16'h7653,4);
TASK_PP(16'h7654,4);
TASK_PP(16'h7655,4);
TASK_PP(16'h7656,4);
TASK_PP(16'h7657,4);
TASK_PP(16'h7658,4);
TASK_PP(16'h7659,4);
TASK_PP(16'h765A,4);
TASK_PP(16'h765B,4);
TASK_PP(16'h765C,4);
TASK_PP(16'h765D,4);
TASK_PP(16'h765E,4);
TASK_PP(16'h765F,4);
TASK_PP(16'h7660,4);
TASK_PP(16'h7661,4);
TASK_PP(16'h7662,4);
TASK_PP(16'h7663,4);
TASK_PP(16'h7664,4);
TASK_PP(16'h7665,4);
TASK_PP(16'h7666,4);
TASK_PP(16'h7667,4);
TASK_PP(16'h7668,4);
TASK_PP(16'h7669,4);
TASK_PP(16'h766A,4);
TASK_PP(16'h766B,4);
TASK_PP(16'h766C,4);
TASK_PP(16'h766D,4);
TASK_PP(16'h766E,4);
TASK_PP(16'h766F,4);
TASK_PP(16'h7670,4);
TASK_PP(16'h7671,4);
TASK_PP(16'h7672,4);
TASK_PP(16'h7673,4);
TASK_PP(16'h7674,4);
TASK_PP(16'h7675,4);
TASK_PP(16'h7676,4);
TASK_PP(16'h7677,4);
TASK_PP(16'h7678,4);
TASK_PP(16'h7679,4);
TASK_PP(16'h767A,4);
TASK_PP(16'h767B,4);
TASK_PP(16'h767C,4);
TASK_PP(16'h767D,4);
TASK_PP(16'h767E,4);
TASK_PP(16'h767F,4);
TASK_PP(16'h7680,4);
TASK_PP(16'h7681,4);
TASK_PP(16'h7682,4);
TASK_PP(16'h7683,4);
TASK_PP(16'h7684,4);
TASK_PP(16'h7685,4);
TASK_PP(16'h7686,4);
TASK_PP(16'h7687,4);
TASK_PP(16'h7688,4);
TASK_PP(16'h7689,4);
TASK_PP(16'h768A,4);
TASK_PP(16'h768B,4);
TASK_PP(16'h768C,4);
TASK_PP(16'h768D,4);
TASK_PP(16'h768E,4);
TASK_PP(16'h768F,4);
TASK_PP(16'h7690,4);
TASK_PP(16'h7691,4);
TASK_PP(16'h7692,4);
TASK_PP(16'h7693,4);
TASK_PP(16'h7694,4);
TASK_PP(16'h7695,4);
TASK_PP(16'h7696,4);
TASK_PP(16'h7697,4);
TASK_PP(16'h7698,4);
TASK_PP(16'h7699,4);
TASK_PP(16'h769A,4);
TASK_PP(16'h769B,4);
TASK_PP(16'h769C,4);
TASK_PP(16'h769D,4);
TASK_PP(16'h769E,4);
TASK_PP(16'h769F,4);
TASK_PP(16'h76A0,4);
TASK_PP(16'h76A1,4);
TASK_PP(16'h76A2,4);
TASK_PP(16'h76A3,4);
TASK_PP(16'h76A4,4);
TASK_PP(16'h76A5,4);
TASK_PP(16'h76A6,4);
TASK_PP(16'h76A7,4);
TASK_PP(16'h76A8,4);
TASK_PP(16'h76A9,4);
TASK_PP(16'h76AA,4);
TASK_PP(16'h76AB,4);
TASK_PP(16'h76AC,4);
TASK_PP(16'h76AD,4);
TASK_PP(16'h76AE,4);
TASK_PP(16'h76AF,4);
TASK_PP(16'h76B0,4);
TASK_PP(16'h76B1,4);
TASK_PP(16'h76B2,4);
TASK_PP(16'h76B3,4);
TASK_PP(16'h76B4,4);
TASK_PP(16'h76B5,4);
TASK_PP(16'h76B6,4);
TASK_PP(16'h76B7,4);
TASK_PP(16'h76B8,4);
TASK_PP(16'h76B9,4);
TASK_PP(16'h76BA,4);
TASK_PP(16'h76BB,4);
TASK_PP(16'h76BC,4);
TASK_PP(16'h76BD,4);
TASK_PP(16'h76BE,4);
TASK_PP(16'h76BF,4);
TASK_PP(16'h76C0,4);
TASK_PP(16'h76C1,4);
TASK_PP(16'h76C2,4);
TASK_PP(16'h76C3,4);
TASK_PP(16'h76C4,4);
TASK_PP(16'h76C5,4);
TASK_PP(16'h76C6,4);
TASK_PP(16'h76C7,4);
TASK_PP(16'h76C8,4);
TASK_PP(16'h76C9,4);
TASK_PP(16'h76CA,4);
TASK_PP(16'h76CB,4);
TASK_PP(16'h76CC,4);
TASK_PP(16'h76CD,4);
TASK_PP(16'h76CE,4);
TASK_PP(16'h76CF,4);
TASK_PP(16'h76D0,4);
TASK_PP(16'h76D1,4);
TASK_PP(16'h76D2,4);
TASK_PP(16'h76D3,4);
TASK_PP(16'h76D4,4);
TASK_PP(16'h76D5,4);
TASK_PP(16'h76D6,4);
TASK_PP(16'h76D7,4);
TASK_PP(16'h76D8,4);
TASK_PP(16'h76D9,4);
TASK_PP(16'h76DA,4);
TASK_PP(16'h76DB,4);
TASK_PP(16'h76DC,4);
TASK_PP(16'h76DD,4);
TASK_PP(16'h76DE,4);
TASK_PP(16'h76DF,4);
TASK_PP(16'h76E0,4);
TASK_PP(16'h76E1,4);
TASK_PP(16'h76E2,4);
TASK_PP(16'h76E3,4);
TASK_PP(16'h76E4,4);
TASK_PP(16'h76E5,4);
TASK_PP(16'h76E6,4);
TASK_PP(16'h76E7,4);
TASK_PP(16'h76E8,4);
TASK_PP(16'h76E9,4);
TASK_PP(16'h76EA,4);
TASK_PP(16'h76EB,4);
TASK_PP(16'h76EC,4);
TASK_PP(16'h76ED,4);
TASK_PP(16'h76EE,4);
TASK_PP(16'h76EF,4);
TASK_PP(16'h76F0,4);
TASK_PP(16'h76F1,4);
TASK_PP(16'h76F2,4);
TASK_PP(16'h76F3,4);
TASK_PP(16'h76F4,4);
TASK_PP(16'h76F5,4);
TASK_PP(16'h76F6,4);
TASK_PP(16'h76F7,4);
TASK_PP(16'h76F8,4);
TASK_PP(16'h76F9,4);
TASK_PP(16'h76FA,4);
TASK_PP(16'h76FB,4);
TASK_PP(16'h76FC,4);
TASK_PP(16'h76FD,4);
TASK_PP(16'h76FE,4);
TASK_PP(16'h76FF,4);
TASK_PP(16'h7700,4);
TASK_PP(16'h7701,4);
TASK_PP(16'h7702,4);
TASK_PP(16'h7703,4);
TASK_PP(16'h7704,4);
TASK_PP(16'h7705,4);
TASK_PP(16'h7706,4);
TASK_PP(16'h7707,4);
TASK_PP(16'h7708,4);
TASK_PP(16'h7709,4);
TASK_PP(16'h770A,4);
TASK_PP(16'h770B,4);
TASK_PP(16'h770C,4);
TASK_PP(16'h770D,4);
TASK_PP(16'h770E,4);
TASK_PP(16'h770F,4);
TASK_PP(16'h7710,4);
TASK_PP(16'h7711,4);
TASK_PP(16'h7712,4);
TASK_PP(16'h7713,4);
TASK_PP(16'h7714,4);
TASK_PP(16'h7715,4);
TASK_PP(16'h7716,4);
TASK_PP(16'h7717,4);
TASK_PP(16'h7718,4);
TASK_PP(16'h7719,4);
TASK_PP(16'h771A,4);
TASK_PP(16'h771B,4);
TASK_PP(16'h771C,4);
TASK_PP(16'h771D,4);
TASK_PP(16'h771E,4);
TASK_PP(16'h771F,4);
TASK_PP(16'h7720,4);
TASK_PP(16'h7721,4);
TASK_PP(16'h7722,4);
TASK_PP(16'h7723,4);
TASK_PP(16'h7724,4);
TASK_PP(16'h7725,4);
TASK_PP(16'h7726,4);
TASK_PP(16'h7727,4);
TASK_PP(16'h7728,4);
TASK_PP(16'h7729,4);
TASK_PP(16'h772A,4);
TASK_PP(16'h772B,4);
TASK_PP(16'h772C,4);
TASK_PP(16'h772D,4);
TASK_PP(16'h772E,4);
TASK_PP(16'h772F,4);
TASK_PP(16'h7730,4);
TASK_PP(16'h7731,4);
TASK_PP(16'h7732,4);
TASK_PP(16'h7733,4);
TASK_PP(16'h7734,4);
TASK_PP(16'h7735,4);
TASK_PP(16'h7736,4);
TASK_PP(16'h7737,4);
TASK_PP(16'h7738,4);
TASK_PP(16'h7739,4);
TASK_PP(16'h773A,4);
TASK_PP(16'h773B,4);
TASK_PP(16'h773C,4);
TASK_PP(16'h773D,4);
TASK_PP(16'h773E,4);
TASK_PP(16'h773F,4);
TASK_PP(16'h7740,4);
TASK_PP(16'h7741,4);
TASK_PP(16'h7742,4);
TASK_PP(16'h7743,4);
TASK_PP(16'h7744,4);
TASK_PP(16'h7745,4);
TASK_PP(16'h7746,4);
TASK_PP(16'h7747,4);
TASK_PP(16'h7748,4);
TASK_PP(16'h7749,4);
TASK_PP(16'h774A,4);
TASK_PP(16'h774B,4);
TASK_PP(16'h774C,4);
TASK_PP(16'h774D,4);
TASK_PP(16'h774E,4);
TASK_PP(16'h774F,4);
TASK_PP(16'h7750,4);
TASK_PP(16'h7751,4);
TASK_PP(16'h7752,4);
TASK_PP(16'h7753,4);
TASK_PP(16'h7754,4);
TASK_PP(16'h7755,4);
TASK_PP(16'h7756,4);
TASK_PP(16'h7757,4);
TASK_PP(16'h7758,4);
TASK_PP(16'h7759,4);
TASK_PP(16'h775A,4);
TASK_PP(16'h775B,4);
TASK_PP(16'h775C,4);
TASK_PP(16'h775D,4);
TASK_PP(16'h775E,4);
TASK_PP(16'h775F,4);
TASK_PP(16'h7760,4);
TASK_PP(16'h7761,4);
TASK_PP(16'h7762,4);
TASK_PP(16'h7763,4);
TASK_PP(16'h7764,4);
TASK_PP(16'h7765,4);
TASK_PP(16'h7766,4);
TASK_PP(16'h7767,4);
TASK_PP(16'h7768,4);
TASK_PP(16'h7769,4);
TASK_PP(16'h776A,4);
TASK_PP(16'h776B,4);
TASK_PP(16'h776C,4);
TASK_PP(16'h776D,4);
TASK_PP(16'h776E,4);
TASK_PP(16'h776F,4);
TASK_PP(16'h7770,4);
TASK_PP(16'h7771,4);
TASK_PP(16'h7772,4);
TASK_PP(16'h7773,4);
TASK_PP(16'h7774,4);
TASK_PP(16'h7775,4);
TASK_PP(16'h7776,4);
TASK_PP(16'h7777,4);
TASK_PP(16'h7778,4);
TASK_PP(16'h7779,4);
TASK_PP(16'h777A,4);
TASK_PP(16'h777B,4);
TASK_PP(16'h777C,4);
TASK_PP(16'h777D,4);
TASK_PP(16'h777E,4);
TASK_PP(16'h777F,4);
TASK_PP(16'h7780,4);
TASK_PP(16'h7781,4);
TASK_PP(16'h7782,4);
TASK_PP(16'h7783,4);
TASK_PP(16'h7784,4);
TASK_PP(16'h7785,4);
TASK_PP(16'h7786,4);
TASK_PP(16'h7787,4);
TASK_PP(16'h7788,4);
TASK_PP(16'h7789,4);
TASK_PP(16'h778A,4);
TASK_PP(16'h778B,4);
TASK_PP(16'h778C,4);
TASK_PP(16'h778D,4);
TASK_PP(16'h778E,4);
TASK_PP(16'h778F,4);
TASK_PP(16'h7790,4);
TASK_PP(16'h7791,4);
TASK_PP(16'h7792,4);
TASK_PP(16'h7793,4);
TASK_PP(16'h7794,4);
TASK_PP(16'h7795,4);
TASK_PP(16'h7796,4);
TASK_PP(16'h7797,4);
TASK_PP(16'h7798,4);
TASK_PP(16'h7799,4);
TASK_PP(16'h779A,4);
TASK_PP(16'h779B,4);
TASK_PP(16'h779C,4);
TASK_PP(16'h779D,4);
TASK_PP(16'h779E,4);
TASK_PP(16'h779F,4);
TASK_PP(16'h77A0,4);
TASK_PP(16'h77A1,4);
TASK_PP(16'h77A2,4);
TASK_PP(16'h77A3,4);
TASK_PP(16'h77A4,4);
TASK_PP(16'h77A5,4);
TASK_PP(16'h77A6,4);
TASK_PP(16'h77A7,4);
TASK_PP(16'h77A8,4);
TASK_PP(16'h77A9,4);
TASK_PP(16'h77AA,4);
TASK_PP(16'h77AB,4);
TASK_PP(16'h77AC,4);
TASK_PP(16'h77AD,4);
TASK_PP(16'h77AE,4);
TASK_PP(16'h77AF,4);
TASK_PP(16'h77B0,4);
TASK_PP(16'h77B1,4);
TASK_PP(16'h77B2,4);
TASK_PP(16'h77B3,4);
TASK_PP(16'h77B4,4);
TASK_PP(16'h77B5,4);
TASK_PP(16'h77B6,4);
TASK_PP(16'h77B7,4);
TASK_PP(16'h77B8,4);
TASK_PP(16'h77B9,4);
TASK_PP(16'h77BA,4);
TASK_PP(16'h77BB,4);
TASK_PP(16'h77BC,4);
TASK_PP(16'h77BD,4);
TASK_PP(16'h77BE,4);
TASK_PP(16'h77BF,4);
TASK_PP(16'h77C0,4);
TASK_PP(16'h77C1,4);
TASK_PP(16'h77C2,4);
TASK_PP(16'h77C3,4);
TASK_PP(16'h77C4,4);
TASK_PP(16'h77C5,4);
TASK_PP(16'h77C6,4);
TASK_PP(16'h77C7,4);
TASK_PP(16'h77C8,4);
TASK_PP(16'h77C9,4);
TASK_PP(16'h77CA,4);
TASK_PP(16'h77CB,4);
TASK_PP(16'h77CC,4);
TASK_PP(16'h77CD,4);
TASK_PP(16'h77CE,4);
TASK_PP(16'h77CF,4);
TASK_PP(16'h77D0,4);
TASK_PP(16'h77D1,4);
TASK_PP(16'h77D2,4);
TASK_PP(16'h77D3,4);
TASK_PP(16'h77D4,4);
TASK_PP(16'h77D5,4);
TASK_PP(16'h77D6,4);
TASK_PP(16'h77D7,4);
TASK_PP(16'h77D8,4);
TASK_PP(16'h77D9,4);
TASK_PP(16'h77DA,4);
TASK_PP(16'h77DB,4);
TASK_PP(16'h77DC,4);
TASK_PP(16'h77DD,4);
TASK_PP(16'h77DE,4);
TASK_PP(16'h77DF,4);
TASK_PP(16'h77E0,4);
TASK_PP(16'h77E1,4);
TASK_PP(16'h77E2,4);
TASK_PP(16'h77E3,4);
TASK_PP(16'h77E4,4);
TASK_PP(16'h77E5,4);
TASK_PP(16'h77E6,4);
TASK_PP(16'h77E7,4);
TASK_PP(16'h77E8,4);
TASK_PP(16'h77E9,4);
TASK_PP(16'h77EA,4);
TASK_PP(16'h77EB,4);
TASK_PP(16'h77EC,4);
TASK_PP(16'h77ED,4);
TASK_PP(16'h77EE,4);
TASK_PP(16'h77EF,4);
TASK_PP(16'h77F0,4);
TASK_PP(16'h77F1,4);
TASK_PP(16'h77F2,4);
TASK_PP(16'h77F3,4);
TASK_PP(16'h77F4,4);
TASK_PP(16'h77F5,4);
TASK_PP(16'h77F6,4);
TASK_PP(16'h77F7,4);
TASK_PP(16'h77F8,4);
TASK_PP(16'h77F9,4);
TASK_PP(16'h77FA,4);
TASK_PP(16'h77FB,4);
TASK_PP(16'h77FC,4);
TASK_PP(16'h77FD,4);
TASK_PP(16'h77FE,4);
TASK_PP(16'h77FF,4);
TASK_PP(16'h7800,4);
TASK_PP(16'h7801,4);
TASK_PP(16'h7802,4);
TASK_PP(16'h7803,4);
TASK_PP(16'h7804,4);
TASK_PP(16'h7805,4);
TASK_PP(16'h7806,4);
TASK_PP(16'h7807,4);
TASK_PP(16'h7808,4);
TASK_PP(16'h7809,4);
TASK_PP(16'h780A,4);
TASK_PP(16'h780B,4);
TASK_PP(16'h780C,4);
TASK_PP(16'h780D,4);
TASK_PP(16'h780E,4);
TASK_PP(16'h780F,4);
TASK_PP(16'h7810,4);
TASK_PP(16'h7811,4);
TASK_PP(16'h7812,4);
TASK_PP(16'h7813,4);
TASK_PP(16'h7814,4);
TASK_PP(16'h7815,4);
TASK_PP(16'h7816,4);
TASK_PP(16'h7817,4);
TASK_PP(16'h7818,4);
TASK_PP(16'h7819,4);
TASK_PP(16'h781A,4);
TASK_PP(16'h781B,4);
TASK_PP(16'h781C,4);
TASK_PP(16'h781D,4);
TASK_PP(16'h781E,4);
TASK_PP(16'h781F,4);
TASK_PP(16'h7820,4);
TASK_PP(16'h7821,4);
TASK_PP(16'h7822,4);
TASK_PP(16'h7823,4);
TASK_PP(16'h7824,4);
TASK_PP(16'h7825,4);
TASK_PP(16'h7826,4);
TASK_PP(16'h7827,4);
TASK_PP(16'h7828,4);
TASK_PP(16'h7829,4);
TASK_PP(16'h782A,4);
TASK_PP(16'h782B,4);
TASK_PP(16'h782C,4);
TASK_PP(16'h782D,4);
TASK_PP(16'h782E,4);
TASK_PP(16'h782F,4);
TASK_PP(16'h7830,4);
TASK_PP(16'h7831,4);
TASK_PP(16'h7832,4);
TASK_PP(16'h7833,4);
TASK_PP(16'h7834,4);
TASK_PP(16'h7835,4);
TASK_PP(16'h7836,4);
TASK_PP(16'h7837,4);
TASK_PP(16'h7838,4);
TASK_PP(16'h7839,4);
TASK_PP(16'h783A,4);
TASK_PP(16'h783B,4);
TASK_PP(16'h783C,4);
TASK_PP(16'h783D,4);
TASK_PP(16'h783E,4);
TASK_PP(16'h783F,4);
TASK_PP(16'h7840,4);
TASK_PP(16'h7841,4);
TASK_PP(16'h7842,4);
TASK_PP(16'h7843,4);
TASK_PP(16'h7844,4);
TASK_PP(16'h7845,4);
TASK_PP(16'h7846,4);
TASK_PP(16'h7847,4);
TASK_PP(16'h7848,4);
TASK_PP(16'h7849,4);
TASK_PP(16'h784A,4);
TASK_PP(16'h784B,4);
TASK_PP(16'h784C,4);
TASK_PP(16'h784D,4);
TASK_PP(16'h784E,4);
TASK_PP(16'h784F,4);
TASK_PP(16'h7850,4);
TASK_PP(16'h7851,4);
TASK_PP(16'h7852,4);
TASK_PP(16'h7853,4);
TASK_PP(16'h7854,4);
TASK_PP(16'h7855,4);
TASK_PP(16'h7856,4);
TASK_PP(16'h7857,4);
TASK_PP(16'h7858,4);
TASK_PP(16'h7859,4);
TASK_PP(16'h785A,4);
TASK_PP(16'h785B,4);
TASK_PP(16'h785C,4);
TASK_PP(16'h785D,4);
TASK_PP(16'h785E,4);
TASK_PP(16'h785F,4);
TASK_PP(16'h7860,4);
TASK_PP(16'h7861,4);
TASK_PP(16'h7862,4);
TASK_PP(16'h7863,4);
TASK_PP(16'h7864,4);
TASK_PP(16'h7865,4);
TASK_PP(16'h7866,4);
TASK_PP(16'h7867,4);
TASK_PP(16'h7868,4);
TASK_PP(16'h7869,4);
TASK_PP(16'h786A,4);
TASK_PP(16'h786B,4);
TASK_PP(16'h786C,4);
TASK_PP(16'h786D,4);
TASK_PP(16'h786E,4);
TASK_PP(16'h786F,4);
TASK_PP(16'h7870,4);
TASK_PP(16'h7871,4);
TASK_PP(16'h7872,4);
TASK_PP(16'h7873,4);
TASK_PP(16'h7874,4);
TASK_PP(16'h7875,4);
TASK_PP(16'h7876,4);
TASK_PP(16'h7877,4);
TASK_PP(16'h7878,4);
TASK_PP(16'h7879,4);
TASK_PP(16'h787A,4);
TASK_PP(16'h787B,4);
TASK_PP(16'h787C,4);
TASK_PP(16'h787D,4);
TASK_PP(16'h787E,4);
TASK_PP(16'h787F,4);
TASK_PP(16'h7880,4);
TASK_PP(16'h7881,4);
TASK_PP(16'h7882,4);
TASK_PP(16'h7883,4);
TASK_PP(16'h7884,4);
TASK_PP(16'h7885,4);
TASK_PP(16'h7886,4);
TASK_PP(16'h7887,4);
TASK_PP(16'h7888,4);
TASK_PP(16'h7889,4);
TASK_PP(16'h788A,4);
TASK_PP(16'h788B,4);
TASK_PP(16'h788C,4);
TASK_PP(16'h788D,4);
TASK_PP(16'h788E,4);
TASK_PP(16'h788F,4);
TASK_PP(16'h7890,4);
TASK_PP(16'h7891,4);
TASK_PP(16'h7892,4);
TASK_PP(16'h7893,4);
TASK_PP(16'h7894,4);
TASK_PP(16'h7895,4);
TASK_PP(16'h7896,4);
TASK_PP(16'h7897,4);
TASK_PP(16'h7898,4);
TASK_PP(16'h7899,4);
TASK_PP(16'h789A,4);
TASK_PP(16'h789B,4);
TASK_PP(16'h789C,4);
TASK_PP(16'h789D,4);
TASK_PP(16'h789E,4);
TASK_PP(16'h789F,4);
TASK_PP(16'h78A0,4);
TASK_PP(16'h78A1,4);
TASK_PP(16'h78A2,4);
TASK_PP(16'h78A3,4);
TASK_PP(16'h78A4,4);
TASK_PP(16'h78A5,4);
TASK_PP(16'h78A6,4);
TASK_PP(16'h78A7,4);
TASK_PP(16'h78A8,4);
TASK_PP(16'h78A9,4);
TASK_PP(16'h78AA,4);
TASK_PP(16'h78AB,4);
TASK_PP(16'h78AC,4);
TASK_PP(16'h78AD,4);
TASK_PP(16'h78AE,4);
TASK_PP(16'h78AF,4);
TASK_PP(16'h78B0,4);
TASK_PP(16'h78B1,4);
TASK_PP(16'h78B2,4);
TASK_PP(16'h78B3,4);
TASK_PP(16'h78B4,4);
TASK_PP(16'h78B5,4);
TASK_PP(16'h78B6,4);
TASK_PP(16'h78B7,4);
TASK_PP(16'h78B8,4);
TASK_PP(16'h78B9,4);
TASK_PP(16'h78BA,4);
TASK_PP(16'h78BB,4);
TASK_PP(16'h78BC,4);
TASK_PP(16'h78BD,4);
TASK_PP(16'h78BE,4);
TASK_PP(16'h78BF,4);
TASK_PP(16'h78C0,4);
TASK_PP(16'h78C1,4);
TASK_PP(16'h78C2,4);
TASK_PP(16'h78C3,4);
TASK_PP(16'h78C4,4);
TASK_PP(16'h78C5,4);
TASK_PP(16'h78C6,4);
TASK_PP(16'h78C7,4);
TASK_PP(16'h78C8,4);
TASK_PP(16'h78C9,4);
TASK_PP(16'h78CA,4);
TASK_PP(16'h78CB,4);
TASK_PP(16'h78CC,4);
TASK_PP(16'h78CD,4);
TASK_PP(16'h78CE,4);
TASK_PP(16'h78CF,4);
TASK_PP(16'h78D0,4);
TASK_PP(16'h78D1,4);
TASK_PP(16'h78D2,4);
TASK_PP(16'h78D3,4);
TASK_PP(16'h78D4,4);
TASK_PP(16'h78D5,4);
TASK_PP(16'h78D6,4);
TASK_PP(16'h78D7,4);
TASK_PP(16'h78D8,4);
TASK_PP(16'h78D9,4);
TASK_PP(16'h78DA,4);
TASK_PP(16'h78DB,4);
TASK_PP(16'h78DC,4);
TASK_PP(16'h78DD,4);
TASK_PP(16'h78DE,4);
TASK_PP(16'h78DF,4);
TASK_PP(16'h78E0,4);
TASK_PP(16'h78E1,4);
TASK_PP(16'h78E2,4);
TASK_PP(16'h78E3,4);
TASK_PP(16'h78E4,4);
TASK_PP(16'h78E5,4);
TASK_PP(16'h78E6,4);
TASK_PP(16'h78E7,4);
TASK_PP(16'h78E8,4);
TASK_PP(16'h78E9,4);
TASK_PP(16'h78EA,4);
TASK_PP(16'h78EB,4);
TASK_PP(16'h78EC,4);
TASK_PP(16'h78ED,4);
TASK_PP(16'h78EE,4);
TASK_PP(16'h78EF,4);
TASK_PP(16'h78F0,4);
TASK_PP(16'h78F1,4);
TASK_PP(16'h78F2,4);
TASK_PP(16'h78F3,4);
TASK_PP(16'h78F4,4);
TASK_PP(16'h78F5,4);
TASK_PP(16'h78F6,4);
TASK_PP(16'h78F7,4);
TASK_PP(16'h78F8,4);
TASK_PP(16'h78F9,4);
TASK_PP(16'h78FA,4);
TASK_PP(16'h78FB,4);
TASK_PP(16'h78FC,4);
TASK_PP(16'h78FD,4);
TASK_PP(16'h78FE,4);
TASK_PP(16'h78FF,4);
TASK_PP(16'h7900,4);
TASK_PP(16'h7901,4);
TASK_PP(16'h7902,4);
TASK_PP(16'h7903,4);
TASK_PP(16'h7904,4);
TASK_PP(16'h7905,4);
TASK_PP(16'h7906,4);
TASK_PP(16'h7907,4);
TASK_PP(16'h7908,4);
TASK_PP(16'h7909,4);
TASK_PP(16'h790A,4);
TASK_PP(16'h790B,4);
TASK_PP(16'h790C,4);
TASK_PP(16'h790D,4);
TASK_PP(16'h790E,4);
TASK_PP(16'h790F,4);
TASK_PP(16'h7910,4);
TASK_PP(16'h7911,4);
TASK_PP(16'h7912,4);
TASK_PP(16'h7913,4);
TASK_PP(16'h7914,4);
TASK_PP(16'h7915,4);
TASK_PP(16'h7916,4);
TASK_PP(16'h7917,4);
TASK_PP(16'h7918,4);
TASK_PP(16'h7919,4);
TASK_PP(16'h791A,4);
TASK_PP(16'h791B,4);
TASK_PP(16'h791C,4);
TASK_PP(16'h791D,4);
TASK_PP(16'h791E,4);
TASK_PP(16'h791F,4);
TASK_PP(16'h7920,4);
TASK_PP(16'h7921,4);
TASK_PP(16'h7922,4);
TASK_PP(16'h7923,4);
TASK_PP(16'h7924,4);
TASK_PP(16'h7925,4);
TASK_PP(16'h7926,4);
TASK_PP(16'h7927,4);
TASK_PP(16'h7928,4);
TASK_PP(16'h7929,4);
TASK_PP(16'h792A,4);
TASK_PP(16'h792B,4);
TASK_PP(16'h792C,4);
TASK_PP(16'h792D,4);
TASK_PP(16'h792E,4);
TASK_PP(16'h792F,4);
TASK_PP(16'h7930,4);
TASK_PP(16'h7931,4);
TASK_PP(16'h7932,4);
TASK_PP(16'h7933,4);
TASK_PP(16'h7934,4);
TASK_PP(16'h7935,4);
TASK_PP(16'h7936,4);
TASK_PP(16'h7937,4);
TASK_PP(16'h7938,4);
TASK_PP(16'h7939,4);
TASK_PP(16'h793A,4);
TASK_PP(16'h793B,4);
TASK_PP(16'h793C,4);
TASK_PP(16'h793D,4);
TASK_PP(16'h793E,4);
TASK_PP(16'h793F,4);
TASK_PP(16'h7940,4);
TASK_PP(16'h7941,4);
TASK_PP(16'h7942,4);
TASK_PP(16'h7943,4);
TASK_PP(16'h7944,4);
TASK_PP(16'h7945,4);
TASK_PP(16'h7946,4);
TASK_PP(16'h7947,4);
TASK_PP(16'h7948,4);
TASK_PP(16'h7949,4);
TASK_PP(16'h794A,4);
TASK_PP(16'h794B,4);
TASK_PP(16'h794C,4);
TASK_PP(16'h794D,4);
TASK_PP(16'h794E,4);
TASK_PP(16'h794F,4);
TASK_PP(16'h7950,4);
TASK_PP(16'h7951,4);
TASK_PP(16'h7952,4);
TASK_PP(16'h7953,4);
TASK_PP(16'h7954,4);
TASK_PP(16'h7955,4);
TASK_PP(16'h7956,4);
TASK_PP(16'h7957,4);
TASK_PP(16'h7958,4);
TASK_PP(16'h7959,4);
TASK_PP(16'h795A,4);
TASK_PP(16'h795B,4);
TASK_PP(16'h795C,4);
TASK_PP(16'h795D,4);
TASK_PP(16'h795E,4);
TASK_PP(16'h795F,4);
TASK_PP(16'h7960,4);
TASK_PP(16'h7961,4);
TASK_PP(16'h7962,4);
TASK_PP(16'h7963,4);
TASK_PP(16'h7964,4);
TASK_PP(16'h7965,4);
TASK_PP(16'h7966,4);
TASK_PP(16'h7967,4);
TASK_PP(16'h7968,4);
TASK_PP(16'h7969,4);
TASK_PP(16'h796A,4);
TASK_PP(16'h796B,4);
TASK_PP(16'h796C,4);
TASK_PP(16'h796D,4);
TASK_PP(16'h796E,4);
TASK_PP(16'h796F,4);
TASK_PP(16'h7970,4);
TASK_PP(16'h7971,4);
TASK_PP(16'h7972,4);
TASK_PP(16'h7973,4);
TASK_PP(16'h7974,4);
TASK_PP(16'h7975,4);
TASK_PP(16'h7976,4);
TASK_PP(16'h7977,4);
TASK_PP(16'h7978,4);
TASK_PP(16'h7979,4);
TASK_PP(16'h797A,4);
TASK_PP(16'h797B,4);
TASK_PP(16'h797C,4);
TASK_PP(16'h797D,4);
TASK_PP(16'h797E,4);
TASK_PP(16'h797F,4);
TASK_PP(16'h7980,4);
TASK_PP(16'h7981,4);
TASK_PP(16'h7982,4);
TASK_PP(16'h7983,4);
TASK_PP(16'h7984,4);
TASK_PP(16'h7985,4);
TASK_PP(16'h7986,4);
TASK_PP(16'h7987,4);
TASK_PP(16'h7988,4);
TASK_PP(16'h7989,4);
TASK_PP(16'h798A,4);
TASK_PP(16'h798B,4);
TASK_PP(16'h798C,4);
TASK_PP(16'h798D,4);
TASK_PP(16'h798E,4);
TASK_PP(16'h798F,4);
TASK_PP(16'h7990,4);
TASK_PP(16'h7991,4);
TASK_PP(16'h7992,4);
TASK_PP(16'h7993,4);
TASK_PP(16'h7994,4);
TASK_PP(16'h7995,4);
TASK_PP(16'h7996,4);
TASK_PP(16'h7997,4);
TASK_PP(16'h7998,4);
TASK_PP(16'h7999,4);
TASK_PP(16'h799A,4);
TASK_PP(16'h799B,4);
TASK_PP(16'h799C,4);
TASK_PP(16'h799D,4);
TASK_PP(16'h799E,4);
TASK_PP(16'h799F,4);
TASK_PP(16'h79A0,4);
TASK_PP(16'h79A1,4);
TASK_PP(16'h79A2,4);
TASK_PP(16'h79A3,4);
TASK_PP(16'h79A4,4);
TASK_PP(16'h79A5,4);
TASK_PP(16'h79A6,4);
TASK_PP(16'h79A7,4);
TASK_PP(16'h79A8,4);
TASK_PP(16'h79A9,4);
TASK_PP(16'h79AA,4);
TASK_PP(16'h79AB,4);
TASK_PP(16'h79AC,4);
TASK_PP(16'h79AD,4);
TASK_PP(16'h79AE,4);
TASK_PP(16'h79AF,4);
TASK_PP(16'h79B0,4);
TASK_PP(16'h79B1,4);
TASK_PP(16'h79B2,4);
TASK_PP(16'h79B3,4);
TASK_PP(16'h79B4,4);
TASK_PP(16'h79B5,4);
TASK_PP(16'h79B6,4);
TASK_PP(16'h79B7,4);
TASK_PP(16'h79B8,4);
TASK_PP(16'h79B9,4);
TASK_PP(16'h79BA,4);
TASK_PP(16'h79BB,4);
TASK_PP(16'h79BC,4);
TASK_PP(16'h79BD,4);
TASK_PP(16'h79BE,4);
TASK_PP(16'h79BF,4);
TASK_PP(16'h79C0,4);
TASK_PP(16'h79C1,4);
TASK_PP(16'h79C2,4);
TASK_PP(16'h79C3,4);
TASK_PP(16'h79C4,4);
TASK_PP(16'h79C5,4);
TASK_PP(16'h79C6,4);
TASK_PP(16'h79C7,4);
TASK_PP(16'h79C8,4);
TASK_PP(16'h79C9,4);
TASK_PP(16'h79CA,4);
TASK_PP(16'h79CB,4);
TASK_PP(16'h79CC,4);
TASK_PP(16'h79CD,4);
TASK_PP(16'h79CE,4);
TASK_PP(16'h79CF,4);
TASK_PP(16'h79D0,4);
TASK_PP(16'h79D1,4);
TASK_PP(16'h79D2,4);
TASK_PP(16'h79D3,4);
TASK_PP(16'h79D4,4);
TASK_PP(16'h79D5,4);
TASK_PP(16'h79D6,4);
TASK_PP(16'h79D7,4);
TASK_PP(16'h79D8,4);
TASK_PP(16'h79D9,4);
TASK_PP(16'h79DA,4);
TASK_PP(16'h79DB,4);
TASK_PP(16'h79DC,4);
TASK_PP(16'h79DD,4);
TASK_PP(16'h79DE,4);
TASK_PP(16'h79DF,4);
TASK_PP(16'h79E0,4);
TASK_PP(16'h79E1,4);
TASK_PP(16'h79E2,4);
TASK_PP(16'h79E3,4);
TASK_PP(16'h79E4,4);
TASK_PP(16'h79E5,4);
TASK_PP(16'h79E6,4);
TASK_PP(16'h79E7,4);
TASK_PP(16'h79E8,4);
TASK_PP(16'h79E9,4);
TASK_PP(16'h79EA,4);
TASK_PP(16'h79EB,4);
TASK_PP(16'h79EC,4);
TASK_PP(16'h79ED,4);
TASK_PP(16'h79EE,4);
TASK_PP(16'h79EF,4);
TASK_PP(16'h79F0,4);
TASK_PP(16'h79F1,4);
TASK_PP(16'h79F2,4);
TASK_PP(16'h79F3,4);
TASK_PP(16'h79F4,4);
TASK_PP(16'h79F5,4);
TASK_PP(16'h79F6,4);
TASK_PP(16'h79F7,4);
TASK_PP(16'h79F8,4);
TASK_PP(16'h79F9,4);
TASK_PP(16'h79FA,4);
TASK_PP(16'h79FB,4);
TASK_PP(16'h79FC,4);
TASK_PP(16'h79FD,4);
TASK_PP(16'h79FE,4);
TASK_PP(16'h79FF,4);
TASK_PP(16'h7A00,4);
TASK_PP(16'h7A01,4);
TASK_PP(16'h7A02,4);
TASK_PP(16'h7A03,4);
TASK_PP(16'h7A04,4);
TASK_PP(16'h7A05,4);
TASK_PP(16'h7A06,4);
TASK_PP(16'h7A07,4);
TASK_PP(16'h7A08,4);
TASK_PP(16'h7A09,4);
TASK_PP(16'h7A0A,4);
TASK_PP(16'h7A0B,4);
TASK_PP(16'h7A0C,4);
TASK_PP(16'h7A0D,4);
TASK_PP(16'h7A0E,4);
TASK_PP(16'h7A0F,4);
TASK_PP(16'h7A10,4);
TASK_PP(16'h7A11,4);
TASK_PP(16'h7A12,4);
TASK_PP(16'h7A13,4);
TASK_PP(16'h7A14,4);
TASK_PP(16'h7A15,4);
TASK_PP(16'h7A16,4);
TASK_PP(16'h7A17,4);
TASK_PP(16'h7A18,4);
TASK_PP(16'h7A19,4);
TASK_PP(16'h7A1A,4);
TASK_PP(16'h7A1B,4);
TASK_PP(16'h7A1C,4);
TASK_PP(16'h7A1D,4);
TASK_PP(16'h7A1E,4);
TASK_PP(16'h7A1F,4);
TASK_PP(16'h7A20,4);
TASK_PP(16'h7A21,4);
TASK_PP(16'h7A22,4);
TASK_PP(16'h7A23,4);
TASK_PP(16'h7A24,4);
TASK_PP(16'h7A25,4);
TASK_PP(16'h7A26,4);
TASK_PP(16'h7A27,4);
TASK_PP(16'h7A28,4);
TASK_PP(16'h7A29,4);
TASK_PP(16'h7A2A,4);
TASK_PP(16'h7A2B,4);
TASK_PP(16'h7A2C,4);
TASK_PP(16'h7A2D,4);
TASK_PP(16'h7A2E,4);
TASK_PP(16'h7A2F,4);
TASK_PP(16'h7A30,4);
TASK_PP(16'h7A31,4);
TASK_PP(16'h7A32,4);
TASK_PP(16'h7A33,4);
TASK_PP(16'h7A34,4);
TASK_PP(16'h7A35,4);
TASK_PP(16'h7A36,4);
TASK_PP(16'h7A37,4);
TASK_PP(16'h7A38,4);
TASK_PP(16'h7A39,4);
TASK_PP(16'h7A3A,4);
TASK_PP(16'h7A3B,4);
TASK_PP(16'h7A3C,4);
TASK_PP(16'h7A3D,4);
TASK_PP(16'h7A3E,4);
TASK_PP(16'h7A3F,4);
TASK_PP(16'h7A40,4);
TASK_PP(16'h7A41,4);
TASK_PP(16'h7A42,4);
TASK_PP(16'h7A43,4);
TASK_PP(16'h7A44,4);
TASK_PP(16'h7A45,4);
TASK_PP(16'h7A46,4);
TASK_PP(16'h7A47,4);
TASK_PP(16'h7A48,4);
TASK_PP(16'h7A49,4);
TASK_PP(16'h7A4A,4);
TASK_PP(16'h7A4B,4);
TASK_PP(16'h7A4C,4);
TASK_PP(16'h7A4D,4);
TASK_PP(16'h7A4E,4);
TASK_PP(16'h7A4F,4);
TASK_PP(16'h7A50,4);
TASK_PP(16'h7A51,4);
TASK_PP(16'h7A52,4);
TASK_PP(16'h7A53,4);
TASK_PP(16'h7A54,4);
TASK_PP(16'h7A55,4);
TASK_PP(16'h7A56,4);
TASK_PP(16'h7A57,4);
TASK_PP(16'h7A58,4);
TASK_PP(16'h7A59,4);
TASK_PP(16'h7A5A,4);
TASK_PP(16'h7A5B,4);
TASK_PP(16'h7A5C,4);
TASK_PP(16'h7A5D,4);
TASK_PP(16'h7A5E,4);
TASK_PP(16'h7A5F,4);
TASK_PP(16'h7A60,4);
TASK_PP(16'h7A61,4);
TASK_PP(16'h7A62,4);
TASK_PP(16'h7A63,4);
TASK_PP(16'h7A64,4);
TASK_PP(16'h7A65,4);
TASK_PP(16'h7A66,4);
TASK_PP(16'h7A67,4);
TASK_PP(16'h7A68,4);
TASK_PP(16'h7A69,4);
TASK_PP(16'h7A6A,4);
TASK_PP(16'h7A6B,4);
TASK_PP(16'h7A6C,4);
TASK_PP(16'h7A6D,4);
TASK_PP(16'h7A6E,4);
TASK_PP(16'h7A6F,4);
TASK_PP(16'h7A70,4);
TASK_PP(16'h7A71,4);
TASK_PP(16'h7A72,4);
TASK_PP(16'h7A73,4);
TASK_PP(16'h7A74,4);
TASK_PP(16'h7A75,4);
TASK_PP(16'h7A76,4);
TASK_PP(16'h7A77,4);
TASK_PP(16'h7A78,4);
TASK_PP(16'h7A79,4);
TASK_PP(16'h7A7A,4);
TASK_PP(16'h7A7B,4);
TASK_PP(16'h7A7C,4);
TASK_PP(16'h7A7D,4);
TASK_PP(16'h7A7E,4);
TASK_PP(16'h7A7F,4);
TASK_PP(16'h7A80,4);
TASK_PP(16'h7A81,4);
TASK_PP(16'h7A82,4);
TASK_PP(16'h7A83,4);
TASK_PP(16'h7A84,4);
TASK_PP(16'h7A85,4);
TASK_PP(16'h7A86,4);
TASK_PP(16'h7A87,4);
TASK_PP(16'h7A88,4);
TASK_PP(16'h7A89,4);
TASK_PP(16'h7A8A,4);
TASK_PP(16'h7A8B,4);
TASK_PP(16'h7A8C,4);
TASK_PP(16'h7A8D,4);
TASK_PP(16'h7A8E,4);
TASK_PP(16'h7A8F,4);
TASK_PP(16'h7A90,4);
TASK_PP(16'h7A91,4);
TASK_PP(16'h7A92,4);
TASK_PP(16'h7A93,4);
TASK_PP(16'h7A94,4);
TASK_PP(16'h7A95,4);
TASK_PP(16'h7A96,4);
TASK_PP(16'h7A97,4);
TASK_PP(16'h7A98,4);
TASK_PP(16'h7A99,4);
TASK_PP(16'h7A9A,4);
TASK_PP(16'h7A9B,4);
TASK_PP(16'h7A9C,4);
TASK_PP(16'h7A9D,4);
TASK_PP(16'h7A9E,4);
TASK_PP(16'h7A9F,4);
TASK_PP(16'h7AA0,4);
TASK_PP(16'h7AA1,4);
TASK_PP(16'h7AA2,4);
TASK_PP(16'h7AA3,4);
TASK_PP(16'h7AA4,4);
TASK_PP(16'h7AA5,4);
TASK_PP(16'h7AA6,4);
TASK_PP(16'h7AA7,4);
TASK_PP(16'h7AA8,4);
TASK_PP(16'h7AA9,4);
TASK_PP(16'h7AAA,4);
TASK_PP(16'h7AAB,4);
TASK_PP(16'h7AAC,4);
TASK_PP(16'h7AAD,4);
TASK_PP(16'h7AAE,4);
TASK_PP(16'h7AAF,4);
TASK_PP(16'h7AB0,4);
TASK_PP(16'h7AB1,4);
TASK_PP(16'h7AB2,4);
TASK_PP(16'h7AB3,4);
TASK_PP(16'h7AB4,4);
TASK_PP(16'h7AB5,4);
TASK_PP(16'h7AB6,4);
TASK_PP(16'h7AB7,4);
TASK_PP(16'h7AB8,4);
TASK_PP(16'h7AB9,4);
TASK_PP(16'h7ABA,4);
TASK_PP(16'h7ABB,4);
TASK_PP(16'h7ABC,4);
TASK_PP(16'h7ABD,4);
TASK_PP(16'h7ABE,4);
TASK_PP(16'h7ABF,4);
TASK_PP(16'h7AC0,4);
TASK_PP(16'h7AC1,4);
TASK_PP(16'h7AC2,4);
TASK_PP(16'h7AC3,4);
TASK_PP(16'h7AC4,4);
TASK_PP(16'h7AC5,4);
TASK_PP(16'h7AC6,4);
TASK_PP(16'h7AC7,4);
TASK_PP(16'h7AC8,4);
TASK_PP(16'h7AC9,4);
TASK_PP(16'h7ACA,4);
TASK_PP(16'h7ACB,4);
TASK_PP(16'h7ACC,4);
TASK_PP(16'h7ACD,4);
TASK_PP(16'h7ACE,4);
TASK_PP(16'h7ACF,4);
TASK_PP(16'h7AD0,4);
TASK_PP(16'h7AD1,4);
TASK_PP(16'h7AD2,4);
TASK_PP(16'h7AD3,4);
TASK_PP(16'h7AD4,4);
TASK_PP(16'h7AD5,4);
TASK_PP(16'h7AD6,4);
TASK_PP(16'h7AD7,4);
TASK_PP(16'h7AD8,4);
TASK_PP(16'h7AD9,4);
TASK_PP(16'h7ADA,4);
TASK_PP(16'h7ADB,4);
TASK_PP(16'h7ADC,4);
TASK_PP(16'h7ADD,4);
TASK_PP(16'h7ADE,4);
TASK_PP(16'h7ADF,4);
TASK_PP(16'h7AE0,4);
TASK_PP(16'h7AE1,4);
TASK_PP(16'h7AE2,4);
TASK_PP(16'h7AE3,4);
TASK_PP(16'h7AE4,4);
TASK_PP(16'h7AE5,4);
TASK_PP(16'h7AE6,4);
TASK_PP(16'h7AE7,4);
TASK_PP(16'h7AE8,4);
TASK_PP(16'h7AE9,4);
TASK_PP(16'h7AEA,4);
TASK_PP(16'h7AEB,4);
TASK_PP(16'h7AEC,4);
TASK_PP(16'h7AED,4);
TASK_PP(16'h7AEE,4);
TASK_PP(16'h7AEF,4);
TASK_PP(16'h7AF0,4);
TASK_PP(16'h7AF1,4);
TASK_PP(16'h7AF2,4);
TASK_PP(16'h7AF3,4);
TASK_PP(16'h7AF4,4);
TASK_PP(16'h7AF5,4);
TASK_PP(16'h7AF6,4);
TASK_PP(16'h7AF7,4);
TASK_PP(16'h7AF8,4);
TASK_PP(16'h7AF9,4);
TASK_PP(16'h7AFA,4);
TASK_PP(16'h7AFB,4);
TASK_PP(16'h7AFC,4);
TASK_PP(16'h7AFD,4);
TASK_PP(16'h7AFE,4);
TASK_PP(16'h7AFF,4);
TASK_PP(16'h7B00,4);
TASK_PP(16'h7B01,4);
TASK_PP(16'h7B02,4);
TASK_PP(16'h7B03,4);
TASK_PP(16'h7B04,4);
TASK_PP(16'h7B05,4);
TASK_PP(16'h7B06,4);
TASK_PP(16'h7B07,4);
TASK_PP(16'h7B08,4);
TASK_PP(16'h7B09,4);
TASK_PP(16'h7B0A,4);
TASK_PP(16'h7B0B,4);
TASK_PP(16'h7B0C,4);
TASK_PP(16'h7B0D,4);
TASK_PP(16'h7B0E,4);
TASK_PP(16'h7B0F,4);
TASK_PP(16'h7B10,4);
TASK_PP(16'h7B11,4);
TASK_PP(16'h7B12,4);
TASK_PP(16'h7B13,4);
TASK_PP(16'h7B14,4);
TASK_PP(16'h7B15,4);
TASK_PP(16'h7B16,4);
TASK_PP(16'h7B17,4);
TASK_PP(16'h7B18,4);
TASK_PP(16'h7B19,4);
TASK_PP(16'h7B1A,4);
TASK_PP(16'h7B1B,4);
TASK_PP(16'h7B1C,4);
TASK_PP(16'h7B1D,4);
TASK_PP(16'h7B1E,4);
TASK_PP(16'h7B1F,4);
TASK_PP(16'h7B20,4);
TASK_PP(16'h7B21,4);
TASK_PP(16'h7B22,4);
TASK_PP(16'h7B23,4);
TASK_PP(16'h7B24,4);
TASK_PP(16'h7B25,4);
TASK_PP(16'h7B26,4);
TASK_PP(16'h7B27,4);
TASK_PP(16'h7B28,4);
TASK_PP(16'h7B29,4);
TASK_PP(16'h7B2A,4);
TASK_PP(16'h7B2B,4);
TASK_PP(16'h7B2C,4);
TASK_PP(16'h7B2D,4);
TASK_PP(16'h7B2E,4);
TASK_PP(16'h7B2F,4);
TASK_PP(16'h7B30,4);
TASK_PP(16'h7B31,4);
TASK_PP(16'h7B32,4);
TASK_PP(16'h7B33,4);
TASK_PP(16'h7B34,4);
TASK_PP(16'h7B35,4);
TASK_PP(16'h7B36,4);
TASK_PP(16'h7B37,4);
TASK_PP(16'h7B38,4);
TASK_PP(16'h7B39,4);
TASK_PP(16'h7B3A,4);
TASK_PP(16'h7B3B,4);
TASK_PP(16'h7B3C,4);
TASK_PP(16'h7B3D,4);
TASK_PP(16'h7B3E,4);
TASK_PP(16'h7B3F,4);
TASK_PP(16'h7B40,4);
TASK_PP(16'h7B41,4);
TASK_PP(16'h7B42,4);
TASK_PP(16'h7B43,4);
TASK_PP(16'h7B44,4);
TASK_PP(16'h7B45,4);
TASK_PP(16'h7B46,4);
TASK_PP(16'h7B47,4);
TASK_PP(16'h7B48,4);
TASK_PP(16'h7B49,4);
TASK_PP(16'h7B4A,4);
TASK_PP(16'h7B4B,4);
TASK_PP(16'h7B4C,4);
TASK_PP(16'h7B4D,4);
TASK_PP(16'h7B4E,4);
TASK_PP(16'h7B4F,4);
TASK_PP(16'h7B50,4);
TASK_PP(16'h7B51,4);
TASK_PP(16'h7B52,4);
TASK_PP(16'h7B53,4);
TASK_PP(16'h7B54,4);
TASK_PP(16'h7B55,4);
TASK_PP(16'h7B56,4);
TASK_PP(16'h7B57,4);
TASK_PP(16'h7B58,4);
TASK_PP(16'h7B59,4);
TASK_PP(16'h7B5A,4);
TASK_PP(16'h7B5B,4);
TASK_PP(16'h7B5C,4);
TASK_PP(16'h7B5D,4);
TASK_PP(16'h7B5E,4);
TASK_PP(16'h7B5F,4);
TASK_PP(16'h7B60,4);
TASK_PP(16'h7B61,4);
TASK_PP(16'h7B62,4);
TASK_PP(16'h7B63,4);
TASK_PP(16'h7B64,4);
TASK_PP(16'h7B65,4);
TASK_PP(16'h7B66,4);
TASK_PP(16'h7B67,4);
TASK_PP(16'h7B68,4);
TASK_PP(16'h7B69,4);
TASK_PP(16'h7B6A,4);
TASK_PP(16'h7B6B,4);
TASK_PP(16'h7B6C,4);
TASK_PP(16'h7B6D,4);
TASK_PP(16'h7B6E,4);
TASK_PP(16'h7B6F,4);
TASK_PP(16'h7B70,4);
TASK_PP(16'h7B71,4);
TASK_PP(16'h7B72,4);
TASK_PP(16'h7B73,4);
TASK_PP(16'h7B74,4);
TASK_PP(16'h7B75,4);
TASK_PP(16'h7B76,4);
TASK_PP(16'h7B77,4);
TASK_PP(16'h7B78,4);
TASK_PP(16'h7B79,4);
TASK_PP(16'h7B7A,4);
TASK_PP(16'h7B7B,4);
TASK_PP(16'h7B7C,4);
TASK_PP(16'h7B7D,4);
TASK_PP(16'h7B7E,4);
TASK_PP(16'h7B7F,4);
TASK_PP(16'h7B80,4);
TASK_PP(16'h7B81,4);
TASK_PP(16'h7B82,4);
TASK_PP(16'h7B83,4);
TASK_PP(16'h7B84,4);
TASK_PP(16'h7B85,4);
TASK_PP(16'h7B86,4);
TASK_PP(16'h7B87,4);
TASK_PP(16'h7B88,4);
TASK_PP(16'h7B89,4);
TASK_PP(16'h7B8A,4);
TASK_PP(16'h7B8B,4);
TASK_PP(16'h7B8C,4);
TASK_PP(16'h7B8D,4);
TASK_PP(16'h7B8E,4);
TASK_PP(16'h7B8F,4);
TASK_PP(16'h7B90,4);
TASK_PP(16'h7B91,4);
TASK_PP(16'h7B92,4);
TASK_PP(16'h7B93,4);
TASK_PP(16'h7B94,4);
TASK_PP(16'h7B95,4);
TASK_PP(16'h7B96,4);
TASK_PP(16'h7B97,4);
TASK_PP(16'h7B98,4);
TASK_PP(16'h7B99,4);
TASK_PP(16'h7B9A,4);
TASK_PP(16'h7B9B,4);
TASK_PP(16'h7B9C,4);
TASK_PP(16'h7B9D,4);
TASK_PP(16'h7B9E,4);
TASK_PP(16'h7B9F,4);
TASK_PP(16'h7BA0,4);
TASK_PP(16'h7BA1,4);
TASK_PP(16'h7BA2,4);
TASK_PP(16'h7BA3,4);
TASK_PP(16'h7BA4,4);
TASK_PP(16'h7BA5,4);
TASK_PP(16'h7BA6,4);
TASK_PP(16'h7BA7,4);
TASK_PP(16'h7BA8,4);
TASK_PP(16'h7BA9,4);
TASK_PP(16'h7BAA,4);
TASK_PP(16'h7BAB,4);
TASK_PP(16'h7BAC,4);
TASK_PP(16'h7BAD,4);
TASK_PP(16'h7BAE,4);
TASK_PP(16'h7BAF,4);
TASK_PP(16'h7BB0,4);
TASK_PP(16'h7BB1,4);
TASK_PP(16'h7BB2,4);
TASK_PP(16'h7BB3,4);
TASK_PP(16'h7BB4,4);
TASK_PP(16'h7BB5,4);
TASK_PP(16'h7BB6,4);
TASK_PP(16'h7BB7,4);
TASK_PP(16'h7BB8,4);
TASK_PP(16'h7BB9,4);
TASK_PP(16'h7BBA,4);
TASK_PP(16'h7BBB,4);
TASK_PP(16'h7BBC,4);
TASK_PP(16'h7BBD,4);
TASK_PP(16'h7BBE,4);
TASK_PP(16'h7BBF,4);
TASK_PP(16'h7BC0,4);
TASK_PP(16'h7BC1,4);
TASK_PP(16'h7BC2,4);
TASK_PP(16'h7BC3,4);
TASK_PP(16'h7BC4,4);
TASK_PP(16'h7BC5,4);
TASK_PP(16'h7BC6,4);
TASK_PP(16'h7BC7,4);
TASK_PP(16'h7BC8,4);
TASK_PP(16'h7BC9,4);
TASK_PP(16'h7BCA,4);
TASK_PP(16'h7BCB,4);
TASK_PP(16'h7BCC,4);
TASK_PP(16'h7BCD,4);
TASK_PP(16'h7BCE,4);
TASK_PP(16'h7BCF,4);
TASK_PP(16'h7BD0,4);
TASK_PP(16'h7BD1,4);
TASK_PP(16'h7BD2,4);
TASK_PP(16'h7BD3,4);
TASK_PP(16'h7BD4,4);
TASK_PP(16'h7BD5,4);
TASK_PP(16'h7BD6,4);
TASK_PP(16'h7BD7,4);
TASK_PP(16'h7BD8,4);
TASK_PP(16'h7BD9,4);
TASK_PP(16'h7BDA,4);
TASK_PP(16'h7BDB,4);
TASK_PP(16'h7BDC,4);
TASK_PP(16'h7BDD,4);
TASK_PP(16'h7BDE,4);
TASK_PP(16'h7BDF,4);
TASK_PP(16'h7BE0,4);
TASK_PP(16'h7BE1,4);
TASK_PP(16'h7BE2,4);
TASK_PP(16'h7BE3,4);
TASK_PP(16'h7BE4,4);
TASK_PP(16'h7BE5,4);
TASK_PP(16'h7BE6,4);
TASK_PP(16'h7BE7,4);
TASK_PP(16'h7BE8,4);
TASK_PP(16'h7BE9,4);
TASK_PP(16'h7BEA,4);
TASK_PP(16'h7BEB,4);
TASK_PP(16'h7BEC,4);
TASK_PP(16'h7BED,4);
TASK_PP(16'h7BEE,4);
TASK_PP(16'h7BEF,4);
TASK_PP(16'h7BF0,4);
TASK_PP(16'h7BF1,4);
TASK_PP(16'h7BF2,4);
TASK_PP(16'h7BF3,4);
TASK_PP(16'h7BF4,4);
TASK_PP(16'h7BF5,4);
TASK_PP(16'h7BF6,4);
TASK_PP(16'h7BF7,4);
TASK_PP(16'h7BF8,4);
TASK_PP(16'h7BF9,4);
TASK_PP(16'h7BFA,4);
TASK_PP(16'h7BFB,4);
TASK_PP(16'h7BFC,4);
TASK_PP(16'h7BFD,4);
TASK_PP(16'h7BFE,4);
TASK_PP(16'h7BFF,4);
TASK_PP(16'h7C00,4);
TASK_PP(16'h7C01,4);
TASK_PP(16'h7C02,4);
TASK_PP(16'h7C03,4);
TASK_PP(16'h7C04,4);
TASK_PP(16'h7C05,4);
TASK_PP(16'h7C06,4);
TASK_PP(16'h7C07,4);
TASK_PP(16'h7C08,4);
TASK_PP(16'h7C09,4);
TASK_PP(16'h7C0A,4);
TASK_PP(16'h7C0B,4);
TASK_PP(16'h7C0C,4);
TASK_PP(16'h7C0D,4);
TASK_PP(16'h7C0E,4);
TASK_PP(16'h7C0F,4);
TASK_PP(16'h7C10,4);
TASK_PP(16'h7C11,4);
TASK_PP(16'h7C12,4);
TASK_PP(16'h7C13,4);
TASK_PP(16'h7C14,4);
TASK_PP(16'h7C15,4);
TASK_PP(16'h7C16,4);
TASK_PP(16'h7C17,4);
TASK_PP(16'h7C18,4);
TASK_PP(16'h7C19,4);
TASK_PP(16'h7C1A,4);
TASK_PP(16'h7C1B,4);
TASK_PP(16'h7C1C,4);
TASK_PP(16'h7C1D,4);
TASK_PP(16'h7C1E,4);
TASK_PP(16'h7C1F,4);
TASK_PP(16'h7C20,4);
TASK_PP(16'h7C21,4);
TASK_PP(16'h7C22,4);
TASK_PP(16'h7C23,4);
TASK_PP(16'h7C24,4);
TASK_PP(16'h7C25,4);
TASK_PP(16'h7C26,4);
TASK_PP(16'h7C27,4);
TASK_PP(16'h7C28,4);
TASK_PP(16'h7C29,4);
TASK_PP(16'h7C2A,4);
TASK_PP(16'h7C2B,4);
TASK_PP(16'h7C2C,4);
TASK_PP(16'h7C2D,4);
TASK_PP(16'h7C2E,4);
TASK_PP(16'h7C2F,4);
TASK_PP(16'h7C30,4);
TASK_PP(16'h7C31,4);
TASK_PP(16'h7C32,4);
TASK_PP(16'h7C33,4);
TASK_PP(16'h7C34,4);
TASK_PP(16'h7C35,4);
TASK_PP(16'h7C36,4);
TASK_PP(16'h7C37,4);
TASK_PP(16'h7C38,4);
TASK_PP(16'h7C39,4);
TASK_PP(16'h7C3A,4);
TASK_PP(16'h7C3B,4);
TASK_PP(16'h7C3C,4);
TASK_PP(16'h7C3D,4);
TASK_PP(16'h7C3E,4);
TASK_PP(16'h7C3F,4);
TASK_PP(16'h7C40,4);
TASK_PP(16'h7C41,4);
TASK_PP(16'h7C42,4);
TASK_PP(16'h7C43,4);
TASK_PP(16'h7C44,4);
TASK_PP(16'h7C45,4);
TASK_PP(16'h7C46,4);
TASK_PP(16'h7C47,4);
TASK_PP(16'h7C48,4);
TASK_PP(16'h7C49,4);
TASK_PP(16'h7C4A,4);
TASK_PP(16'h7C4B,4);
TASK_PP(16'h7C4C,4);
TASK_PP(16'h7C4D,4);
TASK_PP(16'h7C4E,4);
TASK_PP(16'h7C4F,4);
TASK_PP(16'h7C50,4);
TASK_PP(16'h7C51,4);
TASK_PP(16'h7C52,4);
TASK_PP(16'h7C53,4);
TASK_PP(16'h7C54,4);
TASK_PP(16'h7C55,4);
TASK_PP(16'h7C56,4);
TASK_PP(16'h7C57,4);
TASK_PP(16'h7C58,4);
TASK_PP(16'h7C59,4);
TASK_PP(16'h7C5A,4);
TASK_PP(16'h7C5B,4);
TASK_PP(16'h7C5C,4);
TASK_PP(16'h7C5D,4);
TASK_PP(16'h7C5E,4);
TASK_PP(16'h7C5F,4);
TASK_PP(16'h7C60,4);
TASK_PP(16'h7C61,4);
TASK_PP(16'h7C62,4);
TASK_PP(16'h7C63,4);
TASK_PP(16'h7C64,4);
TASK_PP(16'h7C65,4);
TASK_PP(16'h7C66,4);
TASK_PP(16'h7C67,4);
TASK_PP(16'h7C68,4);
TASK_PP(16'h7C69,4);
TASK_PP(16'h7C6A,4);
TASK_PP(16'h7C6B,4);
TASK_PP(16'h7C6C,4);
TASK_PP(16'h7C6D,4);
TASK_PP(16'h7C6E,4);
TASK_PP(16'h7C6F,4);
TASK_PP(16'h7C70,4);
TASK_PP(16'h7C71,4);
TASK_PP(16'h7C72,4);
TASK_PP(16'h7C73,4);
TASK_PP(16'h7C74,4);
TASK_PP(16'h7C75,4);
TASK_PP(16'h7C76,4);
TASK_PP(16'h7C77,4);
TASK_PP(16'h7C78,4);
TASK_PP(16'h7C79,4);
TASK_PP(16'h7C7A,4);
TASK_PP(16'h7C7B,4);
TASK_PP(16'h7C7C,4);
TASK_PP(16'h7C7D,4);
TASK_PP(16'h7C7E,4);
TASK_PP(16'h7C7F,4);
TASK_PP(16'h7C80,4);
TASK_PP(16'h7C81,4);
TASK_PP(16'h7C82,4);
TASK_PP(16'h7C83,4);
TASK_PP(16'h7C84,4);
TASK_PP(16'h7C85,4);
TASK_PP(16'h7C86,4);
TASK_PP(16'h7C87,4);
TASK_PP(16'h7C88,4);
TASK_PP(16'h7C89,4);
TASK_PP(16'h7C8A,4);
TASK_PP(16'h7C8B,4);
TASK_PP(16'h7C8C,4);
TASK_PP(16'h7C8D,4);
TASK_PP(16'h7C8E,4);
TASK_PP(16'h7C8F,4);
TASK_PP(16'h7C90,4);
TASK_PP(16'h7C91,4);
TASK_PP(16'h7C92,4);
TASK_PP(16'h7C93,4);
TASK_PP(16'h7C94,4);
TASK_PP(16'h7C95,4);
TASK_PP(16'h7C96,4);
TASK_PP(16'h7C97,4);
TASK_PP(16'h7C98,4);
TASK_PP(16'h7C99,4);
TASK_PP(16'h7C9A,4);
TASK_PP(16'h7C9B,4);
TASK_PP(16'h7C9C,4);
TASK_PP(16'h7C9D,4);
TASK_PP(16'h7C9E,4);
TASK_PP(16'h7C9F,4);
TASK_PP(16'h7CA0,4);
TASK_PP(16'h7CA1,4);
TASK_PP(16'h7CA2,4);
TASK_PP(16'h7CA3,4);
TASK_PP(16'h7CA4,4);
TASK_PP(16'h7CA5,4);
TASK_PP(16'h7CA6,4);
TASK_PP(16'h7CA7,4);
TASK_PP(16'h7CA8,4);
TASK_PP(16'h7CA9,4);
TASK_PP(16'h7CAA,4);
TASK_PP(16'h7CAB,4);
TASK_PP(16'h7CAC,4);
TASK_PP(16'h7CAD,4);
TASK_PP(16'h7CAE,4);
TASK_PP(16'h7CAF,4);
TASK_PP(16'h7CB0,4);
TASK_PP(16'h7CB1,4);
TASK_PP(16'h7CB2,4);
TASK_PP(16'h7CB3,4);
TASK_PP(16'h7CB4,4);
TASK_PP(16'h7CB5,4);
TASK_PP(16'h7CB6,4);
TASK_PP(16'h7CB7,4);
TASK_PP(16'h7CB8,4);
TASK_PP(16'h7CB9,4);
TASK_PP(16'h7CBA,4);
TASK_PP(16'h7CBB,4);
TASK_PP(16'h7CBC,4);
TASK_PP(16'h7CBD,4);
TASK_PP(16'h7CBE,4);
TASK_PP(16'h7CBF,4);
TASK_PP(16'h7CC0,4);
TASK_PP(16'h7CC1,4);
TASK_PP(16'h7CC2,4);
TASK_PP(16'h7CC3,4);
TASK_PP(16'h7CC4,4);
TASK_PP(16'h7CC5,4);
TASK_PP(16'h7CC6,4);
TASK_PP(16'h7CC7,4);
TASK_PP(16'h7CC8,4);
TASK_PP(16'h7CC9,4);
TASK_PP(16'h7CCA,4);
TASK_PP(16'h7CCB,4);
TASK_PP(16'h7CCC,4);
TASK_PP(16'h7CCD,4);
TASK_PP(16'h7CCE,4);
TASK_PP(16'h7CCF,4);
TASK_PP(16'h7CD0,4);
TASK_PP(16'h7CD1,4);
TASK_PP(16'h7CD2,4);
TASK_PP(16'h7CD3,4);
TASK_PP(16'h7CD4,4);
TASK_PP(16'h7CD5,4);
TASK_PP(16'h7CD6,4);
TASK_PP(16'h7CD7,4);
TASK_PP(16'h7CD8,4);
TASK_PP(16'h7CD9,4);
TASK_PP(16'h7CDA,4);
TASK_PP(16'h7CDB,4);
TASK_PP(16'h7CDC,4);
TASK_PP(16'h7CDD,4);
TASK_PP(16'h7CDE,4);
TASK_PP(16'h7CDF,4);
TASK_PP(16'h7CE0,4);
TASK_PP(16'h7CE1,4);
TASK_PP(16'h7CE2,4);
TASK_PP(16'h7CE3,4);
TASK_PP(16'h7CE4,4);
TASK_PP(16'h7CE5,4);
TASK_PP(16'h7CE6,4);
TASK_PP(16'h7CE7,4);
TASK_PP(16'h7CE8,4);
TASK_PP(16'h7CE9,4);
TASK_PP(16'h7CEA,4);
TASK_PP(16'h7CEB,4);
TASK_PP(16'h7CEC,4);
TASK_PP(16'h7CED,4);
TASK_PP(16'h7CEE,4);
TASK_PP(16'h7CEF,4);
TASK_PP(16'h7CF0,4);
TASK_PP(16'h7CF1,4);
TASK_PP(16'h7CF2,4);
TASK_PP(16'h7CF3,4);
TASK_PP(16'h7CF4,4);
TASK_PP(16'h7CF5,4);
TASK_PP(16'h7CF6,4);
TASK_PP(16'h7CF7,4);
TASK_PP(16'h7CF8,4);
TASK_PP(16'h7CF9,4);
TASK_PP(16'h7CFA,4);
TASK_PP(16'h7CFB,4);
TASK_PP(16'h7CFC,4);
TASK_PP(16'h7CFD,4);
TASK_PP(16'h7CFE,4);
TASK_PP(16'h7CFF,4);
TASK_PP(16'h7D00,4);
TASK_PP(16'h7D01,4);
TASK_PP(16'h7D02,4);
TASK_PP(16'h7D03,4);
TASK_PP(16'h7D04,4);
TASK_PP(16'h7D05,4);
TASK_PP(16'h7D06,4);
TASK_PP(16'h7D07,4);
TASK_PP(16'h7D08,4);
TASK_PP(16'h7D09,4);
TASK_PP(16'h7D0A,4);
TASK_PP(16'h7D0B,4);
TASK_PP(16'h7D0C,4);
TASK_PP(16'h7D0D,4);
TASK_PP(16'h7D0E,4);
TASK_PP(16'h7D0F,4);
TASK_PP(16'h7D10,4);
TASK_PP(16'h7D11,4);
TASK_PP(16'h7D12,4);
TASK_PP(16'h7D13,4);
TASK_PP(16'h7D14,4);
TASK_PP(16'h7D15,4);
TASK_PP(16'h7D16,4);
TASK_PP(16'h7D17,4);
TASK_PP(16'h7D18,4);
TASK_PP(16'h7D19,4);
TASK_PP(16'h7D1A,4);
TASK_PP(16'h7D1B,4);
TASK_PP(16'h7D1C,4);
TASK_PP(16'h7D1D,4);
TASK_PP(16'h7D1E,4);
TASK_PP(16'h7D1F,4);
TASK_PP(16'h7D20,4);
TASK_PP(16'h7D21,4);
TASK_PP(16'h7D22,4);
TASK_PP(16'h7D23,4);
TASK_PP(16'h7D24,4);
TASK_PP(16'h7D25,4);
TASK_PP(16'h7D26,4);
TASK_PP(16'h7D27,4);
TASK_PP(16'h7D28,4);
TASK_PP(16'h7D29,4);
TASK_PP(16'h7D2A,4);
TASK_PP(16'h7D2B,4);
TASK_PP(16'h7D2C,4);
TASK_PP(16'h7D2D,4);
TASK_PP(16'h7D2E,4);
TASK_PP(16'h7D2F,4);
TASK_PP(16'h7D30,4);
TASK_PP(16'h7D31,4);
TASK_PP(16'h7D32,4);
TASK_PP(16'h7D33,4);
TASK_PP(16'h7D34,4);
TASK_PP(16'h7D35,4);
TASK_PP(16'h7D36,4);
TASK_PP(16'h7D37,4);
TASK_PP(16'h7D38,4);
TASK_PP(16'h7D39,4);
TASK_PP(16'h7D3A,4);
TASK_PP(16'h7D3B,4);
TASK_PP(16'h7D3C,4);
TASK_PP(16'h7D3D,4);
TASK_PP(16'h7D3E,4);
TASK_PP(16'h7D3F,4);
TASK_PP(16'h7D40,4);
TASK_PP(16'h7D41,4);
TASK_PP(16'h7D42,4);
TASK_PP(16'h7D43,4);
TASK_PP(16'h7D44,4);
TASK_PP(16'h7D45,4);
TASK_PP(16'h7D46,4);
TASK_PP(16'h7D47,4);
TASK_PP(16'h7D48,4);
TASK_PP(16'h7D49,4);
TASK_PP(16'h7D4A,4);
TASK_PP(16'h7D4B,4);
TASK_PP(16'h7D4C,4);
TASK_PP(16'h7D4D,4);
TASK_PP(16'h7D4E,4);
TASK_PP(16'h7D4F,4);
TASK_PP(16'h7D50,4);
TASK_PP(16'h7D51,4);
TASK_PP(16'h7D52,4);
TASK_PP(16'h7D53,4);
TASK_PP(16'h7D54,4);
TASK_PP(16'h7D55,4);
TASK_PP(16'h7D56,4);
TASK_PP(16'h7D57,4);
TASK_PP(16'h7D58,4);
TASK_PP(16'h7D59,4);
TASK_PP(16'h7D5A,4);
TASK_PP(16'h7D5B,4);
TASK_PP(16'h7D5C,4);
TASK_PP(16'h7D5D,4);
TASK_PP(16'h7D5E,4);
TASK_PP(16'h7D5F,4);
TASK_PP(16'h7D60,4);
TASK_PP(16'h7D61,4);
TASK_PP(16'h7D62,4);
TASK_PP(16'h7D63,4);
TASK_PP(16'h7D64,4);
TASK_PP(16'h7D65,4);
TASK_PP(16'h7D66,4);
TASK_PP(16'h7D67,4);
TASK_PP(16'h7D68,4);
TASK_PP(16'h7D69,4);
TASK_PP(16'h7D6A,4);
TASK_PP(16'h7D6B,4);
TASK_PP(16'h7D6C,4);
TASK_PP(16'h7D6D,4);
TASK_PP(16'h7D6E,4);
TASK_PP(16'h7D6F,4);
TASK_PP(16'h7D70,4);
TASK_PP(16'h7D71,4);
TASK_PP(16'h7D72,4);
TASK_PP(16'h7D73,4);
TASK_PP(16'h7D74,4);
TASK_PP(16'h7D75,4);
TASK_PP(16'h7D76,4);
TASK_PP(16'h7D77,4);
TASK_PP(16'h7D78,4);
TASK_PP(16'h7D79,4);
TASK_PP(16'h7D7A,4);
TASK_PP(16'h7D7B,4);
TASK_PP(16'h7D7C,4);
TASK_PP(16'h7D7D,4);
TASK_PP(16'h7D7E,4);
TASK_PP(16'h7D7F,4);
TASK_PP(16'h7D80,4);
TASK_PP(16'h7D81,4);
TASK_PP(16'h7D82,4);
TASK_PP(16'h7D83,4);
TASK_PP(16'h7D84,4);
TASK_PP(16'h7D85,4);
TASK_PP(16'h7D86,4);
TASK_PP(16'h7D87,4);
TASK_PP(16'h7D88,4);
TASK_PP(16'h7D89,4);
TASK_PP(16'h7D8A,4);
TASK_PP(16'h7D8B,4);
TASK_PP(16'h7D8C,4);
TASK_PP(16'h7D8D,4);
TASK_PP(16'h7D8E,4);
TASK_PP(16'h7D8F,4);
TASK_PP(16'h7D90,4);
TASK_PP(16'h7D91,4);
TASK_PP(16'h7D92,4);
TASK_PP(16'h7D93,4);
TASK_PP(16'h7D94,4);
TASK_PP(16'h7D95,4);
TASK_PP(16'h7D96,4);
TASK_PP(16'h7D97,4);
TASK_PP(16'h7D98,4);
TASK_PP(16'h7D99,4);
TASK_PP(16'h7D9A,4);
TASK_PP(16'h7D9B,4);
TASK_PP(16'h7D9C,4);
TASK_PP(16'h7D9D,4);
TASK_PP(16'h7D9E,4);
TASK_PP(16'h7D9F,4);
TASK_PP(16'h7DA0,4);
TASK_PP(16'h7DA1,4);
TASK_PP(16'h7DA2,4);
TASK_PP(16'h7DA3,4);
TASK_PP(16'h7DA4,4);
TASK_PP(16'h7DA5,4);
TASK_PP(16'h7DA6,4);
TASK_PP(16'h7DA7,4);
TASK_PP(16'h7DA8,4);
TASK_PP(16'h7DA9,4);
TASK_PP(16'h7DAA,4);
TASK_PP(16'h7DAB,4);
TASK_PP(16'h7DAC,4);
TASK_PP(16'h7DAD,4);
TASK_PP(16'h7DAE,4);
TASK_PP(16'h7DAF,4);
TASK_PP(16'h7DB0,4);
TASK_PP(16'h7DB1,4);
TASK_PP(16'h7DB2,4);
TASK_PP(16'h7DB3,4);
TASK_PP(16'h7DB4,4);
TASK_PP(16'h7DB5,4);
TASK_PP(16'h7DB6,4);
TASK_PP(16'h7DB7,4);
TASK_PP(16'h7DB8,4);
TASK_PP(16'h7DB9,4);
TASK_PP(16'h7DBA,4);
TASK_PP(16'h7DBB,4);
TASK_PP(16'h7DBC,4);
TASK_PP(16'h7DBD,4);
TASK_PP(16'h7DBE,4);
TASK_PP(16'h7DBF,4);
TASK_PP(16'h7DC0,4);
TASK_PP(16'h7DC1,4);
TASK_PP(16'h7DC2,4);
TASK_PP(16'h7DC3,4);
TASK_PP(16'h7DC4,4);
TASK_PP(16'h7DC5,4);
TASK_PP(16'h7DC6,4);
TASK_PP(16'h7DC7,4);
TASK_PP(16'h7DC8,4);
TASK_PP(16'h7DC9,4);
TASK_PP(16'h7DCA,4);
TASK_PP(16'h7DCB,4);
TASK_PP(16'h7DCC,4);
TASK_PP(16'h7DCD,4);
TASK_PP(16'h7DCE,4);
TASK_PP(16'h7DCF,4);
TASK_PP(16'h7DD0,4);
TASK_PP(16'h7DD1,4);
TASK_PP(16'h7DD2,4);
TASK_PP(16'h7DD3,4);
TASK_PP(16'h7DD4,4);
TASK_PP(16'h7DD5,4);
TASK_PP(16'h7DD6,4);
TASK_PP(16'h7DD7,4);
TASK_PP(16'h7DD8,4);
TASK_PP(16'h7DD9,4);
TASK_PP(16'h7DDA,4);
TASK_PP(16'h7DDB,4);
TASK_PP(16'h7DDC,4);
TASK_PP(16'h7DDD,4);
TASK_PP(16'h7DDE,4);
TASK_PP(16'h7DDF,4);
TASK_PP(16'h7DE0,4);
TASK_PP(16'h7DE1,4);
TASK_PP(16'h7DE2,4);
TASK_PP(16'h7DE3,4);
TASK_PP(16'h7DE4,4);
TASK_PP(16'h7DE5,4);
TASK_PP(16'h7DE6,4);
TASK_PP(16'h7DE7,4);
TASK_PP(16'h7DE8,4);
TASK_PP(16'h7DE9,4);
TASK_PP(16'h7DEA,4);
TASK_PP(16'h7DEB,4);
TASK_PP(16'h7DEC,4);
TASK_PP(16'h7DED,4);
TASK_PP(16'h7DEE,4);
TASK_PP(16'h7DEF,4);
TASK_PP(16'h7DF0,4);
TASK_PP(16'h7DF1,4);
TASK_PP(16'h7DF2,4);
TASK_PP(16'h7DF3,4);
TASK_PP(16'h7DF4,4);
TASK_PP(16'h7DF5,4);
TASK_PP(16'h7DF6,4);
TASK_PP(16'h7DF7,4);
TASK_PP(16'h7DF8,4);
TASK_PP(16'h7DF9,4);
TASK_PP(16'h7DFA,4);
TASK_PP(16'h7DFB,4);
TASK_PP(16'h7DFC,4);
TASK_PP(16'h7DFD,4);
TASK_PP(16'h7DFE,4);
TASK_PP(16'h7DFF,4);
TASK_PP(16'h7E00,4);
TASK_PP(16'h7E01,4);
TASK_PP(16'h7E02,4);
TASK_PP(16'h7E03,4);
TASK_PP(16'h7E04,4);
TASK_PP(16'h7E05,4);
TASK_PP(16'h7E06,4);
TASK_PP(16'h7E07,4);
TASK_PP(16'h7E08,4);
TASK_PP(16'h7E09,4);
TASK_PP(16'h7E0A,4);
TASK_PP(16'h7E0B,4);
TASK_PP(16'h7E0C,4);
TASK_PP(16'h7E0D,4);
TASK_PP(16'h7E0E,4);
TASK_PP(16'h7E0F,4);
TASK_PP(16'h7E10,4);
TASK_PP(16'h7E11,4);
TASK_PP(16'h7E12,4);
TASK_PP(16'h7E13,4);
TASK_PP(16'h7E14,4);
TASK_PP(16'h7E15,4);
TASK_PP(16'h7E16,4);
TASK_PP(16'h7E17,4);
TASK_PP(16'h7E18,4);
TASK_PP(16'h7E19,4);
TASK_PP(16'h7E1A,4);
TASK_PP(16'h7E1B,4);
TASK_PP(16'h7E1C,4);
TASK_PP(16'h7E1D,4);
TASK_PP(16'h7E1E,4);
TASK_PP(16'h7E1F,4);
TASK_PP(16'h7E20,4);
TASK_PP(16'h7E21,4);
TASK_PP(16'h7E22,4);
TASK_PP(16'h7E23,4);
TASK_PP(16'h7E24,4);
TASK_PP(16'h7E25,4);
TASK_PP(16'h7E26,4);
TASK_PP(16'h7E27,4);
TASK_PP(16'h7E28,4);
TASK_PP(16'h7E29,4);
TASK_PP(16'h7E2A,4);
TASK_PP(16'h7E2B,4);
TASK_PP(16'h7E2C,4);
TASK_PP(16'h7E2D,4);
TASK_PP(16'h7E2E,4);
TASK_PP(16'h7E2F,4);
TASK_PP(16'h7E30,4);
TASK_PP(16'h7E31,4);
TASK_PP(16'h7E32,4);
TASK_PP(16'h7E33,4);
TASK_PP(16'h7E34,4);
TASK_PP(16'h7E35,4);
TASK_PP(16'h7E36,4);
TASK_PP(16'h7E37,4);
TASK_PP(16'h7E38,4);
TASK_PP(16'h7E39,4);
TASK_PP(16'h7E3A,4);
TASK_PP(16'h7E3B,4);
TASK_PP(16'h7E3C,4);
TASK_PP(16'h7E3D,4);
TASK_PP(16'h7E3E,4);
TASK_PP(16'h7E3F,4);
TASK_PP(16'h7E40,4);
TASK_PP(16'h7E41,4);
TASK_PP(16'h7E42,4);
TASK_PP(16'h7E43,4);
TASK_PP(16'h7E44,4);
TASK_PP(16'h7E45,4);
TASK_PP(16'h7E46,4);
TASK_PP(16'h7E47,4);
TASK_PP(16'h7E48,4);
TASK_PP(16'h7E49,4);
TASK_PP(16'h7E4A,4);
TASK_PP(16'h7E4B,4);
TASK_PP(16'h7E4C,4);
TASK_PP(16'h7E4D,4);
TASK_PP(16'h7E4E,4);
TASK_PP(16'h7E4F,4);
TASK_PP(16'h7E50,4);
TASK_PP(16'h7E51,4);
TASK_PP(16'h7E52,4);
TASK_PP(16'h7E53,4);
TASK_PP(16'h7E54,4);
TASK_PP(16'h7E55,4);
TASK_PP(16'h7E56,4);
TASK_PP(16'h7E57,4);
TASK_PP(16'h7E58,4);
TASK_PP(16'h7E59,4);
TASK_PP(16'h7E5A,4);
TASK_PP(16'h7E5B,4);
TASK_PP(16'h7E5C,4);
TASK_PP(16'h7E5D,4);
TASK_PP(16'h7E5E,4);
TASK_PP(16'h7E5F,4);
TASK_PP(16'h7E60,4);
TASK_PP(16'h7E61,4);
TASK_PP(16'h7E62,4);
TASK_PP(16'h7E63,4);
TASK_PP(16'h7E64,4);
TASK_PP(16'h7E65,4);
TASK_PP(16'h7E66,4);
TASK_PP(16'h7E67,4);
TASK_PP(16'h7E68,4);
TASK_PP(16'h7E69,4);
TASK_PP(16'h7E6A,4);
TASK_PP(16'h7E6B,4);
TASK_PP(16'h7E6C,4);
TASK_PP(16'h7E6D,4);
TASK_PP(16'h7E6E,4);
TASK_PP(16'h7E6F,4);
TASK_PP(16'h7E70,4);
TASK_PP(16'h7E71,4);
TASK_PP(16'h7E72,4);
TASK_PP(16'h7E73,4);
TASK_PP(16'h7E74,4);
TASK_PP(16'h7E75,4);
TASK_PP(16'h7E76,4);
TASK_PP(16'h7E77,4);
TASK_PP(16'h7E78,4);
TASK_PP(16'h7E79,4);
TASK_PP(16'h7E7A,4);
TASK_PP(16'h7E7B,4);
TASK_PP(16'h7E7C,4);
TASK_PP(16'h7E7D,4);
TASK_PP(16'h7E7E,4);
TASK_PP(16'h7E7F,4);
TASK_PP(16'h7E80,4);
TASK_PP(16'h7E81,4);
TASK_PP(16'h7E82,4);
TASK_PP(16'h7E83,4);
TASK_PP(16'h7E84,4);
TASK_PP(16'h7E85,4);
TASK_PP(16'h7E86,4);
TASK_PP(16'h7E87,4);
TASK_PP(16'h7E88,4);
TASK_PP(16'h7E89,4);
TASK_PP(16'h7E8A,4);
TASK_PP(16'h7E8B,4);
TASK_PP(16'h7E8C,4);
TASK_PP(16'h7E8D,4);
TASK_PP(16'h7E8E,4);
TASK_PP(16'h7E8F,4);
TASK_PP(16'h7E90,4);
TASK_PP(16'h7E91,4);
TASK_PP(16'h7E92,4);
TASK_PP(16'h7E93,4);
TASK_PP(16'h7E94,4);
TASK_PP(16'h7E95,4);
TASK_PP(16'h7E96,4);
TASK_PP(16'h7E97,4);
TASK_PP(16'h7E98,4);
TASK_PP(16'h7E99,4);
TASK_PP(16'h7E9A,4);
TASK_PP(16'h7E9B,4);
TASK_PP(16'h7E9C,4);
TASK_PP(16'h7E9D,4);
TASK_PP(16'h7E9E,4);
TASK_PP(16'h7E9F,4);
TASK_PP(16'h7EA0,4);
TASK_PP(16'h7EA1,4);
TASK_PP(16'h7EA2,4);
TASK_PP(16'h7EA3,4);
TASK_PP(16'h7EA4,4);
TASK_PP(16'h7EA5,4);
TASK_PP(16'h7EA6,4);
TASK_PP(16'h7EA7,4);
TASK_PP(16'h7EA8,4);
TASK_PP(16'h7EA9,4);
TASK_PP(16'h7EAA,4);
TASK_PP(16'h7EAB,4);
TASK_PP(16'h7EAC,4);
TASK_PP(16'h7EAD,4);
TASK_PP(16'h7EAE,4);
TASK_PP(16'h7EAF,4);
TASK_PP(16'h7EB0,4);
TASK_PP(16'h7EB1,4);
TASK_PP(16'h7EB2,4);
TASK_PP(16'h7EB3,4);
TASK_PP(16'h7EB4,4);
TASK_PP(16'h7EB5,4);
TASK_PP(16'h7EB6,4);
TASK_PP(16'h7EB7,4);
TASK_PP(16'h7EB8,4);
TASK_PP(16'h7EB9,4);
TASK_PP(16'h7EBA,4);
TASK_PP(16'h7EBB,4);
TASK_PP(16'h7EBC,4);
TASK_PP(16'h7EBD,4);
TASK_PP(16'h7EBE,4);
TASK_PP(16'h7EBF,4);
TASK_PP(16'h7EC0,4);
TASK_PP(16'h7EC1,4);
TASK_PP(16'h7EC2,4);
TASK_PP(16'h7EC3,4);
TASK_PP(16'h7EC4,4);
TASK_PP(16'h7EC5,4);
TASK_PP(16'h7EC6,4);
TASK_PP(16'h7EC7,4);
TASK_PP(16'h7EC8,4);
TASK_PP(16'h7EC9,4);
TASK_PP(16'h7ECA,4);
TASK_PP(16'h7ECB,4);
TASK_PP(16'h7ECC,4);
TASK_PP(16'h7ECD,4);
TASK_PP(16'h7ECE,4);
TASK_PP(16'h7ECF,4);
TASK_PP(16'h7ED0,4);
TASK_PP(16'h7ED1,4);
TASK_PP(16'h7ED2,4);
TASK_PP(16'h7ED3,4);
TASK_PP(16'h7ED4,4);
TASK_PP(16'h7ED5,4);
TASK_PP(16'h7ED6,4);
TASK_PP(16'h7ED7,4);
TASK_PP(16'h7ED8,4);
TASK_PP(16'h7ED9,4);
TASK_PP(16'h7EDA,4);
TASK_PP(16'h7EDB,4);
TASK_PP(16'h7EDC,4);
TASK_PP(16'h7EDD,4);
TASK_PP(16'h7EDE,4);
TASK_PP(16'h7EDF,4);
TASK_PP(16'h7EE0,4);
TASK_PP(16'h7EE1,4);
TASK_PP(16'h7EE2,4);
TASK_PP(16'h7EE3,4);
TASK_PP(16'h7EE4,4);
TASK_PP(16'h7EE5,4);
TASK_PP(16'h7EE6,4);
TASK_PP(16'h7EE7,4);
TASK_PP(16'h7EE8,4);
TASK_PP(16'h7EE9,4);
TASK_PP(16'h7EEA,4);
TASK_PP(16'h7EEB,4);
TASK_PP(16'h7EEC,4);
TASK_PP(16'h7EED,4);
TASK_PP(16'h7EEE,4);
TASK_PP(16'h7EEF,4);
TASK_PP(16'h7EF0,4);
TASK_PP(16'h7EF1,4);
TASK_PP(16'h7EF2,4);
TASK_PP(16'h7EF3,4);
TASK_PP(16'h7EF4,4);
TASK_PP(16'h7EF5,4);
TASK_PP(16'h7EF6,4);
TASK_PP(16'h7EF7,4);
TASK_PP(16'h7EF8,4);
TASK_PP(16'h7EF9,4);
TASK_PP(16'h7EFA,4);
TASK_PP(16'h7EFB,4);
TASK_PP(16'h7EFC,4);
TASK_PP(16'h7EFD,4);
TASK_PP(16'h7EFE,4);
TASK_PP(16'h7EFF,4);
TASK_PP(16'h7F00,4);
TASK_PP(16'h7F01,4);
TASK_PP(16'h7F02,4);
TASK_PP(16'h7F03,4);
TASK_PP(16'h7F04,4);
TASK_PP(16'h7F05,4);
TASK_PP(16'h7F06,4);
TASK_PP(16'h7F07,4);
TASK_PP(16'h7F08,4);
TASK_PP(16'h7F09,4);
TASK_PP(16'h7F0A,4);
TASK_PP(16'h7F0B,4);
TASK_PP(16'h7F0C,4);
TASK_PP(16'h7F0D,4);
TASK_PP(16'h7F0E,4);
TASK_PP(16'h7F0F,4);
TASK_PP(16'h7F10,4);
TASK_PP(16'h7F11,4);
TASK_PP(16'h7F12,4);
TASK_PP(16'h7F13,4);
TASK_PP(16'h7F14,4);
TASK_PP(16'h7F15,4);
TASK_PP(16'h7F16,4);
TASK_PP(16'h7F17,4);
TASK_PP(16'h7F18,4);
TASK_PP(16'h7F19,4);
TASK_PP(16'h7F1A,4);
TASK_PP(16'h7F1B,4);
TASK_PP(16'h7F1C,4);
TASK_PP(16'h7F1D,4);
TASK_PP(16'h7F1E,4);
TASK_PP(16'h7F1F,4);
TASK_PP(16'h7F20,4);
TASK_PP(16'h7F21,4);
TASK_PP(16'h7F22,4);
TASK_PP(16'h7F23,4);
TASK_PP(16'h7F24,4);
TASK_PP(16'h7F25,4);
TASK_PP(16'h7F26,4);
TASK_PP(16'h7F27,4);
TASK_PP(16'h7F28,4);
TASK_PP(16'h7F29,4);
TASK_PP(16'h7F2A,4);
TASK_PP(16'h7F2B,4);
TASK_PP(16'h7F2C,4);
TASK_PP(16'h7F2D,4);
TASK_PP(16'h7F2E,4);
TASK_PP(16'h7F2F,4);
TASK_PP(16'h7F30,4);
TASK_PP(16'h7F31,4);
TASK_PP(16'h7F32,4);
TASK_PP(16'h7F33,4);
TASK_PP(16'h7F34,4);
TASK_PP(16'h7F35,4);
TASK_PP(16'h7F36,4);
TASK_PP(16'h7F37,4);
TASK_PP(16'h7F38,4);
TASK_PP(16'h7F39,4);
TASK_PP(16'h7F3A,4);
TASK_PP(16'h7F3B,4);
TASK_PP(16'h7F3C,4);
TASK_PP(16'h7F3D,4);
TASK_PP(16'h7F3E,4);
TASK_PP(16'h7F3F,4);
TASK_PP(16'h7F40,4);
TASK_PP(16'h7F41,4);
TASK_PP(16'h7F42,4);
TASK_PP(16'h7F43,4);
TASK_PP(16'h7F44,4);
TASK_PP(16'h7F45,4);
TASK_PP(16'h7F46,4);
TASK_PP(16'h7F47,4);
TASK_PP(16'h7F48,4);
TASK_PP(16'h7F49,4);
TASK_PP(16'h7F4A,4);
TASK_PP(16'h7F4B,4);
TASK_PP(16'h7F4C,4);
TASK_PP(16'h7F4D,4);
TASK_PP(16'h7F4E,4);
TASK_PP(16'h7F4F,4);
TASK_PP(16'h7F50,4);
TASK_PP(16'h7F51,4);
TASK_PP(16'h7F52,4);
TASK_PP(16'h7F53,4);
TASK_PP(16'h7F54,4);
TASK_PP(16'h7F55,4);
TASK_PP(16'h7F56,4);
TASK_PP(16'h7F57,4);
TASK_PP(16'h7F58,4);
TASK_PP(16'h7F59,4);
TASK_PP(16'h7F5A,4);
TASK_PP(16'h7F5B,4);
TASK_PP(16'h7F5C,4);
TASK_PP(16'h7F5D,4);
TASK_PP(16'h7F5E,4);
TASK_PP(16'h7F5F,4);
TASK_PP(16'h7F60,4);
TASK_PP(16'h7F61,4);
TASK_PP(16'h7F62,4);
TASK_PP(16'h7F63,4);
TASK_PP(16'h7F64,4);
TASK_PP(16'h7F65,4);
TASK_PP(16'h7F66,4);
TASK_PP(16'h7F67,4);
TASK_PP(16'h7F68,4);
TASK_PP(16'h7F69,4);
TASK_PP(16'h7F6A,4);
TASK_PP(16'h7F6B,4);
TASK_PP(16'h7F6C,4);
TASK_PP(16'h7F6D,4);
TASK_PP(16'h7F6E,4);
TASK_PP(16'h7F6F,4);
TASK_PP(16'h7F70,4);
TASK_PP(16'h7F71,4);
TASK_PP(16'h7F72,4);
TASK_PP(16'h7F73,4);
TASK_PP(16'h7F74,4);
TASK_PP(16'h7F75,4);
TASK_PP(16'h7F76,4);
TASK_PP(16'h7F77,4);
TASK_PP(16'h7F78,4);
TASK_PP(16'h7F79,4);
TASK_PP(16'h7F7A,4);
TASK_PP(16'h7F7B,4);
TASK_PP(16'h7F7C,4);
TASK_PP(16'h7F7D,4);
TASK_PP(16'h7F7E,4);
TASK_PP(16'h7F7F,4);
TASK_PP(16'h7F80,4);
TASK_PP(16'h7F81,4);
TASK_PP(16'h7F82,4);
TASK_PP(16'h7F83,4);
TASK_PP(16'h7F84,4);
TASK_PP(16'h7F85,4);
TASK_PP(16'h7F86,4);
TASK_PP(16'h7F87,4);
TASK_PP(16'h7F88,4);
TASK_PP(16'h7F89,4);
TASK_PP(16'h7F8A,4);
TASK_PP(16'h7F8B,4);
TASK_PP(16'h7F8C,4);
TASK_PP(16'h7F8D,4);
TASK_PP(16'h7F8E,4);
TASK_PP(16'h7F8F,4);
TASK_PP(16'h7F90,4);
TASK_PP(16'h7F91,4);
TASK_PP(16'h7F92,4);
TASK_PP(16'h7F93,4);
TASK_PP(16'h7F94,4);
TASK_PP(16'h7F95,4);
TASK_PP(16'h7F96,4);
TASK_PP(16'h7F97,4);
TASK_PP(16'h7F98,4);
TASK_PP(16'h7F99,4);
TASK_PP(16'h7F9A,4);
TASK_PP(16'h7F9B,4);
TASK_PP(16'h7F9C,4);
TASK_PP(16'h7F9D,4);
TASK_PP(16'h7F9E,4);
TASK_PP(16'h7F9F,4);
TASK_PP(16'h7FA0,4);
TASK_PP(16'h7FA1,4);
TASK_PP(16'h7FA2,4);
TASK_PP(16'h7FA3,4);
TASK_PP(16'h7FA4,4);
TASK_PP(16'h7FA5,4);
TASK_PP(16'h7FA6,4);
TASK_PP(16'h7FA7,4);
TASK_PP(16'h7FA8,4);
TASK_PP(16'h7FA9,4);
TASK_PP(16'h7FAA,4);
TASK_PP(16'h7FAB,4);
TASK_PP(16'h7FAC,4);
TASK_PP(16'h7FAD,4);
TASK_PP(16'h7FAE,4);
TASK_PP(16'h7FAF,4);
TASK_PP(16'h7FB0,4);
TASK_PP(16'h7FB1,4);
TASK_PP(16'h7FB2,4);
TASK_PP(16'h7FB3,4);
TASK_PP(16'h7FB4,4);
TASK_PP(16'h7FB5,4);
TASK_PP(16'h7FB6,4);
TASK_PP(16'h7FB7,4);
TASK_PP(16'h7FB8,4);
TASK_PP(16'h7FB9,4);
TASK_PP(16'h7FBA,4);
TASK_PP(16'h7FBB,4);
TASK_PP(16'h7FBC,4);
TASK_PP(16'h7FBD,4);
TASK_PP(16'h7FBE,4);
TASK_PP(16'h7FBF,4);
TASK_PP(16'h7FC0,4);
TASK_PP(16'h7FC1,4);
TASK_PP(16'h7FC2,4);
TASK_PP(16'h7FC3,4);
TASK_PP(16'h7FC4,4);
TASK_PP(16'h7FC5,4);
TASK_PP(16'h7FC6,4);
TASK_PP(16'h7FC7,4);
TASK_PP(16'h7FC8,4);
TASK_PP(16'h7FC9,4);
TASK_PP(16'h7FCA,4);
TASK_PP(16'h7FCB,4);
TASK_PP(16'h7FCC,4);
TASK_PP(16'h7FCD,4);
TASK_PP(16'h7FCE,4);
TASK_PP(16'h7FCF,4);
TASK_PP(16'h7FD0,4);
TASK_PP(16'h7FD1,4);
TASK_PP(16'h7FD2,4);
TASK_PP(16'h7FD3,4);
TASK_PP(16'h7FD4,4);
TASK_PP(16'h7FD5,4);
TASK_PP(16'h7FD6,4);
TASK_PP(16'h7FD7,4);
TASK_PP(16'h7FD8,4);
TASK_PP(16'h7FD9,4);
TASK_PP(16'h7FDA,4);
TASK_PP(16'h7FDB,4);
TASK_PP(16'h7FDC,4);
TASK_PP(16'h7FDD,4);
TASK_PP(16'h7FDE,4);
TASK_PP(16'h7FDF,4);
TASK_PP(16'h7FE0,4);
TASK_PP(16'h7FE1,4);
TASK_PP(16'h7FE2,4);
TASK_PP(16'h7FE3,4);
TASK_PP(16'h7FE4,4);
TASK_PP(16'h7FE5,4);
TASK_PP(16'h7FE6,4);
TASK_PP(16'h7FE7,4);
TASK_PP(16'h7FE8,4);
TASK_PP(16'h7FE9,4);
TASK_PP(16'h7FEA,4);
TASK_PP(16'h7FEB,4);
TASK_PP(16'h7FEC,4);
TASK_PP(16'h7FED,4);
TASK_PP(16'h7FEE,4);
TASK_PP(16'h7FEF,4);
TASK_PP(16'h7FF0,4);
TASK_PP(16'h7FF1,4);
TASK_PP(16'h7FF2,4);
TASK_PP(16'h7FF3,4);
TASK_PP(16'h7FF4,4);
TASK_PP(16'h7FF5,4);
TASK_PP(16'h7FF6,4);
TASK_PP(16'h7FF7,4);
TASK_PP(16'h7FF8,4);
TASK_PP(16'h7FF9,4);
TASK_PP(16'h7FFA,4);
TASK_PP(16'h7FFB,4);
TASK_PP(16'h7FFC,4);
TASK_PP(16'h7FFD,4);
TASK_PP(16'h7FFE,4);
TASK_PP(16'h7FFF,4);
TASK_PP(16'h8000,4);
TASK_PP(16'h8001,4);
TASK_PP(16'h8002,4);
TASK_PP(16'h8003,4);
TASK_PP(16'h8004,4);
TASK_PP(16'h8005,4);
TASK_PP(16'h8006,4);
TASK_PP(16'h8007,4);
TASK_PP(16'h8008,4);
TASK_PP(16'h8009,4);
TASK_PP(16'h800A,4);
TASK_PP(16'h800B,4);
TASK_PP(16'h800C,4);
TASK_PP(16'h800D,4);
TASK_PP(16'h800E,4);
TASK_PP(16'h800F,4);
TASK_PP(16'h8010,4);
TASK_PP(16'h8011,4);
TASK_PP(16'h8012,4);
TASK_PP(16'h8013,4);
TASK_PP(16'h8014,4);
TASK_PP(16'h8015,4);
TASK_PP(16'h8016,4);
TASK_PP(16'h8017,4);
TASK_PP(16'h8018,4);
TASK_PP(16'h8019,4);
TASK_PP(16'h801A,4);
TASK_PP(16'h801B,4);
TASK_PP(16'h801C,4);
TASK_PP(16'h801D,4);
TASK_PP(16'h801E,4);
TASK_PP(16'h801F,4);
TASK_PP(16'h8020,4);
TASK_PP(16'h8021,4);
TASK_PP(16'h8022,4);
TASK_PP(16'h8023,4);
TASK_PP(16'h8024,4);
TASK_PP(16'h8025,4);
TASK_PP(16'h8026,4);
TASK_PP(16'h8027,4);
TASK_PP(16'h8028,4);
TASK_PP(16'h8029,4);
TASK_PP(16'h802A,4);
TASK_PP(16'h802B,4);
TASK_PP(16'h802C,4);
TASK_PP(16'h802D,4);
TASK_PP(16'h802E,4);
TASK_PP(16'h802F,4);
TASK_PP(16'h8030,4);
TASK_PP(16'h8031,4);
TASK_PP(16'h8032,4);
TASK_PP(16'h8033,4);
TASK_PP(16'h8034,4);
TASK_PP(16'h8035,4);
TASK_PP(16'h8036,4);
TASK_PP(16'h8037,4);
TASK_PP(16'h8038,4);
TASK_PP(16'h8039,4);
TASK_PP(16'h803A,4);
TASK_PP(16'h803B,4);
TASK_PP(16'h803C,4);
TASK_PP(16'h803D,4);
TASK_PP(16'h803E,4);
TASK_PP(16'h803F,4);
TASK_PP(16'h8040,4);
TASK_PP(16'h8041,4);
TASK_PP(16'h8042,4);
TASK_PP(16'h8043,4);
TASK_PP(16'h8044,4);
TASK_PP(16'h8045,4);
TASK_PP(16'h8046,4);
TASK_PP(16'h8047,4);
TASK_PP(16'h8048,4);
TASK_PP(16'h8049,4);
TASK_PP(16'h804A,4);
TASK_PP(16'h804B,4);
TASK_PP(16'h804C,4);
TASK_PP(16'h804D,4);
TASK_PP(16'h804E,4);
TASK_PP(16'h804F,4);
TASK_PP(16'h8050,4);
TASK_PP(16'h8051,4);
TASK_PP(16'h8052,4);
TASK_PP(16'h8053,4);
TASK_PP(16'h8054,4);
TASK_PP(16'h8055,4);
TASK_PP(16'h8056,4);
TASK_PP(16'h8057,4);
TASK_PP(16'h8058,4);
TASK_PP(16'h8059,4);
TASK_PP(16'h805A,4);
TASK_PP(16'h805B,4);
TASK_PP(16'h805C,4);
TASK_PP(16'h805D,4);
TASK_PP(16'h805E,4);
TASK_PP(16'h805F,4);
TASK_PP(16'h8060,4);
TASK_PP(16'h8061,4);
TASK_PP(16'h8062,4);
TASK_PP(16'h8063,4);
TASK_PP(16'h8064,4);
TASK_PP(16'h8065,4);
TASK_PP(16'h8066,4);
TASK_PP(16'h8067,4);
TASK_PP(16'h8068,4);
TASK_PP(16'h8069,4);
TASK_PP(16'h806A,4);
TASK_PP(16'h806B,4);
TASK_PP(16'h806C,4);
TASK_PP(16'h806D,4);
TASK_PP(16'h806E,4);
TASK_PP(16'h806F,4);
TASK_PP(16'h8070,4);
TASK_PP(16'h8071,4);
TASK_PP(16'h8072,4);
TASK_PP(16'h8073,4);
TASK_PP(16'h8074,4);
TASK_PP(16'h8075,4);
TASK_PP(16'h8076,4);
TASK_PP(16'h8077,4);
TASK_PP(16'h8078,4);
TASK_PP(16'h8079,4);
TASK_PP(16'h807A,4);
TASK_PP(16'h807B,4);
TASK_PP(16'h807C,4);
TASK_PP(16'h807D,4);
TASK_PP(16'h807E,4);
TASK_PP(16'h807F,4);
TASK_PP(16'h8080,4);
TASK_PP(16'h8081,4);
TASK_PP(16'h8082,4);
TASK_PP(16'h8083,4);
TASK_PP(16'h8084,4);
TASK_PP(16'h8085,4);
TASK_PP(16'h8086,4);
TASK_PP(16'h8087,4);
TASK_PP(16'h8088,4);
TASK_PP(16'h8089,4);
TASK_PP(16'h808A,4);
TASK_PP(16'h808B,4);
TASK_PP(16'h808C,4);
TASK_PP(16'h808D,4);
TASK_PP(16'h808E,4);
TASK_PP(16'h808F,4);
TASK_PP(16'h8090,4);
TASK_PP(16'h8091,4);
TASK_PP(16'h8092,4);
TASK_PP(16'h8093,4);
TASK_PP(16'h8094,4);
TASK_PP(16'h8095,4);
TASK_PP(16'h8096,4);
TASK_PP(16'h8097,4);
TASK_PP(16'h8098,4);
TASK_PP(16'h8099,4);
TASK_PP(16'h809A,4);
TASK_PP(16'h809B,4);
TASK_PP(16'h809C,4);
TASK_PP(16'h809D,4);
TASK_PP(16'h809E,4);
TASK_PP(16'h809F,4);
TASK_PP(16'h80A0,4);
TASK_PP(16'h80A1,4);
TASK_PP(16'h80A2,4);
TASK_PP(16'h80A3,4);
TASK_PP(16'h80A4,4);
TASK_PP(16'h80A5,4);
TASK_PP(16'h80A6,4);
TASK_PP(16'h80A7,4);
TASK_PP(16'h80A8,4);
TASK_PP(16'h80A9,4);
TASK_PP(16'h80AA,4);
TASK_PP(16'h80AB,4);
TASK_PP(16'h80AC,4);
TASK_PP(16'h80AD,4);
TASK_PP(16'h80AE,4);
TASK_PP(16'h80AF,4);
TASK_PP(16'h80B0,4);
TASK_PP(16'h80B1,4);
TASK_PP(16'h80B2,4);
TASK_PP(16'h80B3,4);
TASK_PP(16'h80B4,4);
TASK_PP(16'h80B5,4);
TASK_PP(16'h80B6,4);
TASK_PP(16'h80B7,4);
TASK_PP(16'h80B8,4);
TASK_PP(16'h80B9,4);
TASK_PP(16'h80BA,4);
TASK_PP(16'h80BB,4);
TASK_PP(16'h80BC,4);
TASK_PP(16'h80BD,4);
TASK_PP(16'h80BE,4);
TASK_PP(16'h80BF,4);
TASK_PP(16'h80C0,4);
TASK_PP(16'h80C1,4);
TASK_PP(16'h80C2,4);
TASK_PP(16'h80C3,4);
TASK_PP(16'h80C4,4);
TASK_PP(16'h80C5,4);
TASK_PP(16'h80C6,4);
TASK_PP(16'h80C7,4);
TASK_PP(16'h80C8,4);
TASK_PP(16'h80C9,4);
TASK_PP(16'h80CA,4);
TASK_PP(16'h80CB,4);
TASK_PP(16'h80CC,4);
TASK_PP(16'h80CD,4);
TASK_PP(16'h80CE,4);
TASK_PP(16'h80CF,4);
TASK_PP(16'h80D0,4);
TASK_PP(16'h80D1,4);
TASK_PP(16'h80D2,4);
TASK_PP(16'h80D3,4);
TASK_PP(16'h80D4,4);
TASK_PP(16'h80D5,4);
TASK_PP(16'h80D6,4);
TASK_PP(16'h80D7,4);
TASK_PP(16'h80D8,4);
TASK_PP(16'h80D9,4);
TASK_PP(16'h80DA,4);
TASK_PP(16'h80DB,4);
TASK_PP(16'h80DC,4);
TASK_PP(16'h80DD,4);
TASK_PP(16'h80DE,4);
TASK_PP(16'h80DF,4);
TASK_PP(16'h80E0,4);
TASK_PP(16'h80E1,4);
TASK_PP(16'h80E2,4);
TASK_PP(16'h80E3,4);
TASK_PP(16'h80E4,4);
TASK_PP(16'h80E5,4);
TASK_PP(16'h80E6,4);
TASK_PP(16'h80E7,4);
TASK_PP(16'h80E8,4);
TASK_PP(16'h80E9,4);
TASK_PP(16'h80EA,4);
TASK_PP(16'h80EB,4);
TASK_PP(16'h80EC,4);
TASK_PP(16'h80ED,4);
TASK_PP(16'h80EE,4);
TASK_PP(16'h80EF,4);
TASK_PP(16'h80F0,4);
TASK_PP(16'h80F1,4);
TASK_PP(16'h80F2,4);
TASK_PP(16'h80F3,4);
TASK_PP(16'h80F4,4);
TASK_PP(16'h80F5,4);
TASK_PP(16'h80F6,4);
TASK_PP(16'h80F7,4);
TASK_PP(16'h80F8,4);
TASK_PP(16'h80F9,4);
TASK_PP(16'h80FA,4);
TASK_PP(16'h80FB,4);
TASK_PP(16'h80FC,4);
TASK_PP(16'h80FD,4);
TASK_PP(16'h80FE,4);
TASK_PP(16'h80FF,4);
TASK_PP(16'h8100,4);
TASK_PP(16'h8101,4);
TASK_PP(16'h8102,4);
TASK_PP(16'h8103,4);
TASK_PP(16'h8104,4);
TASK_PP(16'h8105,4);
TASK_PP(16'h8106,4);
TASK_PP(16'h8107,4);
TASK_PP(16'h8108,4);
TASK_PP(16'h8109,4);
TASK_PP(16'h810A,4);
TASK_PP(16'h810B,4);
TASK_PP(16'h810C,4);
TASK_PP(16'h810D,4);
TASK_PP(16'h810E,4);
TASK_PP(16'h810F,4);
TASK_PP(16'h8110,4);
TASK_PP(16'h8111,4);
TASK_PP(16'h8112,4);
TASK_PP(16'h8113,4);
TASK_PP(16'h8114,4);
TASK_PP(16'h8115,4);
TASK_PP(16'h8116,4);
TASK_PP(16'h8117,4);
TASK_PP(16'h8118,4);
TASK_PP(16'h8119,4);
TASK_PP(16'h811A,4);
TASK_PP(16'h811B,4);
TASK_PP(16'h811C,4);
TASK_PP(16'h811D,4);
TASK_PP(16'h811E,4);
TASK_PP(16'h811F,4);
TASK_PP(16'h8120,4);
TASK_PP(16'h8121,4);
TASK_PP(16'h8122,4);
TASK_PP(16'h8123,4);
TASK_PP(16'h8124,4);
TASK_PP(16'h8125,4);
TASK_PP(16'h8126,4);
TASK_PP(16'h8127,4);
TASK_PP(16'h8128,4);
TASK_PP(16'h8129,4);
TASK_PP(16'h812A,4);
TASK_PP(16'h812B,4);
TASK_PP(16'h812C,4);
TASK_PP(16'h812D,4);
TASK_PP(16'h812E,4);
TASK_PP(16'h812F,4);
TASK_PP(16'h8130,4);
TASK_PP(16'h8131,4);
TASK_PP(16'h8132,4);
TASK_PP(16'h8133,4);
TASK_PP(16'h8134,4);
TASK_PP(16'h8135,4);
TASK_PP(16'h8136,4);
TASK_PP(16'h8137,4);
TASK_PP(16'h8138,4);
TASK_PP(16'h8139,4);
TASK_PP(16'h813A,4);
TASK_PP(16'h813B,4);
TASK_PP(16'h813C,4);
TASK_PP(16'h813D,4);
TASK_PP(16'h813E,4);
TASK_PP(16'h813F,4);
TASK_PP(16'h8140,4);
TASK_PP(16'h8141,4);
TASK_PP(16'h8142,4);
TASK_PP(16'h8143,4);
TASK_PP(16'h8144,4);
TASK_PP(16'h8145,4);
TASK_PP(16'h8146,4);
TASK_PP(16'h8147,4);
TASK_PP(16'h8148,4);
TASK_PP(16'h8149,4);
TASK_PP(16'h814A,4);
TASK_PP(16'h814B,4);
TASK_PP(16'h814C,4);
TASK_PP(16'h814D,4);
TASK_PP(16'h814E,4);
TASK_PP(16'h814F,4);
TASK_PP(16'h8150,4);
TASK_PP(16'h8151,4);
TASK_PP(16'h8152,4);
TASK_PP(16'h8153,4);
TASK_PP(16'h8154,4);
TASK_PP(16'h8155,4);
TASK_PP(16'h8156,4);
TASK_PP(16'h8157,4);
TASK_PP(16'h8158,4);
TASK_PP(16'h8159,4);
TASK_PP(16'h815A,4);
TASK_PP(16'h815B,4);
TASK_PP(16'h815C,4);
TASK_PP(16'h815D,4);
TASK_PP(16'h815E,4);
TASK_PP(16'h815F,4);
TASK_PP(16'h8160,4);
TASK_PP(16'h8161,4);
TASK_PP(16'h8162,4);
TASK_PP(16'h8163,4);
TASK_PP(16'h8164,4);
TASK_PP(16'h8165,4);
TASK_PP(16'h8166,4);
TASK_PP(16'h8167,4);
TASK_PP(16'h8168,4);
TASK_PP(16'h8169,4);
TASK_PP(16'h816A,4);
TASK_PP(16'h816B,4);
TASK_PP(16'h816C,4);
TASK_PP(16'h816D,4);
TASK_PP(16'h816E,4);
TASK_PP(16'h816F,4);
TASK_PP(16'h8170,4);
TASK_PP(16'h8171,4);
TASK_PP(16'h8172,4);
TASK_PP(16'h8173,4);
TASK_PP(16'h8174,4);
TASK_PP(16'h8175,4);
TASK_PP(16'h8176,4);
TASK_PP(16'h8177,4);
TASK_PP(16'h8178,4);
TASK_PP(16'h8179,4);
TASK_PP(16'h817A,4);
TASK_PP(16'h817B,4);
TASK_PP(16'h817C,4);
TASK_PP(16'h817D,4);
TASK_PP(16'h817E,4);
TASK_PP(16'h817F,4);
TASK_PP(16'h8180,4);
TASK_PP(16'h8181,4);
TASK_PP(16'h8182,4);
TASK_PP(16'h8183,4);
TASK_PP(16'h8184,4);
TASK_PP(16'h8185,4);
TASK_PP(16'h8186,4);
TASK_PP(16'h8187,4);
TASK_PP(16'h8188,4);
TASK_PP(16'h8189,4);
TASK_PP(16'h818A,4);
TASK_PP(16'h818B,4);
TASK_PP(16'h818C,4);
TASK_PP(16'h818D,4);
TASK_PP(16'h818E,4);
TASK_PP(16'h818F,4);
TASK_PP(16'h8190,4);
TASK_PP(16'h8191,4);
TASK_PP(16'h8192,4);
TASK_PP(16'h8193,4);
TASK_PP(16'h8194,4);
TASK_PP(16'h8195,4);
TASK_PP(16'h8196,4);
TASK_PP(16'h8197,4);
TASK_PP(16'h8198,4);
TASK_PP(16'h8199,4);
TASK_PP(16'h819A,4);
TASK_PP(16'h819B,4);
TASK_PP(16'h819C,4);
TASK_PP(16'h819D,4);
TASK_PP(16'h819E,4);
TASK_PP(16'h819F,4);
TASK_PP(16'h81A0,4);
TASK_PP(16'h81A1,4);
TASK_PP(16'h81A2,4);
TASK_PP(16'h81A3,4);
TASK_PP(16'h81A4,4);
TASK_PP(16'h81A5,4);
TASK_PP(16'h81A6,4);
TASK_PP(16'h81A7,4);
TASK_PP(16'h81A8,4);
TASK_PP(16'h81A9,4);
TASK_PP(16'h81AA,4);
TASK_PP(16'h81AB,4);
TASK_PP(16'h81AC,4);
TASK_PP(16'h81AD,4);
TASK_PP(16'h81AE,4);
TASK_PP(16'h81AF,4);
TASK_PP(16'h81B0,4);
TASK_PP(16'h81B1,4);
TASK_PP(16'h81B2,4);
TASK_PP(16'h81B3,4);
TASK_PP(16'h81B4,4);
TASK_PP(16'h81B5,4);
TASK_PP(16'h81B6,4);
TASK_PP(16'h81B7,4);
TASK_PP(16'h81B8,4);
TASK_PP(16'h81B9,4);
TASK_PP(16'h81BA,4);
TASK_PP(16'h81BB,4);
TASK_PP(16'h81BC,4);
TASK_PP(16'h81BD,4);
TASK_PP(16'h81BE,4);
TASK_PP(16'h81BF,4);
TASK_PP(16'h81C0,4);
TASK_PP(16'h81C1,4);
TASK_PP(16'h81C2,4);
TASK_PP(16'h81C3,4);
TASK_PP(16'h81C4,4);
TASK_PP(16'h81C5,4);
TASK_PP(16'h81C6,4);
TASK_PP(16'h81C7,4);
TASK_PP(16'h81C8,4);
TASK_PP(16'h81C9,4);
TASK_PP(16'h81CA,4);
TASK_PP(16'h81CB,4);
TASK_PP(16'h81CC,4);
TASK_PP(16'h81CD,4);
TASK_PP(16'h81CE,4);
TASK_PP(16'h81CF,4);
TASK_PP(16'h81D0,4);
TASK_PP(16'h81D1,4);
TASK_PP(16'h81D2,4);
TASK_PP(16'h81D3,4);
TASK_PP(16'h81D4,4);
TASK_PP(16'h81D5,4);
TASK_PP(16'h81D6,4);
TASK_PP(16'h81D7,4);
TASK_PP(16'h81D8,4);
TASK_PP(16'h81D9,4);
TASK_PP(16'h81DA,4);
TASK_PP(16'h81DB,4);
TASK_PP(16'h81DC,4);
TASK_PP(16'h81DD,4);
TASK_PP(16'h81DE,4);
TASK_PP(16'h81DF,4);
TASK_PP(16'h81E0,4);
TASK_PP(16'h81E1,4);
TASK_PP(16'h81E2,4);
TASK_PP(16'h81E3,4);
TASK_PP(16'h81E4,4);
TASK_PP(16'h81E5,4);
TASK_PP(16'h81E6,4);
TASK_PP(16'h81E7,4);
TASK_PP(16'h81E8,4);
TASK_PP(16'h81E9,4);
TASK_PP(16'h81EA,4);
TASK_PP(16'h81EB,4);
TASK_PP(16'h81EC,4);
TASK_PP(16'h81ED,4);
TASK_PP(16'h81EE,4);
TASK_PP(16'h81EF,4);
TASK_PP(16'h81F0,4);
TASK_PP(16'h81F1,4);
TASK_PP(16'h81F2,4);
TASK_PP(16'h81F3,4);
TASK_PP(16'h81F4,4);
TASK_PP(16'h81F5,4);
TASK_PP(16'h81F6,4);
TASK_PP(16'h81F7,4);
TASK_PP(16'h81F8,4);
TASK_PP(16'h81F9,4);
TASK_PP(16'h81FA,4);
TASK_PP(16'h81FB,4);
TASK_PP(16'h81FC,4);
TASK_PP(16'h81FD,4);
TASK_PP(16'h81FE,4);
TASK_PP(16'h81FF,4);
TASK_PP(16'h8200,4);
TASK_PP(16'h8201,4);
TASK_PP(16'h8202,4);
TASK_PP(16'h8203,4);
TASK_PP(16'h8204,4);
TASK_PP(16'h8205,4);
TASK_PP(16'h8206,4);
TASK_PP(16'h8207,4);
TASK_PP(16'h8208,4);
TASK_PP(16'h8209,4);
TASK_PP(16'h820A,4);
TASK_PP(16'h820B,4);
TASK_PP(16'h820C,4);
TASK_PP(16'h820D,4);
TASK_PP(16'h820E,4);
TASK_PP(16'h820F,4);
TASK_PP(16'h8210,4);
TASK_PP(16'h8211,4);
TASK_PP(16'h8212,4);
TASK_PP(16'h8213,4);
TASK_PP(16'h8214,4);
TASK_PP(16'h8215,4);
TASK_PP(16'h8216,4);
TASK_PP(16'h8217,4);
TASK_PP(16'h8218,4);
TASK_PP(16'h8219,4);
TASK_PP(16'h821A,4);
TASK_PP(16'h821B,4);
TASK_PP(16'h821C,4);
TASK_PP(16'h821D,4);
TASK_PP(16'h821E,4);
TASK_PP(16'h821F,4);
TASK_PP(16'h8220,4);
TASK_PP(16'h8221,4);
TASK_PP(16'h8222,4);
TASK_PP(16'h8223,4);
TASK_PP(16'h8224,4);
TASK_PP(16'h8225,4);
TASK_PP(16'h8226,4);
TASK_PP(16'h8227,4);
TASK_PP(16'h8228,4);
TASK_PP(16'h8229,4);
TASK_PP(16'h822A,4);
TASK_PP(16'h822B,4);
TASK_PP(16'h822C,4);
TASK_PP(16'h822D,4);
TASK_PP(16'h822E,4);
TASK_PP(16'h822F,4);
TASK_PP(16'h8230,4);
TASK_PP(16'h8231,4);
TASK_PP(16'h8232,4);
TASK_PP(16'h8233,4);
TASK_PP(16'h8234,4);
TASK_PP(16'h8235,4);
TASK_PP(16'h8236,4);
TASK_PP(16'h8237,4);
TASK_PP(16'h8238,4);
TASK_PP(16'h8239,4);
TASK_PP(16'h823A,4);
TASK_PP(16'h823B,4);
TASK_PP(16'h823C,4);
TASK_PP(16'h823D,4);
TASK_PP(16'h823E,4);
TASK_PP(16'h823F,4);
TASK_PP(16'h8240,4);
TASK_PP(16'h8241,4);
TASK_PP(16'h8242,4);
TASK_PP(16'h8243,4);
TASK_PP(16'h8244,4);
TASK_PP(16'h8245,4);
TASK_PP(16'h8246,4);
TASK_PP(16'h8247,4);
TASK_PP(16'h8248,4);
TASK_PP(16'h8249,4);
TASK_PP(16'h824A,4);
TASK_PP(16'h824B,4);
TASK_PP(16'h824C,4);
TASK_PP(16'h824D,4);
TASK_PP(16'h824E,4);
TASK_PP(16'h824F,4);
TASK_PP(16'h8250,4);
TASK_PP(16'h8251,4);
TASK_PP(16'h8252,4);
TASK_PP(16'h8253,4);
TASK_PP(16'h8254,4);
TASK_PP(16'h8255,4);
TASK_PP(16'h8256,4);
TASK_PP(16'h8257,4);
TASK_PP(16'h8258,4);
TASK_PP(16'h8259,4);
TASK_PP(16'h825A,4);
TASK_PP(16'h825B,4);
TASK_PP(16'h825C,4);
TASK_PP(16'h825D,4);
TASK_PP(16'h825E,4);
TASK_PP(16'h825F,4);
TASK_PP(16'h8260,4);
TASK_PP(16'h8261,4);
TASK_PP(16'h8262,4);
TASK_PP(16'h8263,4);
TASK_PP(16'h8264,4);
TASK_PP(16'h8265,4);
TASK_PP(16'h8266,4);
TASK_PP(16'h8267,4);
TASK_PP(16'h8268,4);
TASK_PP(16'h8269,4);
TASK_PP(16'h826A,4);
TASK_PP(16'h826B,4);
TASK_PP(16'h826C,4);
TASK_PP(16'h826D,4);
TASK_PP(16'h826E,4);
TASK_PP(16'h826F,4);
TASK_PP(16'h8270,4);
TASK_PP(16'h8271,4);
TASK_PP(16'h8272,4);
TASK_PP(16'h8273,4);
TASK_PP(16'h8274,4);
TASK_PP(16'h8275,4);
TASK_PP(16'h8276,4);
TASK_PP(16'h8277,4);
TASK_PP(16'h8278,4);
TASK_PP(16'h8279,4);
TASK_PP(16'h827A,4);
TASK_PP(16'h827B,4);
TASK_PP(16'h827C,4);
TASK_PP(16'h827D,4);
TASK_PP(16'h827E,4);
TASK_PP(16'h827F,4);
TASK_PP(16'h8280,4);
TASK_PP(16'h8281,4);
TASK_PP(16'h8282,4);
TASK_PP(16'h8283,4);
TASK_PP(16'h8284,4);
TASK_PP(16'h8285,4);
TASK_PP(16'h8286,4);
TASK_PP(16'h8287,4);
TASK_PP(16'h8288,4);
TASK_PP(16'h8289,4);
TASK_PP(16'h828A,4);
TASK_PP(16'h828B,4);
TASK_PP(16'h828C,4);
TASK_PP(16'h828D,4);
TASK_PP(16'h828E,4);
TASK_PP(16'h828F,4);
TASK_PP(16'h8290,4);
TASK_PP(16'h8291,4);
TASK_PP(16'h8292,4);
TASK_PP(16'h8293,4);
TASK_PP(16'h8294,4);
TASK_PP(16'h8295,4);
TASK_PP(16'h8296,4);
TASK_PP(16'h8297,4);
TASK_PP(16'h8298,4);
TASK_PP(16'h8299,4);
TASK_PP(16'h829A,4);
TASK_PP(16'h829B,4);
TASK_PP(16'h829C,4);
TASK_PP(16'h829D,4);
TASK_PP(16'h829E,4);
TASK_PP(16'h829F,4);
TASK_PP(16'h82A0,4);
TASK_PP(16'h82A1,4);
TASK_PP(16'h82A2,4);
TASK_PP(16'h82A3,4);
TASK_PP(16'h82A4,4);
TASK_PP(16'h82A5,4);
TASK_PP(16'h82A6,4);
TASK_PP(16'h82A7,4);
TASK_PP(16'h82A8,4);
TASK_PP(16'h82A9,4);
TASK_PP(16'h82AA,4);
TASK_PP(16'h82AB,4);
TASK_PP(16'h82AC,4);
TASK_PP(16'h82AD,4);
TASK_PP(16'h82AE,4);
TASK_PP(16'h82AF,4);
TASK_PP(16'h82B0,4);
TASK_PP(16'h82B1,4);
TASK_PP(16'h82B2,4);
TASK_PP(16'h82B3,4);
TASK_PP(16'h82B4,4);
TASK_PP(16'h82B5,4);
TASK_PP(16'h82B6,4);
TASK_PP(16'h82B7,4);
TASK_PP(16'h82B8,4);
TASK_PP(16'h82B9,4);
TASK_PP(16'h82BA,4);
TASK_PP(16'h82BB,4);
TASK_PP(16'h82BC,4);
TASK_PP(16'h82BD,4);
TASK_PP(16'h82BE,4);
TASK_PP(16'h82BF,4);
TASK_PP(16'h82C0,4);
TASK_PP(16'h82C1,4);
TASK_PP(16'h82C2,4);
TASK_PP(16'h82C3,4);
TASK_PP(16'h82C4,4);
TASK_PP(16'h82C5,4);
TASK_PP(16'h82C6,4);
TASK_PP(16'h82C7,4);
TASK_PP(16'h82C8,4);
TASK_PP(16'h82C9,4);
TASK_PP(16'h82CA,4);
TASK_PP(16'h82CB,4);
TASK_PP(16'h82CC,4);
TASK_PP(16'h82CD,4);
TASK_PP(16'h82CE,4);
TASK_PP(16'h82CF,4);
TASK_PP(16'h82D0,4);
TASK_PP(16'h82D1,4);
TASK_PP(16'h82D2,4);
TASK_PP(16'h82D3,4);
TASK_PP(16'h82D4,4);
TASK_PP(16'h82D5,4);
TASK_PP(16'h82D6,4);
TASK_PP(16'h82D7,4);
TASK_PP(16'h82D8,4);
TASK_PP(16'h82D9,4);
TASK_PP(16'h82DA,4);
TASK_PP(16'h82DB,4);
TASK_PP(16'h82DC,4);
TASK_PP(16'h82DD,4);
TASK_PP(16'h82DE,4);
TASK_PP(16'h82DF,4);
TASK_PP(16'h82E0,4);
TASK_PP(16'h82E1,4);
TASK_PP(16'h82E2,4);
TASK_PP(16'h82E3,4);
TASK_PP(16'h82E4,4);
TASK_PP(16'h82E5,4);
TASK_PP(16'h82E6,4);
TASK_PP(16'h82E7,4);
TASK_PP(16'h82E8,4);
TASK_PP(16'h82E9,4);
TASK_PP(16'h82EA,4);
TASK_PP(16'h82EB,4);
TASK_PP(16'h82EC,4);
TASK_PP(16'h82ED,4);
TASK_PP(16'h82EE,4);
TASK_PP(16'h82EF,4);
TASK_PP(16'h82F0,4);
TASK_PP(16'h82F1,4);
TASK_PP(16'h82F2,4);
TASK_PP(16'h82F3,4);
TASK_PP(16'h82F4,4);
TASK_PP(16'h82F5,4);
TASK_PP(16'h82F6,4);
TASK_PP(16'h82F7,4);
TASK_PP(16'h82F8,4);
TASK_PP(16'h82F9,4);
TASK_PP(16'h82FA,4);
TASK_PP(16'h82FB,4);
TASK_PP(16'h82FC,4);
TASK_PP(16'h82FD,4);
TASK_PP(16'h82FE,4);
TASK_PP(16'h82FF,4);
TASK_PP(16'h8300,4);
TASK_PP(16'h8301,4);
TASK_PP(16'h8302,4);
TASK_PP(16'h8303,4);
TASK_PP(16'h8304,4);
TASK_PP(16'h8305,4);
TASK_PP(16'h8306,4);
TASK_PP(16'h8307,4);
TASK_PP(16'h8308,4);
TASK_PP(16'h8309,4);
TASK_PP(16'h830A,4);
TASK_PP(16'h830B,4);
TASK_PP(16'h830C,4);
TASK_PP(16'h830D,4);
TASK_PP(16'h830E,4);
TASK_PP(16'h830F,4);
TASK_PP(16'h8310,4);
TASK_PP(16'h8311,4);
TASK_PP(16'h8312,4);
TASK_PP(16'h8313,4);
TASK_PP(16'h8314,4);
TASK_PP(16'h8315,4);
TASK_PP(16'h8316,4);
TASK_PP(16'h8317,4);
TASK_PP(16'h8318,4);
TASK_PP(16'h8319,4);
TASK_PP(16'h831A,4);
TASK_PP(16'h831B,4);
TASK_PP(16'h831C,4);
TASK_PP(16'h831D,4);
TASK_PP(16'h831E,4);
TASK_PP(16'h831F,4);
TASK_PP(16'h8320,4);
TASK_PP(16'h8321,4);
TASK_PP(16'h8322,4);
TASK_PP(16'h8323,4);
TASK_PP(16'h8324,4);
TASK_PP(16'h8325,4);
TASK_PP(16'h8326,4);
TASK_PP(16'h8327,4);
TASK_PP(16'h8328,4);
TASK_PP(16'h8329,4);
TASK_PP(16'h832A,4);
TASK_PP(16'h832B,4);
TASK_PP(16'h832C,4);
TASK_PP(16'h832D,4);
TASK_PP(16'h832E,4);
TASK_PP(16'h832F,4);
TASK_PP(16'h8330,4);
TASK_PP(16'h8331,4);
TASK_PP(16'h8332,4);
TASK_PP(16'h8333,4);
TASK_PP(16'h8334,4);
TASK_PP(16'h8335,4);
TASK_PP(16'h8336,4);
TASK_PP(16'h8337,4);
TASK_PP(16'h8338,4);
TASK_PP(16'h8339,4);
TASK_PP(16'h833A,4);
TASK_PP(16'h833B,4);
TASK_PP(16'h833C,4);
TASK_PP(16'h833D,4);
TASK_PP(16'h833E,4);
TASK_PP(16'h833F,4);
TASK_PP(16'h8340,4);
TASK_PP(16'h8341,4);
TASK_PP(16'h8342,4);
TASK_PP(16'h8343,4);
TASK_PP(16'h8344,4);
TASK_PP(16'h8345,4);
TASK_PP(16'h8346,4);
TASK_PP(16'h8347,4);
TASK_PP(16'h8348,4);
TASK_PP(16'h8349,4);
TASK_PP(16'h834A,4);
TASK_PP(16'h834B,4);
TASK_PP(16'h834C,4);
TASK_PP(16'h834D,4);
TASK_PP(16'h834E,4);
TASK_PP(16'h834F,4);
TASK_PP(16'h8350,4);
TASK_PP(16'h8351,4);
TASK_PP(16'h8352,4);
TASK_PP(16'h8353,4);
TASK_PP(16'h8354,4);
TASK_PP(16'h8355,4);
TASK_PP(16'h8356,4);
TASK_PP(16'h8357,4);
TASK_PP(16'h8358,4);
TASK_PP(16'h8359,4);
TASK_PP(16'h835A,4);
TASK_PP(16'h835B,4);
TASK_PP(16'h835C,4);
TASK_PP(16'h835D,4);
TASK_PP(16'h835E,4);
TASK_PP(16'h835F,4);
TASK_PP(16'h8360,4);
TASK_PP(16'h8361,4);
TASK_PP(16'h8362,4);
TASK_PP(16'h8363,4);
TASK_PP(16'h8364,4);
TASK_PP(16'h8365,4);
TASK_PP(16'h8366,4);
TASK_PP(16'h8367,4);
TASK_PP(16'h8368,4);
TASK_PP(16'h8369,4);
TASK_PP(16'h836A,4);
TASK_PP(16'h836B,4);
TASK_PP(16'h836C,4);
TASK_PP(16'h836D,4);
TASK_PP(16'h836E,4);
TASK_PP(16'h836F,4);
TASK_PP(16'h8370,4);
TASK_PP(16'h8371,4);
TASK_PP(16'h8372,4);
TASK_PP(16'h8373,4);
TASK_PP(16'h8374,4);
TASK_PP(16'h8375,4);
TASK_PP(16'h8376,4);
TASK_PP(16'h8377,4);
TASK_PP(16'h8378,4);
TASK_PP(16'h8379,4);
TASK_PP(16'h837A,4);
TASK_PP(16'h837B,4);
TASK_PP(16'h837C,4);
TASK_PP(16'h837D,4);
TASK_PP(16'h837E,4);
TASK_PP(16'h837F,4);
TASK_PP(16'h8380,4);
TASK_PP(16'h8381,4);
TASK_PP(16'h8382,4);
TASK_PP(16'h8383,4);
TASK_PP(16'h8384,4);
TASK_PP(16'h8385,4);
TASK_PP(16'h8386,4);
TASK_PP(16'h8387,4);
TASK_PP(16'h8388,4);
TASK_PP(16'h8389,4);
TASK_PP(16'h838A,4);
TASK_PP(16'h838B,4);
TASK_PP(16'h838C,4);
TASK_PP(16'h838D,4);
TASK_PP(16'h838E,4);
TASK_PP(16'h838F,4);
TASK_PP(16'h8390,4);
TASK_PP(16'h8391,4);
TASK_PP(16'h8392,4);
TASK_PP(16'h8393,4);
TASK_PP(16'h8394,4);
TASK_PP(16'h8395,4);
TASK_PP(16'h8396,4);
TASK_PP(16'h8397,4);
TASK_PP(16'h8398,4);
TASK_PP(16'h8399,4);
TASK_PP(16'h839A,4);
TASK_PP(16'h839B,4);
TASK_PP(16'h839C,4);
TASK_PP(16'h839D,4);
TASK_PP(16'h839E,4);
TASK_PP(16'h839F,4);
TASK_PP(16'h83A0,4);
TASK_PP(16'h83A1,4);
TASK_PP(16'h83A2,4);
TASK_PP(16'h83A3,4);
TASK_PP(16'h83A4,4);
TASK_PP(16'h83A5,4);
TASK_PP(16'h83A6,4);
TASK_PP(16'h83A7,4);
TASK_PP(16'h83A8,4);
TASK_PP(16'h83A9,4);
TASK_PP(16'h83AA,4);
TASK_PP(16'h83AB,4);
TASK_PP(16'h83AC,4);
TASK_PP(16'h83AD,4);
TASK_PP(16'h83AE,4);
TASK_PP(16'h83AF,4);
TASK_PP(16'h83B0,4);
TASK_PP(16'h83B1,4);
TASK_PP(16'h83B2,4);
TASK_PP(16'h83B3,4);
TASK_PP(16'h83B4,4);
TASK_PP(16'h83B5,4);
TASK_PP(16'h83B6,4);
TASK_PP(16'h83B7,4);
TASK_PP(16'h83B8,4);
TASK_PP(16'h83B9,4);
TASK_PP(16'h83BA,4);
TASK_PP(16'h83BB,4);
TASK_PP(16'h83BC,4);
TASK_PP(16'h83BD,4);
TASK_PP(16'h83BE,4);
TASK_PP(16'h83BF,4);
TASK_PP(16'h83C0,4);
TASK_PP(16'h83C1,4);
TASK_PP(16'h83C2,4);
TASK_PP(16'h83C3,4);
TASK_PP(16'h83C4,4);
TASK_PP(16'h83C5,4);
TASK_PP(16'h83C6,4);
TASK_PP(16'h83C7,4);
TASK_PP(16'h83C8,4);
TASK_PP(16'h83C9,4);
TASK_PP(16'h83CA,4);
TASK_PP(16'h83CB,4);
TASK_PP(16'h83CC,4);
TASK_PP(16'h83CD,4);
TASK_PP(16'h83CE,4);
TASK_PP(16'h83CF,4);
TASK_PP(16'h83D0,4);
TASK_PP(16'h83D1,4);
TASK_PP(16'h83D2,4);
TASK_PP(16'h83D3,4);
TASK_PP(16'h83D4,4);
TASK_PP(16'h83D5,4);
TASK_PP(16'h83D6,4);
TASK_PP(16'h83D7,4);
TASK_PP(16'h83D8,4);
TASK_PP(16'h83D9,4);
TASK_PP(16'h83DA,4);
TASK_PP(16'h83DB,4);
TASK_PP(16'h83DC,4);
TASK_PP(16'h83DD,4);
TASK_PP(16'h83DE,4);
TASK_PP(16'h83DF,4);
TASK_PP(16'h83E0,4);
TASK_PP(16'h83E1,4);
TASK_PP(16'h83E2,4);
TASK_PP(16'h83E3,4);
TASK_PP(16'h83E4,4);
TASK_PP(16'h83E5,4);
TASK_PP(16'h83E6,4);
TASK_PP(16'h83E7,4);
TASK_PP(16'h83E8,4);
TASK_PP(16'h83E9,4);
TASK_PP(16'h83EA,4);
TASK_PP(16'h83EB,4);
TASK_PP(16'h83EC,4);
TASK_PP(16'h83ED,4);
TASK_PP(16'h83EE,4);
TASK_PP(16'h83EF,4);
TASK_PP(16'h83F0,4);
TASK_PP(16'h83F1,4);
TASK_PP(16'h83F2,4);
TASK_PP(16'h83F3,4);
TASK_PP(16'h83F4,4);
TASK_PP(16'h83F5,4);
TASK_PP(16'h83F6,4);
TASK_PP(16'h83F7,4);
TASK_PP(16'h83F8,4);
TASK_PP(16'h83F9,4);
TASK_PP(16'h83FA,4);
TASK_PP(16'h83FB,4);
TASK_PP(16'h83FC,4);
TASK_PP(16'h83FD,4);
TASK_PP(16'h83FE,4);
TASK_PP(16'h83FF,4);
TASK_PP(16'h8400,4);
TASK_PP(16'h8401,4);
TASK_PP(16'h8402,4);
TASK_PP(16'h8403,4);
TASK_PP(16'h8404,4);
TASK_PP(16'h8405,4);
TASK_PP(16'h8406,4);
TASK_PP(16'h8407,4);
TASK_PP(16'h8408,4);
TASK_PP(16'h8409,4);
TASK_PP(16'h840A,4);
TASK_PP(16'h840B,4);
TASK_PP(16'h840C,4);
TASK_PP(16'h840D,4);
TASK_PP(16'h840E,4);
TASK_PP(16'h840F,4);
TASK_PP(16'h8410,4);
TASK_PP(16'h8411,4);
TASK_PP(16'h8412,4);
TASK_PP(16'h8413,4);
TASK_PP(16'h8414,4);
TASK_PP(16'h8415,4);
TASK_PP(16'h8416,4);
TASK_PP(16'h8417,4);
TASK_PP(16'h8418,4);
TASK_PP(16'h8419,4);
TASK_PP(16'h841A,4);
TASK_PP(16'h841B,4);
TASK_PP(16'h841C,4);
TASK_PP(16'h841D,4);
TASK_PP(16'h841E,4);
TASK_PP(16'h841F,4);
TASK_PP(16'h8420,4);
TASK_PP(16'h8421,4);
TASK_PP(16'h8422,4);
TASK_PP(16'h8423,4);
TASK_PP(16'h8424,4);
TASK_PP(16'h8425,4);
TASK_PP(16'h8426,4);
TASK_PP(16'h8427,4);
TASK_PP(16'h8428,4);
TASK_PP(16'h8429,4);
TASK_PP(16'h842A,4);
TASK_PP(16'h842B,4);
TASK_PP(16'h842C,4);
TASK_PP(16'h842D,4);
TASK_PP(16'h842E,4);
TASK_PP(16'h842F,4);
TASK_PP(16'h8430,4);
TASK_PP(16'h8431,4);
TASK_PP(16'h8432,4);
TASK_PP(16'h8433,4);
TASK_PP(16'h8434,4);
TASK_PP(16'h8435,4);
TASK_PP(16'h8436,4);
TASK_PP(16'h8437,4);
TASK_PP(16'h8438,4);
TASK_PP(16'h8439,4);
TASK_PP(16'h843A,4);
TASK_PP(16'h843B,4);
TASK_PP(16'h843C,4);
TASK_PP(16'h843D,4);
TASK_PP(16'h843E,4);
TASK_PP(16'h843F,4);
TASK_PP(16'h8440,4);
TASK_PP(16'h8441,4);
TASK_PP(16'h8442,4);
TASK_PP(16'h8443,4);
TASK_PP(16'h8444,4);
TASK_PP(16'h8445,4);
TASK_PP(16'h8446,4);
TASK_PP(16'h8447,4);
TASK_PP(16'h8448,4);
TASK_PP(16'h8449,4);
TASK_PP(16'h844A,4);
TASK_PP(16'h844B,4);
TASK_PP(16'h844C,4);
TASK_PP(16'h844D,4);
TASK_PP(16'h844E,4);
TASK_PP(16'h844F,4);
TASK_PP(16'h8450,4);
TASK_PP(16'h8451,4);
TASK_PP(16'h8452,4);
TASK_PP(16'h8453,4);
TASK_PP(16'h8454,4);
TASK_PP(16'h8455,4);
TASK_PP(16'h8456,4);
TASK_PP(16'h8457,4);
TASK_PP(16'h8458,4);
TASK_PP(16'h8459,4);
TASK_PP(16'h845A,4);
TASK_PP(16'h845B,4);
TASK_PP(16'h845C,4);
TASK_PP(16'h845D,4);
TASK_PP(16'h845E,4);
TASK_PP(16'h845F,4);
TASK_PP(16'h8460,4);
TASK_PP(16'h8461,4);
TASK_PP(16'h8462,4);
TASK_PP(16'h8463,4);
TASK_PP(16'h8464,4);
TASK_PP(16'h8465,4);
TASK_PP(16'h8466,4);
TASK_PP(16'h8467,4);
TASK_PP(16'h8468,4);
TASK_PP(16'h8469,4);
TASK_PP(16'h846A,4);
TASK_PP(16'h846B,4);
TASK_PP(16'h846C,4);
TASK_PP(16'h846D,4);
TASK_PP(16'h846E,4);
TASK_PP(16'h846F,4);
TASK_PP(16'h8470,4);
TASK_PP(16'h8471,4);
TASK_PP(16'h8472,4);
TASK_PP(16'h8473,4);
TASK_PP(16'h8474,4);
TASK_PP(16'h8475,4);
TASK_PP(16'h8476,4);
TASK_PP(16'h8477,4);
TASK_PP(16'h8478,4);
TASK_PP(16'h8479,4);
TASK_PP(16'h847A,4);
TASK_PP(16'h847B,4);
TASK_PP(16'h847C,4);
TASK_PP(16'h847D,4);
TASK_PP(16'h847E,4);
TASK_PP(16'h847F,4);
TASK_PP(16'h8480,4);
TASK_PP(16'h8481,4);
TASK_PP(16'h8482,4);
TASK_PP(16'h8483,4);
TASK_PP(16'h8484,4);
TASK_PP(16'h8485,4);
TASK_PP(16'h8486,4);
TASK_PP(16'h8487,4);
TASK_PP(16'h8488,4);
TASK_PP(16'h8489,4);
TASK_PP(16'h848A,4);
TASK_PP(16'h848B,4);
TASK_PP(16'h848C,4);
TASK_PP(16'h848D,4);
TASK_PP(16'h848E,4);
TASK_PP(16'h848F,4);
TASK_PP(16'h8490,4);
TASK_PP(16'h8491,4);
TASK_PP(16'h8492,4);
TASK_PP(16'h8493,4);
TASK_PP(16'h8494,4);
TASK_PP(16'h8495,4);
TASK_PP(16'h8496,4);
TASK_PP(16'h8497,4);
TASK_PP(16'h8498,4);
TASK_PP(16'h8499,4);
TASK_PP(16'h849A,4);
TASK_PP(16'h849B,4);
TASK_PP(16'h849C,4);
TASK_PP(16'h849D,4);
TASK_PP(16'h849E,4);
TASK_PP(16'h849F,4);
TASK_PP(16'h84A0,4);
TASK_PP(16'h84A1,4);
TASK_PP(16'h84A2,4);
TASK_PP(16'h84A3,4);
TASK_PP(16'h84A4,4);
TASK_PP(16'h84A5,4);
TASK_PP(16'h84A6,4);
TASK_PP(16'h84A7,4);
TASK_PP(16'h84A8,4);
TASK_PP(16'h84A9,4);
TASK_PP(16'h84AA,4);
TASK_PP(16'h84AB,4);
TASK_PP(16'h84AC,4);
TASK_PP(16'h84AD,4);
TASK_PP(16'h84AE,4);
TASK_PP(16'h84AF,4);
TASK_PP(16'h84B0,4);
TASK_PP(16'h84B1,4);
TASK_PP(16'h84B2,4);
TASK_PP(16'h84B3,4);
TASK_PP(16'h84B4,4);
TASK_PP(16'h84B5,4);
TASK_PP(16'h84B6,4);
TASK_PP(16'h84B7,4);
TASK_PP(16'h84B8,4);
TASK_PP(16'h84B9,4);
TASK_PP(16'h84BA,4);
TASK_PP(16'h84BB,4);
TASK_PP(16'h84BC,4);
TASK_PP(16'h84BD,4);
TASK_PP(16'h84BE,4);
TASK_PP(16'h84BF,4);
TASK_PP(16'h84C0,4);
TASK_PP(16'h84C1,4);
TASK_PP(16'h84C2,4);
TASK_PP(16'h84C3,4);
TASK_PP(16'h84C4,4);
TASK_PP(16'h84C5,4);
TASK_PP(16'h84C6,4);
TASK_PP(16'h84C7,4);
TASK_PP(16'h84C8,4);
TASK_PP(16'h84C9,4);
TASK_PP(16'h84CA,4);
TASK_PP(16'h84CB,4);
TASK_PP(16'h84CC,4);
TASK_PP(16'h84CD,4);
TASK_PP(16'h84CE,4);
TASK_PP(16'h84CF,4);
TASK_PP(16'h84D0,4);
TASK_PP(16'h84D1,4);
TASK_PP(16'h84D2,4);
TASK_PP(16'h84D3,4);
TASK_PP(16'h84D4,4);
TASK_PP(16'h84D5,4);
TASK_PP(16'h84D6,4);
TASK_PP(16'h84D7,4);
TASK_PP(16'h84D8,4);
TASK_PP(16'h84D9,4);
TASK_PP(16'h84DA,4);
TASK_PP(16'h84DB,4);
TASK_PP(16'h84DC,4);
TASK_PP(16'h84DD,4);
TASK_PP(16'h84DE,4);
TASK_PP(16'h84DF,4);
TASK_PP(16'h84E0,4);
TASK_PP(16'h84E1,4);
TASK_PP(16'h84E2,4);
TASK_PP(16'h84E3,4);
TASK_PP(16'h84E4,4);
TASK_PP(16'h84E5,4);
TASK_PP(16'h84E6,4);
TASK_PP(16'h84E7,4);
TASK_PP(16'h84E8,4);
TASK_PP(16'h84E9,4);
TASK_PP(16'h84EA,4);
TASK_PP(16'h84EB,4);
TASK_PP(16'h84EC,4);
TASK_PP(16'h84ED,4);
TASK_PP(16'h84EE,4);
TASK_PP(16'h84EF,4);
TASK_PP(16'h84F0,4);
TASK_PP(16'h84F1,4);
TASK_PP(16'h84F2,4);
TASK_PP(16'h84F3,4);
TASK_PP(16'h84F4,4);
TASK_PP(16'h84F5,4);
TASK_PP(16'h84F6,4);
TASK_PP(16'h84F7,4);
TASK_PP(16'h84F8,4);
TASK_PP(16'h84F9,4);
TASK_PP(16'h84FA,4);
TASK_PP(16'h84FB,4);
TASK_PP(16'h84FC,4);
TASK_PP(16'h84FD,4);
TASK_PP(16'h84FE,4);
TASK_PP(16'h84FF,4);
TASK_PP(16'h8500,4);
TASK_PP(16'h8501,4);
TASK_PP(16'h8502,4);
TASK_PP(16'h8503,4);
TASK_PP(16'h8504,4);
TASK_PP(16'h8505,4);
TASK_PP(16'h8506,4);
TASK_PP(16'h8507,4);
TASK_PP(16'h8508,4);
TASK_PP(16'h8509,4);
TASK_PP(16'h850A,4);
TASK_PP(16'h850B,4);
TASK_PP(16'h850C,4);
TASK_PP(16'h850D,4);
TASK_PP(16'h850E,4);
TASK_PP(16'h850F,4);
TASK_PP(16'h8510,4);
TASK_PP(16'h8511,4);
TASK_PP(16'h8512,4);
TASK_PP(16'h8513,4);
TASK_PP(16'h8514,4);
TASK_PP(16'h8515,4);
TASK_PP(16'h8516,4);
TASK_PP(16'h8517,4);
TASK_PP(16'h8518,4);
TASK_PP(16'h8519,4);
TASK_PP(16'h851A,4);
TASK_PP(16'h851B,4);
TASK_PP(16'h851C,4);
TASK_PP(16'h851D,4);
TASK_PP(16'h851E,4);
TASK_PP(16'h851F,4);
TASK_PP(16'h8520,4);
TASK_PP(16'h8521,4);
TASK_PP(16'h8522,4);
TASK_PP(16'h8523,4);
TASK_PP(16'h8524,4);
TASK_PP(16'h8525,4);
TASK_PP(16'h8526,4);
TASK_PP(16'h8527,4);
TASK_PP(16'h8528,4);
TASK_PP(16'h8529,4);
TASK_PP(16'h852A,4);
TASK_PP(16'h852B,4);
TASK_PP(16'h852C,4);
TASK_PP(16'h852D,4);
TASK_PP(16'h852E,4);
TASK_PP(16'h852F,4);
TASK_PP(16'h8530,4);
TASK_PP(16'h8531,4);
TASK_PP(16'h8532,4);
TASK_PP(16'h8533,4);
TASK_PP(16'h8534,4);
TASK_PP(16'h8535,4);
TASK_PP(16'h8536,4);
TASK_PP(16'h8537,4);
TASK_PP(16'h8538,4);
TASK_PP(16'h8539,4);
TASK_PP(16'h853A,4);
TASK_PP(16'h853B,4);
TASK_PP(16'h853C,4);
TASK_PP(16'h853D,4);
TASK_PP(16'h853E,4);
TASK_PP(16'h853F,4);
TASK_PP(16'h8540,4);
TASK_PP(16'h8541,4);
TASK_PP(16'h8542,4);
TASK_PP(16'h8543,4);
TASK_PP(16'h8544,4);
TASK_PP(16'h8545,4);
TASK_PP(16'h8546,4);
TASK_PP(16'h8547,4);
TASK_PP(16'h8548,4);
TASK_PP(16'h8549,4);
TASK_PP(16'h854A,4);
TASK_PP(16'h854B,4);
TASK_PP(16'h854C,4);
TASK_PP(16'h854D,4);
TASK_PP(16'h854E,4);
TASK_PP(16'h854F,4);
TASK_PP(16'h8550,4);
TASK_PP(16'h8551,4);
TASK_PP(16'h8552,4);
TASK_PP(16'h8553,4);
TASK_PP(16'h8554,4);
TASK_PP(16'h8555,4);
TASK_PP(16'h8556,4);
TASK_PP(16'h8557,4);
TASK_PP(16'h8558,4);
TASK_PP(16'h8559,4);
TASK_PP(16'h855A,4);
TASK_PP(16'h855B,4);
TASK_PP(16'h855C,4);
TASK_PP(16'h855D,4);
TASK_PP(16'h855E,4);
TASK_PP(16'h855F,4);
TASK_PP(16'h8560,4);
TASK_PP(16'h8561,4);
TASK_PP(16'h8562,4);
TASK_PP(16'h8563,4);
TASK_PP(16'h8564,4);
TASK_PP(16'h8565,4);
TASK_PP(16'h8566,4);
TASK_PP(16'h8567,4);
TASK_PP(16'h8568,4);
TASK_PP(16'h8569,4);
TASK_PP(16'h856A,4);
TASK_PP(16'h856B,4);
TASK_PP(16'h856C,4);
TASK_PP(16'h856D,4);
TASK_PP(16'h856E,4);
TASK_PP(16'h856F,4);
TASK_PP(16'h8570,4);
TASK_PP(16'h8571,4);
TASK_PP(16'h8572,4);
TASK_PP(16'h8573,4);
TASK_PP(16'h8574,4);
TASK_PP(16'h8575,4);
TASK_PP(16'h8576,4);
TASK_PP(16'h8577,4);
TASK_PP(16'h8578,4);
TASK_PP(16'h8579,4);
TASK_PP(16'h857A,4);
TASK_PP(16'h857B,4);
TASK_PP(16'h857C,4);
TASK_PP(16'h857D,4);
TASK_PP(16'h857E,4);
TASK_PP(16'h857F,4);
TASK_PP(16'h8580,4);
TASK_PP(16'h8581,4);
TASK_PP(16'h8582,4);
TASK_PP(16'h8583,4);
TASK_PP(16'h8584,4);
TASK_PP(16'h8585,4);
TASK_PP(16'h8586,4);
TASK_PP(16'h8587,4);
TASK_PP(16'h8588,4);
TASK_PP(16'h8589,4);
TASK_PP(16'h858A,4);
TASK_PP(16'h858B,4);
TASK_PP(16'h858C,4);
TASK_PP(16'h858D,4);
TASK_PP(16'h858E,4);
TASK_PP(16'h858F,4);
TASK_PP(16'h8590,4);
TASK_PP(16'h8591,4);
TASK_PP(16'h8592,4);
TASK_PP(16'h8593,4);
TASK_PP(16'h8594,4);
TASK_PP(16'h8595,4);
TASK_PP(16'h8596,4);
TASK_PP(16'h8597,4);
TASK_PP(16'h8598,4);
TASK_PP(16'h8599,4);
TASK_PP(16'h859A,4);
TASK_PP(16'h859B,4);
TASK_PP(16'h859C,4);
TASK_PP(16'h859D,4);
TASK_PP(16'h859E,4);
TASK_PP(16'h859F,4);
TASK_PP(16'h85A0,4);
TASK_PP(16'h85A1,4);
TASK_PP(16'h85A2,4);
TASK_PP(16'h85A3,4);
TASK_PP(16'h85A4,4);
TASK_PP(16'h85A5,4);
TASK_PP(16'h85A6,4);
TASK_PP(16'h85A7,4);
TASK_PP(16'h85A8,4);
TASK_PP(16'h85A9,4);
TASK_PP(16'h85AA,4);
TASK_PP(16'h85AB,4);
TASK_PP(16'h85AC,4);
TASK_PP(16'h85AD,4);
TASK_PP(16'h85AE,4);
TASK_PP(16'h85AF,4);
TASK_PP(16'h85B0,4);
TASK_PP(16'h85B1,4);
TASK_PP(16'h85B2,4);
TASK_PP(16'h85B3,4);
TASK_PP(16'h85B4,4);
TASK_PP(16'h85B5,4);
TASK_PP(16'h85B6,4);
TASK_PP(16'h85B7,4);
TASK_PP(16'h85B8,4);
TASK_PP(16'h85B9,4);
TASK_PP(16'h85BA,4);
TASK_PP(16'h85BB,4);
TASK_PP(16'h85BC,4);
TASK_PP(16'h85BD,4);
TASK_PP(16'h85BE,4);
TASK_PP(16'h85BF,4);
TASK_PP(16'h85C0,4);
TASK_PP(16'h85C1,4);
TASK_PP(16'h85C2,4);
TASK_PP(16'h85C3,4);
TASK_PP(16'h85C4,4);
TASK_PP(16'h85C5,4);
TASK_PP(16'h85C6,4);
TASK_PP(16'h85C7,4);
TASK_PP(16'h85C8,4);
TASK_PP(16'h85C9,4);
TASK_PP(16'h85CA,4);
TASK_PP(16'h85CB,4);
TASK_PP(16'h85CC,4);
TASK_PP(16'h85CD,4);
TASK_PP(16'h85CE,4);
TASK_PP(16'h85CF,4);
TASK_PP(16'h85D0,4);
TASK_PP(16'h85D1,4);
TASK_PP(16'h85D2,4);
TASK_PP(16'h85D3,4);
TASK_PP(16'h85D4,4);
TASK_PP(16'h85D5,4);
TASK_PP(16'h85D6,4);
TASK_PP(16'h85D7,4);
TASK_PP(16'h85D8,4);
TASK_PP(16'h85D9,4);
TASK_PP(16'h85DA,4);
TASK_PP(16'h85DB,4);
TASK_PP(16'h85DC,4);
TASK_PP(16'h85DD,4);
TASK_PP(16'h85DE,4);
TASK_PP(16'h85DF,4);
TASK_PP(16'h85E0,4);
TASK_PP(16'h85E1,4);
TASK_PP(16'h85E2,4);
TASK_PP(16'h85E3,4);
TASK_PP(16'h85E4,4);
TASK_PP(16'h85E5,4);
TASK_PP(16'h85E6,4);
TASK_PP(16'h85E7,4);
TASK_PP(16'h85E8,4);
TASK_PP(16'h85E9,4);
TASK_PP(16'h85EA,4);
TASK_PP(16'h85EB,4);
TASK_PP(16'h85EC,4);
TASK_PP(16'h85ED,4);
TASK_PP(16'h85EE,4);
TASK_PP(16'h85EF,4);
TASK_PP(16'h85F0,4);
TASK_PP(16'h85F1,4);
TASK_PP(16'h85F2,4);
TASK_PP(16'h85F3,4);
TASK_PP(16'h85F4,4);
TASK_PP(16'h85F5,4);
TASK_PP(16'h85F6,4);
TASK_PP(16'h85F7,4);
TASK_PP(16'h85F8,4);
TASK_PP(16'h85F9,4);
TASK_PP(16'h85FA,4);
TASK_PP(16'h85FB,4);
TASK_PP(16'h85FC,4);
TASK_PP(16'h85FD,4);
TASK_PP(16'h85FE,4);
TASK_PP(16'h85FF,4);
TASK_PP(16'h8600,4);
TASK_PP(16'h8601,4);
TASK_PP(16'h8602,4);
TASK_PP(16'h8603,4);
TASK_PP(16'h8604,4);
TASK_PP(16'h8605,4);
TASK_PP(16'h8606,4);
TASK_PP(16'h8607,4);
TASK_PP(16'h8608,4);
TASK_PP(16'h8609,4);
TASK_PP(16'h860A,4);
TASK_PP(16'h860B,4);
TASK_PP(16'h860C,4);
TASK_PP(16'h860D,4);
TASK_PP(16'h860E,4);
TASK_PP(16'h860F,4);
TASK_PP(16'h8610,4);
TASK_PP(16'h8611,4);
TASK_PP(16'h8612,4);
TASK_PP(16'h8613,4);
TASK_PP(16'h8614,4);
TASK_PP(16'h8615,4);
TASK_PP(16'h8616,4);
TASK_PP(16'h8617,4);
TASK_PP(16'h8618,4);
TASK_PP(16'h8619,4);
TASK_PP(16'h861A,4);
TASK_PP(16'h861B,4);
TASK_PP(16'h861C,4);
TASK_PP(16'h861D,4);
TASK_PP(16'h861E,4);
TASK_PP(16'h861F,4);
TASK_PP(16'h8620,4);
TASK_PP(16'h8621,4);
TASK_PP(16'h8622,4);
TASK_PP(16'h8623,4);
TASK_PP(16'h8624,4);
TASK_PP(16'h8625,4);
TASK_PP(16'h8626,4);
TASK_PP(16'h8627,4);
TASK_PP(16'h8628,4);
TASK_PP(16'h8629,4);
TASK_PP(16'h862A,4);
TASK_PP(16'h862B,4);
TASK_PP(16'h862C,4);
TASK_PP(16'h862D,4);
TASK_PP(16'h862E,4);
TASK_PP(16'h862F,4);
TASK_PP(16'h8630,4);
TASK_PP(16'h8631,4);
TASK_PP(16'h8632,4);
TASK_PP(16'h8633,4);
TASK_PP(16'h8634,4);
TASK_PP(16'h8635,4);
TASK_PP(16'h8636,4);
TASK_PP(16'h8637,4);
TASK_PP(16'h8638,4);
TASK_PP(16'h8639,4);
TASK_PP(16'h863A,4);
TASK_PP(16'h863B,4);
TASK_PP(16'h863C,4);
TASK_PP(16'h863D,4);
TASK_PP(16'h863E,4);
TASK_PP(16'h863F,4);
TASK_PP(16'h8640,4);
TASK_PP(16'h8641,4);
TASK_PP(16'h8642,4);
TASK_PP(16'h8643,4);
TASK_PP(16'h8644,4);
TASK_PP(16'h8645,4);
TASK_PP(16'h8646,4);
TASK_PP(16'h8647,4);
TASK_PP(16'h8648,4);
TASK_PP(16'h8649,4);
TASK_PP(16'h864A,4);
TASK_PP(16'h864B,4);
TASK_PP(16'h864C,4);
TASK_PP(16'h864D,4);
TASK_PP(16'h864E,4);
TASK_PP(16'h864F,4);
TASK_PP(16'h8650,4);
TASK_PP(16'h8651,4);
TASK_PP(16'h8652,4);
TASK_PP(16'h8653,4);
TASK_PP(16'h8654,4);
TASK_PP(16'h8655,4);
TASK_PP(16'h8656,4);
TASK_PP(16'h8657,4);
TASK_PP(16'h8658,4);
TASK_PP(16'h8659,4);
TASK_PP(16'h865A,4);
TASK_PP(16'h865B,4);
TASK_PP(16'h865C,4);
TASK_PP(16'h865D,4);
TASK_PP(16'h865E,4);
TASK_PP(16'h865F,4);
TASK_PP(16'h8660,4);
TASK_PP(16'h8661,4);
TASK_PP(16'h8662,4);
TASK_PP(16'h8663,4);
TASK_PP(16'h8664,4);
TASK_PP(16'h8665,4);
TASK_PP(16'h8666,4);
TASK_PP(16'h8667,4);
TASK_PP(16'h8668,4);
TASK_PP(16'h8669,4);
TASK_PP(16'h866A,4);
TASK_PP(16'h866B,4);
TASK_PP(16'h866C,4);
TASK_PP(16'h866D,4);
TASK_PP(16'h866E,4);
TASK_PP(16'h866F,4);
TASK_PP(16'h8670,4);
TASK_PP(16'h8671,4);
TASK_PP(16'h8672,4);
TASK_PP(16'h8673,4);
TASK_PP(16'h8674,4);
TASK_PP(16'h8675,4);
TASK_PP(16'h8676,4);
TASK_PP(16'h8677,4);
TASK_PP(16'h8678,4);
TASK_PP(16'h8679,4);
TASK_PP(16'h867A,4);
TASK_PP(16'h867B,4);
TASK_PP(16'h867C,4);
TASK_PP(16'h867D,4);
TASK_PP(16'h867E,4);
TASK_PP(16'h867F,4);
TASK_PP(16'h8680,4);
TASK_PP(16'h8681,4);
TASK_PP(16'h8682,4);
TASK_PP(16'h8683,4);
TASK_PP(16'h8684,4);
TASK_PP(16'h8685,4);
TASK_PP(16'h8686,4);
TASK_PP(16'h8687,4);
TASK_PP(16'h8688,4);
TASK_PP(16'h8689,4);
TASK_PP(16'h868A,4);
TASK_PP(16'h868B,4);
TASK_PP(16'h868C,4);
TASK_PP(16'h868D,4);
TASK_PP(16'h868E,4);
TASK_PP(16'h868F,4);
TASK_PP(16'h8690,4);
TASK_PP(16'h8691,4);
TASK_PP(16'h8692,4);
TASK_PP(16'h8693,4);
TASK_PP(16'h8694,4);
TASK_PP(16'h8695,4);
TASK_PP(16'h8696,4);
TASK_PP(16'h8697,4);
TASK_PP(16'h8698,4);
TASK_PP(16'h8699,4);
TASK_PP(16'h869A,4);
TASK_PP(16'h869B,4);
TASK_PP(16'h869C,4);
TASK_PP(16'h869D,4);
TASK_PP(16'h869E,4);
TASK_PP(16'h869F,4);
TASK_PP(16'h86A0,4);
TASK_PP(16'h86A1,4);
TASK_PP(16'h86A2,4);
TASK_PP(16'h86A3,4);
TASK_PP(16'h86A4,4);
TASK_PP(16'h86A5,4);
TASK_PP(16'h86A6,4);
TASK_PP(16'h86A7,4);
TASK_PP(16'h86A8,4);
TASK_PP(16'h86A9,4);
TASK_PP(16'h86AA,4);
TASK_PP(16'h86AB,4);
TASK_PP(16'h86AC,4);
TASK_PP(16'h86AD,4);
TASK_PP(16'h86AE,4);
TASK_PP(16'h86AF,4);
TASK_PP(16'h86B0,4);
TASK_PP(16'h86B1,4);
TASK_PP(16'h86B2,4);
TASK_PP(16'h86B3,4);
TASK_PP(16'h86B4,4);
TASK_PP(16'h86B5,4);
TASK_PP(16'h86B6,4);
TASK_PP(16'h86B7,4);
TASK_PP(16'h86B8,4);
TASK_PP(16'h86B9,4);
TASK_PP(16'h86BA,4);
TASK_PP(16'h86BB,4);
TASK_PP(16'h86BC,4);
TASK_PP(16'h86BD,4);
TASK_PP(16'h86BE,4);
TASK_PP(16'h86BF,4);
TASK_PP(16'h86C0,4);
TASK_PP(16'h86C1,4);
TASK_PP(16'h86C2,4);
TASK_PP(16'h86C3,4);
TASK_PP(16'h86C4,4);
TASK_PP(16'h86C5,4);
TASK_PP(16'h86C6,4);
TASK_PP(16'h86C7,4);
TASK_PP(16'h86C8,4);
TASK_PP(16'h86C9,4);
TASK_PP(16'h86CA,4);
TASK_PP(16'h86CB,4);
TASK_PP(16'h86CC,4);
TASK_PP(16'h86CD,4);
TASK_PP(16'h86CE,4);
TASK_PP(16'h86CF,4);
TASK_PP(16'h86D0,4);
TASK_PP(16'h86D1,4);
TASK_PP(16'h86D2,4);
TASK_PP(16'h86D3,4);
TASK_PP(16'h86D4,4);
TASK_PP(16'h86D5,4);
TASK_PP(16'h86D6,4);
TASK_PP(16'h86D7,4);
TASK_PP(16'h86D8,4);
TASK_PP(16'h86D9,4);
TASK_PP(16'h86DA,4);
TASK_PP(16'h86DB,4);
TASK_PP(16'h86DC,4);
TASK_PP(16'h86DD,4);
TASK_PP(16'h86DE,4);
TASK_PP(16'h86DF,4);
TASK_PP(16'h86E0,4);
TASK_PP(16'h86E1,4);
TASK_PP(16'h86E2,4);
TASK_PP(16'h86E3,4);
TASK_PP(16'h86E4,4);
TASK_PP(16'h86E5,4);
TASK_PP(16'h86E6,4);
TASK_PP(16'h86E7,4);
TASK_PP(16'h86E8,4);
TASK_PP(16'h86E9,4);
TASK_PP(16'h86EA,4);
TASK_PP(16'h86EB,4);
TASK_PP(16'h86EC,4);
TASK_PP(16'h86ED,4);
TASK_PP(16'h86EE,4);
TASK_PP(16'h86EF,4);
TASK_PP(16'h86F0,4);
TASK_PP(16'h86F1,4);
TASK_PP(16'h86F2,4);
TASK_PP(16'h86F3,4);
TASK_PP(16'h86F4,4);
TASK_PP(16'h86F5,4);
TASK_PP(16'h86F6,4);
TASK_PP(16'h86F7,4);
TASK_PP(16'h86F8,4);
TASK_PP(16'h86F9,4);
TASK_PP(16'h86FA,4);
TASK_PP(16'h86FB,4);
TASK_PP(16'h86FC,4);
TASK_PP(16'h86FD,4);
TASK_PP(16'h86FE,4);
TASK_PP(16'h86FF,4);
TASK_PP(16'h8700,4);
TASK_PP(16'h8701,4);
TASK_PP(16'h8702,4);
TASK_PP(16'h8703,4);
TASK_PP(16'h8704,4);
TASK_PP(16'h8705,4);
TASK_PP(16'h8706,4);
TASK_PP(16'h8707,4);
TASK_PP(16'h8708,4);
TASK_PP(16'h8709,4);
TASK_PP(16'h870A,4);
TASK_PP(16'h870B,4);
TASK_PP(16'h870C,4);
TASK_PP(16'h870D,4);
TASK_PP(16'h870E,4);
TASK_PP(16'h870F,4);
TASK_PP(16'h8710,4);
TASK_PP(16'h8711,4);
TASK_PP(16'h8712,4);
TASK_PP(16'h8713,4);
TASK_PP(16'h8714,4);
TASK_PP(16'h8715,4);
TASK_PP(16'h8716,4);
TASK_PP(16'h8717,4);
TASK_PP(16'h8718,4);
TASK_PP(16'h8719,4);
TASK_PP(16'h871A,4);
TASK_PP(16'h871B,4);
TASK_PP(16'h871C,4);
TASK_PP(16'h871D,4);
TASK_PP(16'h871E,4);
TASK_PP(16'h871F,4);
TASK_PP(16'h8720,4);
TASK_PP(16'h8721,4);
TASK_PP(16'h8722,4);
TASK_PP(16'h8723,4);
TASK_PP(16'h8724,4);
TASK_PP(16'h8725,4);
TASK_PP(16'h8726,4);
TASK_PP(16'h8727,4);
TASK_PP(16'h8728,4);
TASK_PP(16'h8729,4);
TASK_PP(16'h872A,4);
TASK_PP(16'h872B,4);
TASK_PP(16'h872C,4);
TASK_PP(16'h872D,4);
TASK_PP(16'h872E,4);
TASK_PP(16'h872F,4);
TASK_PP(16'h8730,4);
TASK_PP(16'h8731,4);
TASK_PP(16'h8732,4);
TASK_PP(16'h8733,4);
TASK_PP(16'h8734,4);
TASK_PP(16'h8735,4);
TASK_PP(16'h8736,4);
TASK_PP(16'h8737,4);
TASK_PP(16'h8738,4);
TASK_PP(16'h8739,4);
TASK_PP(16'h873A,4);
TASK_PP(16'h873B,4);
TASK_PP(16'h873C,4);
TASK_PP(16'h873D,4);
TASK_PP(16'h873E,4);
TASK_PP(16'h873F,4);
TASK_PP(16'h8740,4);
TASK_PP(16'h8741,4);
TASK_PP(16'h8742,4);
TASK_PP(16'h8743,4);
TASK_PP(16'h8744,4);
TASK_PP(16'h8745,4);
TASK_PP(16'h8746,4);
TASK_PP(16'h8747,4);
TASK_PP(16'h8748,4);
TASK_PP(16'h8749,4);
TASK_PP(16'h874A,4);
TASK_PP(16'h874B,4);
TASK_PP(16'h874C,4);
TASK_PP(16'h874D,4);
TASK_PP(16'h874E,4);
TASK_PP(16'h874F,4);
TASK_PP(16'h8750,4);
TASK_PP(16'h8751,4);
TASK_PP(16'h8752,4);
TASK_PP(16'h8753,4);
TASK_PP(16'h8754,4);
TASK_PP(16'h8755,4);
TASK_PP(16'h8756,4);
TASK_PP(16'h8757,4);
TASK_PP(16'h8758,4);
TASK_PP(16'h8759,4);
TASK_PP(16'h875A,4);
TASK_PP(16'h875B,4);
TASK_PP(16'h875C,4);
TASK_PP(16'h875D,4);
TASK_PP(16'h875E,4);
TASK_PP(16'h875F,4);
TASK_PP(16'h8760,4);
TASK_PP(16'h8761,4);
TASK_PP(16'h8762,4);
TASK_PP(16'h8763,4);
TASK_PP(16'h8764,4);
TASK_PP(16'h8765,4);
TASK_PP(16'h8766,4);
TASK_PP(16'h8767,4);
TASK_PP(16'h8768,4);
TASK_PP(16'h8769,4);
TASK_PP(16'h876A,4);
TASK_PP(16'h876B,4);
TASK_PP(16'h876C,4);
TASK_PP(16'h876D,4);
TASK_PP(16'h876E,4);
TASK_PP(16'h876F,4);
TASK_PP(16'h8770,4);
TASK_PP(16'h8771,4);
TASK_PP(16'h8772,4);
TASK_PP(16'h8773,4);
TASK_PP(16'h8774,4);
TASK_PP(16'h8775,4);
TASK_PP(16'h8776,4);
TASK_PP(16'h8777,4);
TASK_PP(16'h8778,4);
TASK_PP(16'h8779,4);
TASK_PP(16'h877A,4);
TASK_PP(16'h877B,4);
TASK_PP(16'h877C,4);
TASK_PP(16'h877D,4);
TASK_PP(16'h877E,4);
TASK_PP(16'h877F,4);
TASK_PP(16'h8780,4);
TASK_PP(16'h8781,4);
TASK_PP(16'h8782,4);
TASK_PP(16'h8783,4);
TASK_PP(16'h8784,4);
TASK_PP(16'h8785,4);
TASK_PP(16'h8786,4);
TASK_PP(16'h8787,4);
TASK_PP(16'h8788,4);
TASK_PP(16'h8789,4);
TASK_PP(16'h878A,4);
TASK_PP(16'h878B,4);
TASK_PP(16'h878C,4);
TASK_PP(16'h878D,4);
TASK_PP(16'h878E,4);
TASK_PP(16'h878F,4);
TASK_PP(16'h8790,4);
TASK_PP(16'h8791,4);
TASK_PP(16'h8792,4);
TASK_PP(16'h8793,4);
TASK_PP(16'h8794,4);
TASK_PP(16'h8795,4);
TASK_PP(16'h8796,4);
TASK_PP(16'h8797,4);
TASK_PP(16'h8798,4);
TASK_PP(16'h8799,4);
TASK_PP(16'h879A,4);
TASK_PP(16'h879B,4);
TASK_PP(16'h879C,4);
TASK_PP(16'h879D,4);
TASK_PP(16'h879E,4);
TASK_PP(16'h879F,4);
TASK_PP(16'h87A0,4);
TASK_PP(16'h87A1,4);
TASK_PP(16'h87A2,4);
TASK_PP(16'h87A3,4);
TASK_PP(16'h87A4,4);
TASK_PP(16'h87A5,4);
TASK_PP(16'h87A6,4);
TASK_PP(16'h87A7,4);
TASK_PP(16'h87A8,4);
TASK_PP(16'h87A9,4);
TASK_PP(16'h87AA,4);
TASK_PP(16'h87AB,4);
TASK_PP(16'h87AC,4);
TASK_PP(16'h87AD,4);
TASK_PP(16'h87AE,4);
TASK_PP(16'h87AF,4);
TASK_PP(16'h87B0,4);
TASK_PP(16'h87B1,4);
TASK_PP(16'h87B2,4);
TASK_PP(16'h87B3,4);
TASK_PP(16'h87B4,4);
TASK_PP(16'h87B5,4);
TASK_PP(16'h87B6,4);
TASK_PP(16'h87B7,4);
TASK_PP(16'h87B8,4);
TASK_PP(16'h87B9,4);
TASK_PP(16'h87BA,4);
TASK_PP(16'h87BB,4);
TASK_PP(16'h87BC,4);
TASK_PP(16'h87BD,4);
TASK_PP(16'h87BE,4);
TASK_PP(16'h87BF,4);
TASK_PP(16'h87C0,4);
TASK_PP(16'h87C1,4);
TASK_PP(16'h87C2,4);
TASK_PP(16'h87C3,4);
TASK_PP(16'h87C4,4);
TASK_PP(16'h87C5,4);
TASK_PP(16'h87C6,4);
TASK_PP(16'h87C7,4);
TASK_PP(16'h87C8,4);
TASK_PP(16'h87C9,4);
TASK_PP(16'h87CA,4);
TASK_PP(16'h87CB,4);
TASK_PP(16'h87CC,4);
TASK_PP(16'h87CD,4);
TASK_PP(16'h87CE,4);
TASK_PP(16'h87CF,4);
TASK_PP(16'h87D0,4);
TASK_PP(16'h87D1,4);
TASK_PP(16'h87D2,4);
TASK_PP(16'h87D3,4);
TASK_PP(16'h87D4,4);
TASK_PP(16'h87D5,4);
TASK_PP(16'h87D6,4);
TASK_PP(16'h87D7,4);
TASK_PP(16'h87D8,4);
TASK_PP(16'h87D9,4);
TASK_PP(16'h87DA,4);
TASK_PP(16'h87DB,4);
TASK_PP(16'h87DC,4);
TASK_PP(16'h87DD,4);
TASK_PP(16'h87DE,4);
TASK_PP(16'h87DF,4);
TASK_PP(16'h87E0,4);
TASK_PP(16'h87E1,4);
TASK_PP(16'h87E2,4);
TASK_PP(16'h87E3,4);
TASK_PP(16'h87E4,4);
TASK_PP(16'h87E5,4);
TASK_PP(16'h87E6,4);
TASK_PP(16'h87E7,4);
TASK_PP(16'h87E8,4);
TASK_PP(16'h87E9,4);
TASK_PP(16'h87EA,4);
TASK_PP(16'h87EB,4);
TASK_PP(16'h87EC,4);
TASK_PP(16'h87ED,4);
TASK_PP(16'h87EE,4);
TASK_PP(16'h87EF,4);
TASK_PP(16'h87F0,4);
TASK_PP(16'h87F1,4);
TASK_PP(16'h87F2,4);
TASK_PP(16'h87F3,4);
TASK_PP(16'h87F4,4);
TASK_PP(16'h87F5,4);
TASK_PP(16'h87F6,4);
TASK_PP(16'h87F7,4);
TASK_PP(16'h87F8,4);
TASK_PP(16'h87F9,4);
TASK_PP(16'h87FA,4);
TASK_PP(16'h87FB,4);
TASK_PP(16'h87FC,4);
TASK_PP(16'h87FD,4);
TASK_PP(16'h87FE,4);
TASK_PP(16'h87FF,4);
TASK_PP(16'h8800,4);
TASK_PP(16'h8801,4);
TASK_PP(16'h8802,4);
TASK_PP(16'h8803,4);
TASK_PP(16'h8804,4);
TASK_PP(16'h8805,4);
TASK_PP(16'h8806,4);
TASK_PP(16'h8807,4);
TASK_PP(16'h8808,4);
TASK_PP(16'h8809,4);
TASK_PP(16'h880A,4);
TASK_PP(16'h880B,4);
TASK_PP(16'h880C,4);
TASK_PP(16'h880D,4);
TASK_PP(16'h880E,4);
TASK_PP(16'h880F,4);
TASK_PP(16'h8810,4);
TASK_PP(16'h8811,4);
TASK_PP(16'h8812,4);
TASK_PP(16'h8813,4);
TASK_PP(16'h8814,4);
TASK_PP(16'h8815,4);
TASK_PP(16'h8816,4);
TASK_PP(16'h8817,4);
TASK_PP(16'h8818,4);
TASK_PP(16'h8819,4);
TASK_PP(16'h881A,4);
TASK_PP(16'h881B,4);
TASK_PP(16'h881C,4);
TASK_PP(16'h881D,4);
TASK_PP(16'h881E,4);
TASK_PP(16'h881F,4);
TASK_PP(16'h8820,4);
TASK_PP(16'h8821,4);
TASK_PP(16'h8822,4);
TASK_PP(16'h8823,4);
TASK_PP(16'h8824,4);
TASK_PP(16'h8825,4);
TASK_PP(16'h8826,4);
TASK_PP(16'h8827,4);
TASK_PP(16'h8828,4);
TASK_PP(16'h8829,4);
TASK_PP(16'h882A,4);
TASK_PP(16'h882B,4);
TASK_PP(16'h882C,4);
TASK_PP(16'h882D,4);
TASK_PP(16'h882E,4);
TASK_PP(16'h882F,4);
TASK_PP(16'h8830,4);
TASK_PP(16'h8831,4);
TASK_PP(16'h8832,4);
TASK_PP(16'h8833,4);
TASK_PP(16'h8834,4);
TASK_PP(16'h8835,4);
TASK_PP(16'h8836,4);
TASK_PP(16'h8837,4);
TASK_PP(16'h8838,4);
TASK_PP(16'h8839,4);
TASK_PP(16'h883A,4);
TASK_PP(16'h883B,4);
TASK_PP(16'h883C,4);
TASK_PP(16'h883D,4);
TASK_PP(16'h883E,4);
TASK_PP(16'h883F,4);
TASK_PP(16'h8840,4);
TASK_PP(16'h8841,4);
TASK_PP(16'h8842,4);
TASK_PP(16'h8843,4);
TASK_PP(16'h8844,4);
TASK_PP(16'h8845,4);
TASK_PP(16'h8846,4);
TASK_PP(16'h8847,4);
TASK_PP(16'h8848,4);
TASK_PP(16'h8849,4);
TASK_PP(16'h884A,4);
TASK_PP(16'h884B,4);
TASK_PP(16'h884C,4);
TASK_PP(16'h884D,4);
TASK_PP(16'h884E,4);
TASK_PP(16'h884F,4);
TASK_PP(16'h8850,4);
TASK_PP(16'h8851,4);
TASK_PP(16'h8852,4);
TASK_PP(16'h8853,4);
TASK_PP(16'h8854,4);
TASK_PP(16'h8855,4);
TASK_PP(16'h8856,4);
TASK_PP(16'h8857,4);
TASK_PP(16'h8858,4);
TASK_PP(16'h8859,4);
TASK_PP(16'h885A,4);
TASK_PP(16'h885B,4);
TASK_PP(16'h885C,4);
TASK_PP(16'h885D,4);
TASK_PP(16'h885E,4);
TASK_PP(16'h885F,4);
TASK_PP(16'h8860,4);
TASK_PP(16'h8861,4);
TASK_PP(16'h8862,4);
TASK_PP(16'h8863,4);
TASK_PP(16'h8864,4);
TASK_PP(16'h8865,4);
TASK_PP(16'h8866,4);
TASK_PP(16'h8867,4);
TASK_PP(16'h8868,4);
TASK_PP(16'h8869,4);
TASK_PP(16'h886A,4);
TASK_PP(16'h886B,4);
TASK_PP(16'h886C,4);
TASK_PP(16'h886D,4);
TASK_PP(16'h886E,4);
TASK_PP(16'h886F,4);
TASK_PP(16'h8870,4);
TASK_PP(16'h8871,4);
TASK_PP(16'h8872,4);
TASK_PP(16'h8873,4);
TASK_PP(16'h8874,4);
TASK_PP(16'h8875,4);
TASK_PP(16'h8876,4);
TASK_PP(16'h8877,4);
TASK_PP(16'h8878,4);
TASK_PP(16'h8879,4);
TASK_PP(16'h887A,4);
TASK_PP(16'h887B,4);
TASK_PP(16'h887C,4);
TASK_PP(16'h887D,4);
TASK_PP(16'h887E,4);
TASK_PP(16'h887F,4);
TASK_PP(16'h8880,4);
TASK_PP(16'h8881,4);
TASK_PP(16'h8882,4);
TASK_PP(16'h8883,4);
TASK_PP(16'h8884,4);
TASK_PP(16'h8885,4);
TASK_PP(16'h8886,4);
TASK_PP(16'h8887,4);
TASK_PP(16'h8888,4);
TASK_PP(16'h8889,4);
TASK_PP(16'h888A,4);
TASK_PP(16'h888B,4);
TASK_PP(16'h888C,4);
TASK_PP(16'h888D,4);
TASK_PP(16'h888E,4);
TASK_PP(16'h888F,4);
TASK_PP(16'h8890,4);
TASK_PP(16'h8891,4);
TASK_PP(16'h8892,4);
TASK_PP(16'h8893,4);
TASK_PP(16'h8894,4);
TASK_PP(16'h8895,4);
TASK_PP(16'h8896,4);
TASK_PP(16'h8897,4);
TASK_PP(16'h8898,4);
TASK_PP(16'h8899,4);
TASK_PP(16'h889A,4);
TASK_PP(16'h889B,4);
TASK_PP(16'h889C,4);
TASK_PP(16'h889D,4);
TASK_PP(16'h889E,4);
TASK_PP(16'h889F,4);
TASK_PP(16'h88A0,4);
TASK_PP(16'h88A1,4);
TASK_PP(16'h88A2,4);
TASK_PP(16'h88A3,4);
TASK_PP(16'h88A4,4);
TASK_PP(16'h88A5,4);
TASK_PP(16'h88A6,4);
TASK_PP(16'h88A7,4);
TASK_PP(16'h88A8,4);
TASK_PP(16'h88A9,4);
TASK_PP(16'h88AA,4);
TASK_PP(16'h88AB,4);
TASK_PP(16'h88AC,4);
TASK_PP(16'h88AD,4);
TASK_PP(16'h88AE,4);
TASK_PP(16'h88AF,4);
TASK_PP(16'h88B0,4);
TASK_PP(16'h88B1,4);
TASK_PP(16'h88B2,4);
TASK_PP(16'h88B3,4);
TASK_PP(16'h88B4,4);
TASK_PP(16'h88B5,4);
TASK_PP(16'h88B6,4);
TASK_PP(16'h88B7,4);
TASK_PP(16'h88B8,4);
TASK_PP(16'h88B9,4);
TASK_PP(16'h88BA,4);
TASK_PP(16'h88BB,4);
TASK_PP(16'h88BC,4);
TASK_PP(16'h88BD,4);
TASK_PP(16'h88BE,4);
TASK_PP(16'h88BF,4);
TASK_PP(16'h88C0,4);
TASK_PP(16'h88C1,4);
TASK_PP(16'h88C2,4);
TASK_PP(16'h88C3,4);
TASK_PP(16'h88C4,4);
TASK_PP(16'h88C5,4);
TASK_PP(16'h88C6,4);
TASK_PP(16'h88C7,4);
TASK_PP(16'h88C8,4);
TASK_PP(16'h88C9,4);
TASK_PP(16'h88CA,4);
TASK_PP(16'h88CB,4);
TASK_PP(16'h88CC,4);
TASK_PP(16'h88CD,4);
TASK_PP(16'h88CE,4);
TASK_PP(16'h88CF,4);
TASK_PP(16'h88D0,4);
TASK_PP(16'h88D1,4);
TASK_PP(16'h88D2,4);
TASK_PP(16'h88D3,4);
TASK_PP(16'h88D4,4);
TASK_PP(16'h88D5,4);
TASK_PP(16'h88D6,4);
TASK_PP(16'h88D7,4);
TASK_PP(16'h88D8,4);
TASK_PP(16'h88D9,4);
TASK_PP(16'h88DA,4);
TASK_PP(16'h88DB,4);
TASK_PP(16'h88DC,4);
TASK_PP(16'h88DD,4);
TASK_PP(16'h88DE,4);
TASK_PP(16'h88DF,4);
TASK_PP(16'h88E0,4);
TASK_PP(16'h88E1,4);
TASK_PP(16'h88E2,4);
TASK_PP(16'h88E3,4);
TASK_PP(16'h88E4,4);
TASK_PP(16'h88E5,4);
TASK_PP(16'h88E6,4);
TASK_PP(16'h88E7,4);
TASK_PP(16'h88E8,4);
TASK_PP(16'h88E9,4);
TASK_PP(16'h88EA,4);
TASK_PP(16'h88EB,4);
TASK_PP(16'h88EC,4);
TASK_PP(16'h88ED,4);
TASK_PP(16'h88EE,4);
TASK_PP(16'h88EF,4);
TASK_PP(16'h88F0,4);
TASK_PP(16'h88F1,4);
TASK_PP(16'h88F2,4);
TASK_PP(16'h88F3,4);
TASK_PP(16'h88F4,4);
TASK_PP(16'h88F5,4);
TASK_PP(16'h88F6,4);
TASK_PP(16'h88F7,4);
TASK_PP(16'h88F8,4);
TASK_PP(16'h88F9,4);
TASK_PP(16'h88FA,4);
TASK_PP(16'h88FB,4);
TASK_PP(16'h88FC,4);
TASK_PP(16'h88FD,4);
TASK_PP(16'h88FE,4);
TASK_PP(16'h88FF,4);
TASK_PP(16'h8900,4);
TASK_PP(16'h8901,4);
TASK_PP(16'h8902,4);
TASK_PP(16'h8903,4);
TASK_PP(16'h8904,4);
TASK_PP(16'h8905,4);
TASK_PP(16'h8906,4);
TASK_PP(16'h8907,4);
TASK_PP(16'h8908,4);
TASK_PP(16'h8909,4);
TASK_PP(16'h890A,4);
TASK_PP(16'h890B,4);
TASK_PP(16'h890C,4);
TASK_PP(16'h890D,4);
TASK_PP(16'h890E,4);
TASK_PP(16'h890F,4);
TASK_PP(16'h8910,4);
TASK_PP(16'h8911,4);
TASK_PP(16'h8912,4);
TASK_PP(16'h8913,4);
TASK_PP(16'h8914,4);
TASK_PP(16'h8915,4);
TASK_PP(16'h8916,4);
TASK_PP(16'h8917,4);
TASK_PP(16'h8918,4);
TASK_PP(16'h8919,4);
TASK_PP(16'h891A,4);
TASK_PP(16'h891B,4);
TASK_PP(16'h891C,4);
TASK_PP(16'h891D,4);
TASK_PP(16'h891E,4);
TASK_PP(16'h891F,4);
TASK_PP(16'h8920,4);
TASK_PP(16'h8921,4);
TASK_PP(16'h8922,4);
TASK_PP(16'h8923,4);
TASK_PP(16'h8924,4);
TASK_PP(16'h8925,4);
TASK_PP(16'h8926,4);
TASK_PP(16'h8927,4);
TASK_PP(16'h8928,4);
TASK_PP(16'h8929,4);
TASK_PP(16'h892A,4);
TASK_PP(16'h892B,4);
TASK_PP(16'h892C,4);
TASK_PP(16'h892D,4);
TASK_PP(16'h892E,4);
TASK_PP(16'h892F,4);
TASK_PP(16'h8930,4);
TASK_PP(16'h8931,4);
TASK_PP(16'h8932,4);
TASK_PP(16'h8933,4);
TASK_PP(16'h8934,4);
TASK_PP(16'h8935,4);
TASK_PP(16'h8936,4);
TASK_PP(16'h8937,4);
TASK_PP(16'h8938,4);
TASK_PP(16'h8939,4);
TASK_PP(16'h893A,4);
TASK_PP(16'h893B,4);
TASK_PP(16'h893C,4);
TASK_PP(16'h893D,4);
TASK_PP(16'h893E,4);
TASK_PP(16'h893F,4);
TASK_PP(16'h8940,4);
TASK_PP(16'h8941,4);
TASK_PP(16'h8942,4);
TASK_PP(16'h8943,4);
TASK_PP(16'h8944,4);
TASK_PP(16'h8945,4);
TASK_PP(16'h8946,4);
TASK_PP(16'h8947,4);
TASK_PP(16'h8948,4);
TASK_PP(16'h8949,4);
TASK_PP(16'h894A,4);
TASK_PP(16'h894B,4);
TASK_PP(16'h894C,4);
TASK_PP(16'h894D,4);
TASK_PP(16'h894E,4);
TASK_PP(16'h894F,4);
TASK_PP(16'h8950,4);
TASK_PP(16'h8951,4);
TASK_PP(16'h8952,4);
TASK_PP(16'h8953,4);
TASK_PP(16'h8954,4);
TASK_PP(16'h8955,4);
TASK_PP(16'h8956,4);
TASK_PP(16'h8957,4);
TASK_PP(16'h8958,4);
TASK_PP(16'h8959,4);
TASK_PP(16'h895A,4);
TASK_PP(16'h895B,4);
TASK_PP(16'h895C,4);
TASK_PP(16'h895D,4);
TASK_PP(16'h895E,4);
TASK_PP(16'h895F,4);
TASK_PP(16'h8960,4);
TASK_PP(16'h8961,4);
TASK_PP(16'h8962,4);
TASK_PP(16'h8963,4);
TASK_PP(16'h8964,4);
TASK_PP(16'h8965,4);
TASK_PP(16'h8966,4);
TASK_PP(16'h8967,4);
TASK_PP(16'h8968,4);
TASK_PP(16'h8969,4);
TASK_PP(16'h896A,4);
TASK_PP(16'h896B,4);
TASK_PP(16'h896C,4);
TASK_PP(16'h896D,4);
TASK_PP(16'h896E,4);
TASK_PP(16'h896F,4);
TASK_PP(16'h8970,4);
TASK_PP(16'h8971,4);
TASK_PP(16'h8972,4);
TASK_PP(16'h8973,4);
TASK_PP(16'h8974,4);
TASK_PP(16'h8975,4);
TASK_PP(16'h8976,4);
TASK_PP(16'h8977,4);
TASK_PP(16'h8978,4);
TASK_PP(16'h8979,4);
TASK_PP(16'h897A,4);
TASK_PP(16'h897B,4);
TASK_PP(16'h897C,4);
TASK_PP(16'h897D,4);
TASK_PP(16'h897E,4);
TASK_PP(16'h897F,4);
TASK_PP(16'h8980,4);
TASK_PP(16'h8981,4);
TASK_PP(16'h8982,4);
TASK_PP(16'h8983,4);
TASK_PP(16'h8984,4);
TASK_PP(16'h8985,4);
TASK_PP(16'h8986,4);
TASK_PP(16'h8987,4);
TASK_PP(16'h8988,4);
TASK_PP(16'h8989,4);
TASK_PP(16'h898A,4);
TASK_PP(16'h898B,4);
TASK_PP(16'h898C,4);
TASK_PP(16'h898D,4);
TASK_PP(16'h898E,4);
TASK_PP(16'h898F,4);
TASK_PP(16'h8990,4);
TASK_PP(16'h8991,4);
TASK_PP(16'h8992,4);
TASK_PP(16'h8993,4);
TASK_PP(16'h8994,4);
TASK_PP(16'h8995,4);
TASK_PP(16'h8996,4);
TASK_PP(16'h8997,4);
TASK_PP(16'h8998,4);
TASK_PP(16'h8999,4);
TASK_PP(16'h899A,4);
TASK_PP(16'h899B,4);
TASK_PP(16'h899C,4);
TASK_PP(16'h899D,4);
TASK_PP(16'h899E,4);
TASK_PP(16'h899F,4);
TASK_PP(16'h89A0,4);
TASK_PP(16'h89A1,4);
TASK_PP(16'h89A2,4);
TASK_PP(16'h89A3,4);
TASK_PP(16'h89A4,4);
TASK_PP(16'h89A5,4);
TASK_PP(16'h89A6,4);
TASK_PP(16'h89A7,4);
TASK_PP(16'h89A8,4);
TASK_PP(16'h89A9,4);
TASK_PP(16'h89AA,4);
TASK_PP(16'h89AB,4);
TASK_PP(16'h89AC,4);
TASK_PP(16'h89AD,4);
TASK_PP(16'h89AE,4);
TASK_PP(16'h89AF,4);
TASK_PP(16'h89B0,4);
TASK_PP(16'h89B1,4);
TASK_PP(16'h89B2,4);
TASK_PP(16'h89B3,4);
TASK_PP(16'h89B4,4);
TASK_PP(16'h89B5,4);
TASK_PP(16'h89B6,4);
TASK_PP(16'h89B7,4);
TASK_PP(16'h89B8,4);
TASK_PP(16'h89B9,4);
TASK_PP(16'h89BA,4);
TASK_PP(16'h89BB,4);
TASK_PP(16'h89BC,4);
TASK_PP(16'h89BD,4);
TASK_PP(16'h89BE,4);
TASK_PP(16'h89BF,4);
TASK_PP(16'h89C0,4);
TASK_PP(16'h89C1,4);
TASK_PP(16'h89C2,4);
TASK_PP(16'h89C3,4);
TASK_PP(16'h89C4,4);
TASK_PP(16'h89C5,4);
TASK_PP(16'h89C6,4);
TASK_PP(16'h89C7,4);
TASK_PP(16'h89C8,4);
TASK_PP(16'h89C9,4);
TASK_PP(16'h89CA,4);
TASK_PP(16'h89CB,4);
TASK_PP(16'h89CC,4);
TASK_PP(16'h89CD,4);
TASK_PP(16'h89CE,4);
TASK_PP(16'h89CF,4);
TASK_PP(16'h89D0,4);
TASK_PP(16'h89D1,4);
TASK_PP(16'h89D2,4);
TASK_PP(16'h89D3,4);
TASK_PP(16'h89D4,4);
TASK_PP(16'h89D5,4);
TASK_PP(16'h89D6,4);
TASK_PP(16'h89D7,4);
TASK_PP(16'h89D8,4);
TASK_PP(16'h89D9,4);
TASK_PP(16'h89DA,4);
TASK_PP(16'h89DB,4);
TASK_PP(16'h89DC,4);
TASK_PP(16'h89DD,4);
TASK_PP(16'h89DE,4);
TASK_PP(16'h89DF,4);
TASK_PP(16'h89E0,4);
TASK_PP(16'h89E1,4);
TASK_PP(16'h89E2,4);
TASK_PP(16'h89E3,4);
TASK_PP(16'h89E4,4);
TASK_PP(16'h89E5,4);
TASK_PP(16'h89E6,4);
TASK_PP(16'h89E7,4);
TASK_PP(16'h89E8,4);
TASK_PP(16'h89E9,4);
TASK_PP(16'h89EA,4);
TASK_PP(16'h89EB,4);
TASK_PP(16'h89EC,4);
TASK_PP(16'h89ED,4);
TASK_PP(16'h89EE,4);
TASK_PP(16'h89EF,4);
TASK_PP(16'h89F0,4);
TASK_PP(16'h89F1,4);
TASK_PP(16'h89F2,4);
TASK_PP(16'h89F3,4);
TASK_PP(16'h89F4,4);
TASK_PP(16'h89F5,4);
TASK_PP(16'h89F6,4);
TASK_PP(16'h89F7,4);
TASK_PP(16'h89F8,4);
TASK_PP(16'h89F9,4);
TASK_PP(16'h89FA,4);
TASK_PP(16'h89FB,4);
TASK_PP(16'h89FC,4);
TASK_PP(16'h89FD,4);
TASK_PP(16'h89FE,4);
TASK_PP(16'h89FF,4);
TASK_PP(16'h8A00,4);
TASK_PP(16'h8A01,4);
TASK_PP(16'h8A02,4);
TASK_PP(16'h8A03,4);
TASK_PP(16'h8A04,4);
TASK_PP(16'h8A05,4);
TASK_PP(16'h8A06,4);
TASK_PP(16'h8A07,4);
TASK_PP(16'h8A08,4);
TASK_PP(16'h8A09,4);
TASK_PP(16'h8A0A,4);
TASK_PP(16'h8A0B,4);
TASK_PP(16'h8A0C,4);
TASK_PP(16'h8A0D,4);
TASK_PP(16'h8A0E,4);
TASK_PP(16'h8A0F,4);
TASK_PP(16'h8A10,4);
TASK_PP(16'h8A11,4);
TASK_PP(16'h8A12,4);
TASK_PP(16'h8A13,4);
TASK_PP(16'h8A14,4);
TASK_PP(16'h8A15,4);
TASK_PP(16'h8A16,4);
TASK_PP(16'h8A17,4);
TASK_PP(16'h8A18,4);
TASK_PP(16'h8A19,4);
TASK_PP(16'h8A1A,4);
TASK_PP(16'h8A1B,4);
TASK_PP(16'h8A1C,4);
TASK_PP(16'h8A1D,4);
TASK_PP(16'h8A1E,4);
TASK_PP(16'h8A1F,4);
TASK_PP(16'h8A20,4);
TASK_PP(16'h8A21,4);
TASK_PP(16'h8A22,4);
TASK_PP(16'h8A23,4);
TASK_PP(16'h8A24,4);
TASK_PP(16'h8A25,4);
TASK_PP(16'h8A26,4);
TASK_PP(16'h8A27,4);
TASK_PP(16'h8A28,4);
TASK_PP(16'h8A29,4);
TASK_PP(16'h8A2A,4);
TASK_PP(16'h8A2B,4);
TASK_PP(16'h8A2C,4);
TASK_PP(16'h8A2D,4);
TASK_PP(16'h8A2E,4);
TASK_PP(16'h8A2F,4);
TASK_PP(16'h8A30,4);
TASK_PP(16'h8A31,4);
TASK_PP(16'h8A32,4);
TASK_PP(16'h8A33,4);
TASK_PP(16'h8A34,4);
TASK_PP(16'h8A35,4);
TASK_PP(16'h8A36,4);
TASK_PP(16'h8A37,4);
TASK_PP(16'h8A38,4);
TASK_PP(16'h8A39,4);
TASK_PP(16'h8A3A,4);
TASK_PP(16'h8A3B,4);
TASK_PP(16'h8A3C,4);
TASK_PP(16'h8A3D,4);
TASK_PP(16'h8A3E,4);
TASK_PP(16'h8A3F,4);
TASK_PP(16'h8A40,4);
TASK_PP(16'h8A41,4);
TASK_PP(16'h8A42,4);
TASK_PP(16'h8A43,4);
TASK_PP(16'h8A44,4);
TASK_PP(16'h8A45,4);
TASK_PP(16'h8A46,4);
TASK_PP(16'h8A47,4);
TASK_PP(16'h8A48,4);
TASK_PP(16'h8A49,4);
TASK_PP(16'h8A4A,4);
TASK_PP(16'h8A4B,4);
TASK_PP(16'h8A4C,4);
TASK_PP(16'h8A4D,4);
TASK_PP(16'h8A4E,4);
TASK_PP(16'h8A4F,4);
TASK_PP(16'h8A50,4);
TASK_PP(16'h8A51,4);
TASK_PP(16'h8A52,4);
TASK_PP(16'h8A53,4);
TASK_PP(16'h8A54,4);
TASK_PP(16'h8A55,4);
TASK_PP(16'h8A56,4);
TASK_PP(16'h8A57,4);
TASK_PP(16'h8A58,4);
TASK_PP(16'h8A59,4);
TASK_PP(16'h8A5A,4);
TASK_PP(16'h8A5B,4);
TASK_PP(16'h8A5C,4);
TASK_PP(16'h8A5D,4);
TASK_PP(16'h8A5E,4);
TASK_PP(16'h8A5F,4);
TASK_PP(16'h8A60,4);
TASK_PP(16'h8A61,4);
TASK_PP(16'h8A62,4);
TASK_PP(16'h8A63,4);
TASK_PP(16'h8A64,4);
TASK_PP(16'h8A65,4);
TASK_PP(16'h8A66,4);
TASK_PP(16'h8A67,4);
TASK_PP(16'h8A68,4);
TASK_PP(16'h8A69,4);
TASK_PP(16'h8A6A,4);
TASK_PP(16'h8A6B,4);
TASK_PP(16'h8A6C,4);
TASK_PP(16'h8A6D,4);
TASK_PP(16'h8A6E,4);
TASK_PP(16'h8A6F,4);
TASK_PP(16'h8A70,4);
TASK_PP(16'h8A71,4);
TASK_PP(16'h8A72,4);
TASK_PP(16'h8A73,4);
TASK_PP(16'h8A74,4);
TASK_PP(16'h8A75,4);
TASK_PP(16'h8A76,4);
TASK_PP(16'h8A77,4);
TASK_PP(16'h8A78,4);
TASK_PP(16'h8A79,4);
TASK_PP(16'h8A7A,4);
TASK_PP(16'h8A7B,4);
TASK_PP(16'h8A7C,4);
TASK_PP(16'h8A7D,4);
TASK_PP(16'h8A7E,4);
TASK_PP(16'h8A7F,4);
TASK_PP(16'h8A80,4);
TASK_PP(16'h8A81,4);
TASK_PP(16'h8A82,4);
TASK_PP(16'h8A83,4);
TASK_PP(16'h8A84,4);
TASK_PP(16'h8A85,4);
TASK_PP(16'h8A86,4);
TASK_PP(16'h8A87,4);
TASK_PP(16'h8A88,4);
TASK_PP(16'h8A89,4);
TASK_PP(16'h8A8A,4);
TASK_PP(16'h8A8B,4);
TASK_PP(16'h8A8C,4);
TASK_PP(16'h8A8D,4);
TASK_PP(16'h8A8E,4);
TASK_PP(16'h8A8F,4);
TASK_PP(16'h8A90,4);
TASK_PP(16'h8A91,4);
TASK_PP(16'h8A92,4);
TASK_PP(16'h8A93,4);
TASK_PP(16'h8A94,4);
TASK_PP(16'h8A95,4);
TASK_PP(16'h8A96,4);
TASK_PP(16'h8A97,4);
TASK_PP(16'h8A98,4);
TASK_PP(16'h8A99,4);
TASK_PP(16'h8A9A,4);
TASK_PP(16'h8A9B,4);
TASK_PP(16'h8A9C,4);
TASK_PP(16'h8A9D,4);
TASK_PP(16'h8A9E,4);
TASK_PP(16'h8A9F,4);
TASK_PP(16'h8AA0,4);
TASK_PP(16'h8AA1,4);
TASK_PP(16'h8AA2,4);
TASK_PP(16'h8AA3,4);
TASK_PP(16'h8AA4,4);
TASK_PP(16'h8AA5,4);
TASK_PP(16'h8AA6,4);
TASK_PP(16'h8AA7,4);
TASK_PP(16'h8AA8,4);
TASK_PP(16'h8AA9,4);
TASK_PP(16'h8AAA,4);
TASK_PP(16'h8AAB,4);
TASK_PP(16'h8AAC,4);
TASK_PP(16'h8AAD,4);
TASK_PP(16'h8AAE,4);
TASK_PP(16'h8AAF,4);
TASK_PP(16'h8AB0,4);
TASK_PP(16'h8AB1,4);
TASK_PP(16'h8AB2,4);
TASK_PP(16'h8AB3,4);
TASK_PP(16'h8AB4,4);
TASK_PP(16'h8AB5,4);
TASK_PP(16'h8AB6,4);
TASK_PP(16'h8AB7,4);
TASK_PP(16'h8AB8,4);
TASK_PP(16'h8AB9,4);
TASK_PP(16'h8ABA,4);
TASK_PP(16'h8ABB,4);
TASK_PP(16'h8ABC,4);
TASK_PP(16'h8ABD,4);
TASK_PP(16'h8ABE,4);
TASK_PP(16'h8ABF,4);
TASK_PP(16'h8AC0,4);
TASK_PP(16'h8AC1,4);
TASK_PP(16'h8AC2,4);
TASK_PP(16'h8AC3,4);
TASK_PP(16'h8AC4,4);
TASK_PP(16'h8AC5,4);
TASK_PP(16'h8AC6,4);
TASK_PP(16'h8AC7,4);
TASK_PP(16'h8AC8,4);
TASK_PP(16'h8AC9,4);
TASK_PP(16'h8ACA,4);
TASK_PP(16'h8ACB,4);
TASK_PP(16'h8ACC,4);
TASK_PP(16'h8ACD,4);
TASK_PP(16'h8ACE,4);
TASK_PP(16'h8ACF,4);
TASK_PP(16'h8AD0,4);
TASK_PP(16'h8AD1,4);
TASK_PP(16'h8AD2,4);
TASK_PP(16'h8AD3,4);
TASK_PP(16'h8AD4,4);
TASK_PP(16'h8AD5,4);
TASK_PP(16'h8AD6,4);
TASK_PP(16'h8AD7,4);
TASK_PP(16'h8AD8,4);
TASK_PP(16'h8AD9,4);
TASK_PP(16'h8ADA,4);
TASK_PP(16'h8ADB,4);
TASK_PP(16'h8ADC,4);
TASK_PP(16'h8ADD,4);
TASK_PP(16'h8ADE,4);
TASK_PP(16'h8ADF,4);
TASK_PP(16'h8AE0,4);
TASK_PP(16'h8AE1,4);
TASK_PP(16'h8AE2,4);
TASK_PP(16'h8AE3,4);
TASK_PP(16'h8AE4,4);
TASK_PP(16'h8AE5,4);
TASK_PP(16'h8AE6,4);
TASK_PP(16'h8AE7,4);
TASK_PP(16'h8AE8,4);
TASK_PP(16'h8AE9,4);
TASK_PP(16'h8AEA,4);
TASK_PP(16'h8AEB,4);
TASK_PP(16'h8AEC,4);
TASK_PP(16'h8AED,4);
TASK_PP(16'h8AEE,4);
TASK_PP(16'h8AEF,4);
TASK_PP(16'h8AF0,4);
TASK_PP(16'h8AF1,4);
TASK_PP(16'h8AF2,4);
TASK_PP(16'h8AF3,4);
TASK_PP(16'h8AF4,4);
TASK_PP(16'h8AF5,4);
TASK_PP(16'h8AF6,4);
TASK_PP(16'h8AF7,4);
TASK_PP(16'h8AF8,4);
TASK_PP(16'h8AF9,4);
TASK_PP(16'h8AFA,4);
TASK_PP(16'h8AFB,4);
TASK_PP(16'h8AFC,4);
TASK_PP(16'h8AFD,4);
TASK_PP(16'h8AFE,4);
TASK_PP(16'h8AFF,4);
TASK_PP(16'h8B00,4);
TASK_PP(16'h8B01,4);
TASK_PP(16'h8B02,4);
TASK_PP(16'h8B03,4);
TASK_PP(16'h8B04,4);
TASK_PP(16'h8B05,4);
TASK_PP(16'h8B06,4);
TASK_PP(16'h8B07,4);
TASK_PP(16'h8B08,4);
TASK_PP(16'h8B09,4);
TASK_PP(16'h8B0A,4);
TASK_PP(16'h8B0B,4);
TASK_PP(16'h8B0C,4);
TASK_PP(16'h8B0D,4);
TASK_PP(16'h8B0E,4);
TASK_PP(16'h8B0F,4);
TASK_PP(16'h8B10,4);
TASK_PP(16'h8B11,4);
TASK_PP(16'h8B12,4);
TASK_PP(16'h8B13,4);
TASK_PP(16'h8B14,4);
TASK_PP(16'h8B15,4);
TASK_PP(16'h8B16,4);
TASK_PP(16'h8B17,4);
TASK_PP(16'h8B18,4);
TASK_PP(16'h8B19,4);
TASK_PP(16'h8B1A,4);
TASK_PP(16'h8B1B,4);
TASK_PP(16'h8B1C,4);
TASK_PP(16'h8B1D,4);
TASK_PP(16'h8B1E,4);
TASK_PP(16'h8B1F,4);
TASK_PP(16'h8B20,4);
TASK_PP(16'h8B21,4);
TASK_PP(16'h8B22,4);
TASK_PP(16'h8B23,4);
TASK_PP(16'h8B24,4);
TASK_PP(16'h8B25,4);
TASK_PP(16'h8B26,4);
TASK_PP(16'h8B27,4);
TASK_PP(16'h8B28,4);
TASK_PP(16'h8B29,4);
TASK_PP(16'h8B2A,4);
TASK_PP(16'h8B2B,4);
TASK_PP(16'h8B2C,4);
TASK_PP(16'h8B2D,4);
TASK_PP(16'h8B2E,4);
TASK_PP(16'h8B2F,4);
TASK_PP(16'h8B30,4);
TASK_PP(16'h8B31,4);
TASK_PP(16'h8B32,4);
TASK_PP(16'h8B33,4);
TASK_PP(16'h8B34,4);
TASK_PP(16'h8B35,4);
TASK_PP(16'h8B36,4);
TASK_PP(16'h8B37,4);
TASK_PP(16'h8B38,4);
TASK_PP(16'h8B39,4);
TASK_PP(16'h8B3A,4);
TASK_PP(16'h8B3B,4);
TASK_PP(16'h8B3C,4);
TASK_PP(16'h8B3D,4);
TASK_PP(16'h8B3E,4);
TASK_PP(16'h8B3F,4);
TASK_PP(16'h8B40,4);
TASK_PP(16'h8B41,4);
TASK_PP(16'h8B42,4);
TASK_PP(16'h8B43,4);
TASK_PP(16'h8B44,4);
TASK_PP(16'h8B45,4);
TASK_PP(16'h8B46,4);
TASK_PP(16'h8B47,4);
TASK_PP(16'h8B48,4);
TASK_PP(16'h8B49,4);
TASK_PP(16'h8B4A,4);
TASK_PP(16'h8B4B,4);
TASK_PP(16'h8B4C,4);
TASK_PP(16'h8B4D,4);
TASK_PP(16'h8B4E,4);
TASK_PP(16'h8B4F,4);
TASK_PP(16'h8B50,4);
TASK_PP(16'h8B51,4);
TASK_PP(16'h8B52,4);
TASK_PP(16'h8B53,4);
TASK_PP(16'h8B54,4);
TASK_PP(16'h8B55,4);
TASK_PP(16'h8B56,4);
TASK_PP(16'h8B57,4);
TASK_PP(16'h8B58,4);
TASK_PP(16'h8B59,4);
TASK_PP(16'h8B5A,4);
TASK_PP(16'h8B5B,4);
TASK_PP(16'h8B5C,4);
TASK_PP(16'h8B5D,4);
TASK_PP(16'h8B5E,4);
TASK_PP(16'h8B5F,4);
TASK_PP(16'h8B60,4);
TASK_PP(16'h8B61,4);
TASK_PP(16'h8B62,4);
TASK_PP(16'h8B63,4);
TASK_PP(16'h8B64,4);
TASK_PP(16'h8B65,4);
TASK_PP(16'h8B66,4);
TASK_PP(16'h8B67,4);
TASK_PP(16'h8B68,4);
TASK_PP(16'h8B69,4);
TASK_PP(16'h8B6A,4);
TASK_PP(16'h8B6B,4);
TASK_PP(16'h8B6C,4);
TASK_PP(16'h8B6D,4);
TASK_PP(16'h8B6E,4);
TASK_PP(16'h8B6F,4);
TASK_PP(16'h8B70,4);
TASK_PP(16'h8B71,4);
TASK_PP(16'h8B72,4);
TASK_PP(16'h8B73,4);
TASK_PP(16'h8B74,4);
TASK_PP(16'h8B75,4);
TASK_PP(16'h8B76,4);
TASK_PP(16'h8B77,4);
TASK_PP(16'h8B78,4);
TASK_PP(16'h8B79,4);
TASK_PP(16'h8B7A,4);
TASK_PP(16'h8B7B,4);
TASK_PP(16'h8B7C,4);
TASK_PP(16'h8B7D,4);
TASK_PP(16'h8B7E,4);
TASK_PP(16'h8B7F,4);
TASK_PP(16'h8B80,4);
TASK_PP(16'h8B81,4);
TASK_PP(16'h8B82,4);
TASK_PP(16'h8B83,4);
TASK_PP(16'h8B84,4);
TASK_PP(16'h8B85,4);
TASK_PP(16'h8B86,4);
TASK_PP(16'h8B87,4);
TASK_PP(16'h8B88,4);
TASK_PP(16'h8B89,4);
TASK_PP(16'h8B8A,4);
TASK_PP(16'h8B8B,4);
TASK_PP(16'h8B8C,4);
TASK_PP(16'h8B8D,4);
TASK_PP(16'h8B8E,4);
TASK_PP(16'h8B8F,4);
TASK_PP(16'h8B90,4);
TASK_PP(16'h8B91,4);
TASK_PP(16'h8B92,4);
TASK_PP(16'h8B93,4);
TASK_PP(16'h8B94,4);
TASK_PP(16'h8B95,4);
TASK_PP(16'h8B96,4);
TASK_PP(16'h8B97,4);
TASK_PP(16'h8B98,4);
TASK_PP(16'h8B99,4);
TASK_PP(16'h8B9A,4);
TASK_PP(16'h8B9B,4);
TASK_PP(16'h8B9C,4);
TASK_PP(16'h8B9D,4);
TASK_PP(16'h8B9E,4);
TASK_PP(16'h8B9F,4);
TASK_PP(16'h8BA0,4);
TASK_PP(16'h8BA1,4);
TASK_PP(16'h8BA2,4);
TASK_PP(16'h8BA3,4);
TASK_PP(16'h8BA4,4);
TASK_PP(16'h8BA5,4);
TASK_PP(16'h8BA6,4);
TASK_PP(16'h8BA7,4);
TASK_PP(16'h8BA8,4);
TASK_PP(16'h8BA9,4);
TASK_PP(16'h8BAA,4);
TASK_PP(16'h8BAB,4);
TASK_PP(16'h8BAC,4);
TASK_PP(16'h8BAD,4);
TASK_PP(16'h8BAE,4);
TASK_PP(16'h8BAF,4);
TASK_PP(16'h8BB0,4);
TASK_PP(16'h8BB1,4);
TASK_PP(16'h8BB2,4);
TASK_PP(16'h8BB3,4);
TASK_PP(16'h8BB4,4);
TASK_PP(16'h8BB5,4);
TASK_PP(16'h8BB6,4);
TASK_PP(16'h8BB7,4);
TASK_PP(16'h8BB8,4);
TASK_PP(16'h8BB9,4);
TASK_PP(16'h8BBA,4);
TASK_PP(16'h8BBB,4);
TASK_PP(16'h8BBC,4);
TASK_PP(16'h8BBD,4);
TASK_PP(16'h8BBE,4);
TASK_PP(16'h8BBF,4);
TASK_PP(16'h8BC0,4);
TASK_PP(16'h8BC1,4);
TASK_PP(16'h8BC2,4);
TASK_PP(16'h8BC3,4);
TASK_PP(16'h8BC4,4);
TASK_PP(16'h8BC5,4);
TASK_PP(16'h8BC6,4);
TASK_PP(16'h8BC7,4);
TASK_PP(16'h8BC8,4);
TASK_PP(16'h8BC9,4);
TASK_PP(16'h8BCA,4);
TASK_PP(16'h8BCB,4);
TASK_PP(16'h8BCC,4);
TASK_PP(16'h8BCD,4);
TASK_PP(16'h8BCE,4);
TASK_PP(16'h8BCF,4);
TASK_PP(16'h8BD0,4);
TASK_PP(16'h8BD1,4);
TASK_PP(16'h8BD2,4);
TASK_PP(16'h8BD3,4);
TASK_PP(16'h8BD4,4);
TASK_PP(16'h8BD5,4);
TASK_PP(16'h8BD6,4);
TASK_PP(16'h8BD7,4);
TASK_PP(16'h8BD8,4);
TASK_PP(16'h8BD9,4);
TASK_PP(16'h8BDA,4);
TASK_PP(16'h8BDB,4);
TASK_PP(16'h8BDC,4);
TASK_PP(16'h8BDD,4);
TASK_PP(16'h8BDE,4);
TASK_PP(16'h8BDF,4);
TASK_PP(16'h8BE0,4);
TASK_PP(16'h8BE1,4);
TASK_PP(16'h8BE2,4);
TASK_PP(16'h8BE3,4);
TASK_PP(16'h8BE4,4);
TASK_PP(16'h8BE5,4);
TASK_PP(16'h8BE6,4);
TASK_PP(16'h8BE7,4);
TASK_PP(16'h8BE8,4);
TASK_PP(16'h8BE9,4);
TASK_PP(16'h8BEA,4);
TASK_PP(16'h8BEB,4);
TASK_PP(16'h8BEC,4);
TASK_PP(16'h8BED,4);
TASK_PP(16'h8BEE,4);
TASK_PP(16'h8BEF,4);
TASK_PP(16'h8BF0,4);
TASK_PP(16'h8BF1,4);
TASK_PP(16'h8BF2,4);
TASK_PP(16'h8BF3,4);
TASK_PP(16'h8BF4,4);
TASK_PP(16'h8BF5,4);
TASK_PP(16'h8BF6,4);
TASK_PP(16'h8BF7,4);
TASK_PP(16'h8BF8,4);
TASK_PP(16'h8BF9,4);
TASK_PP(16'h8BFA,4);
TASK_PP(16'h8BFB,4);
TASK_PP(16'h8BFC,4);
TASK_PP(16'h8BFD,4);
TASK_PP(16'h8BFE,4);
TASK_PP(16'h8BFF,4);
TASK_PP(16'h8C00,4);
TASK_PP(16'h8C01,4);
TASK_PP(16'h8C02,4);
TASK_PP(16'h8C03,4);
TASK_PP(16'h8C04,4);
TASK_PP(16'h8C05,4);
TASK_PP(16'h8C06,4);
TASK_PP(16'h8C07,4);
TASK_PP(16'h8C08,4);
TASK_PP(16'h8C09,4);
TASK_PP(16'h8C0A,4);
TASK_PP(16'h8C0B,4);
TASK_PP(16'h8C0C,4);
TASK_PP(16'h8C0D,4);
TASK_PP(16'h8C0E,4);
TASK_PP(16'h8C0F,4);
TASK_PP(16'h8C10,4);
TASK_PP(16'h8C11,4);
TASK_PP(16'h8C12,4);
TASK_PP(16'h8C13,4);
TASK_PP(16'h8C14,4);
TASK_PP(16'h8C15,4);
TASK_PP(16'h8C16,4);
TASK_PP(16'h8C17,4);
TASK_PP(16'h8C18,4);
TASK_PP(16'h8C19,4);
TASK_PP(16'h8C1A,4);
TASK_PP(16'h8C1B,4);
TASK_PP(16'h8C1C,4);
TASK_PP(16'h8C1D,4);
TASK_PP(16'h8C1E,4);
TASK_PP(16'h8C1F,4);
TASK_PP(16'h8C20,4);
TASK_PP(16'h8C21,4);
TASK_PP(16'h8C22,4);
TASK_PP(16'h8C23,4);
TASK_PP(16'h8C24,4);
TASK_PP(16'h8C25,4);
TASK_PP(16'h8C26,4);
TASK_PP(16'h8C27,4);
TASK_PP(16'h8C28,4);
TASK_PP(16'h8C29,4);
TASK_PP(16'h8C2A,4);
TASK_PP(16'h8C2B,4);
TASK_PP(16'h8C2C,4);
TASK_PP(16'h8C2D,4);
TASK_PP(16'h8C2E,4);
TASK_PP(16'h8C2F,4);
TASK_PP(16'h8C30,4);
TASK_PP(16'h8C31,4);
TASK_PP(16'h8C32,4);
TASK_PP(16'h8C33,4);
TASK_PP(16'h8C34,4);
TASK_PP(16'h8C35,4);
TASK_PP(16'h8C36,4);
TASK_PP(16'h8C37,4);
TASK_PP(16'h8C38,4);
TASK_PP(16'h8C39,4);
TASK_PP(16'h8C3A,4);
TASK_PP(16'h8C3B,4);
TASK_PP(16'h8C3C,4);
TASK_PP(16'h8C3D,4);
TASK_PP(16'h8C3E,4);
TASK_PP(16'h8C3F,4);
TASK_PP(16'h8C40,4);
TASK_PP(16'h8C41,4);
TASK_PP(16'h8C42,4);
TASK_PP(16'h8C43,4);
TASK_PP(16'h8C44,4);
TASK_PP(16'h8C45,4);
TASK_PP(16'h8C46,4);
TASK_PP(16'h8C47,4);
TASK_PP(16'h8C48,4);
TASK_PP(16'h8C49,4);
TASK_PP(16'h8C4A,4);
TASK_PP(16'h8C4B,4);
TASK_PP(16'h8C4C,4);
TASK_PP(16'h8C4D,4);
TASK_PP(16'h8C4E,4);
TASK_PP(16'h8C4F,4);
TASK_PP(16'h8C50,4);
TASK_PP(16'h8C51,4);
TASK_PP(16'h8C52,4);
TASK_PP(16'h8C53,4);
TASK_PP(16'h8C54,4);
TASK_PP(16'h8C55,4);
TASK_PP(16'h8C56,4);
TASK_PP(16'h8C57,4);
TASK_PP(16'h8C58,4);
TASK_PP(16'h8C59,4);
TASK_PP(16'h8C5A,4);
TASK_PP(16'h8C5B,4);
TASK_PP(16'h8C5C,4);
TASK_PP(16'h8C5D,4);
TASK_PP(16'h8C5E,4);
TASK_PP(16'h8C5F,4);
TASK_PP(16'h8C60,4);
TASK_PP(16'h8C61,4);
TASK_PP(16'h8C62,4);
TASK_PP(16'h8C63,4);
TASK_PP(16'h8C64,4);
TASK_PP(16'h8C65,4);
TASK_PP(16'h8C66,4);
TASK_PP(16'h8C67,4);
TASK_PP(16'h8C68,4);
TASK_PP(16'h8C69,4);
TASK_PP(16'h8C6A,4);
TASK_PP(16'h8C6B,4);
TASK_PP(16'h8C6C,4);
TASK_PP(16'h8C6D,4);
TASK_PP(16'h8C6E,4);
TASK_PP(16'h8C6F,4);
TASK_PP(16'h8C70,4);
TASK_PP(16'h8C71,4);
TASK_PP(16'h8C72,4);
TASK_PP(16'h8C73,4);
TASK_PP(16'h8C74,4);
TASK_PP(16'h8C75,4);
TASK_PP(16'h8C76,4);
TASK_PP(16'h8C77,4);
TASK_PP(16'h8C78,4);
TASK_PP(16'h8C79,4);
TASK_PP(16'h8C7A,4);
TASK_PP(16'h8C7B,4);
TASK_PP(16'h8C7C,4);
TASK_PP(16'h8C7D,4);
TASK_PP(16'h8C7E,4);
TASK_PP(16'h8C7F,4);
TASK_PP(16'h8C80,4);
TASK_PP(16'h8C81,4);
TASK_PP(16'h8C82,4);
TASK_PP(16'h8C83,4);
TASK_PP(16'h8C84,4);
TASK_PP(16'h8C85,4);
TASK_PP(16'h8C86,4);
TASK_PP(16'h8C87,4);
TASK_PP(16'h8C88,4);
TASK_PP(16'h8C89,4);
TASK_PP(16'h8C8A,4);
TASK_PP(16'h8C8B,4);
TASK_PP(16'h8C8C,4);
TASK_PP(16'h8C8D,4);
TASK_PP(16'h8C8E,4);
TASK_PP(16'h8C8F,4);
TASK_PP(16'h8C90,4);
TASK_PP(16'h8C91,4);
TASK_PP(16'h8C92,4);
TASK_PP(16'h8C93,4);
TASK_PP(16'h8C94,4);
TASK_PP(16'h8C95,4);
TASK_PP(16'h8C96,4);
TASK_PP(16'h8C97,4);
TASK_PP(16'h8C98,4);
TASK_PP(16'h8C99,4);
TASK_PP(16'h8C9A,4);
TASK_PP(16'h8C9B,4);
TASK_PP(16'h8C9C,4);
TASK_PP(16'h8C9D,4);
TASK_PP(16'h8C9E,4);
TASK_PP(16'h8C9F,4);
TASK_PP(16'h8CA0,4);
TASK_PP(16'h8CA1,4);
TASK_PP(16'h8CA2,4);
TASK_PP(16'h8CA3,4);
TASK_PP(16'h8CA4,4);
TASK_PP(16'h8CA5,4);
TASK_PP(16'h8CA6,4);
TASK_PP(16'h8CA7,4);
TASK_PP(16'h8CA8,4);
TASK_PP(16'h8CA9,4);
TASK_PP(16'h8CAA,4);
TASK_PP(16'h8CAB,4);
TASK_PP(16'h8CAC,4);
TASK_PP(16'h8CAD,4);
TASK_PP(16'h8CAE,4);
TASK_PP(16'h8CAF,4);
TASK_PP(16'h8CB0,4);
TASK_PP(16'h8CB1,4);
TASK_PP(16'h8CB2,4);
TASK_PP(16'h8CB3,4);
TASK_PP(16'h8CB4,4);
TASK_PP(16'h8CB5,4);
TASK_PP(16'h8CB6,4);
TASK_PP(16'h8CB7,4);
TASK_PP(16'h8CB8,4);
TASK_PP(16'h8CB9,4);
TASK_PP(16'h8CBA,4);
TASK_PP(16'h8CBB,4);
TASK_PP(16'h8CBC,4);
TASK_PP(16'h8CBD,4);
TASK_PP(16'h8CBE,4);
TASK_PP(16'h8CBF,4);
TASK_PP(16'h8CC0,4);
TASK_PP(16'h8CC1,4);
TASK_PP(16'h8CC2,4);
TASK_PP(16'h8CC3,4);
TASK_PP(16'h8CC4,4);
TASK_PP(16'h8CC5,4);
TASK_PP(16'h8CC6,4);
TASK_PP(16'h8CC7,4);
TASK_PP(16'h8CC8,4);
TASK_PP(16'h8CC9,4);
TASK_PP(16'h8CCA,4);
TASK_PP(16'h8CCB,4);
TASK_PP(16'h8CCC,4);
TASK_PP(16'h8CCD,4);
TASK_PP(16'h8CCE,4);
TASK_PP(16'h8CCF,4);
TASK_PP(16'h8CD0,4);
TASK_PP(16'h8CD1,4);
TASK_PP(16'h8CD2,4);
TASK_PP(16'h8CD3,4);
TASK_PP(16'h8CD4,4);
TASK_PP(16'h8CD5,4);
TASK_PP(16'h8CD6,4);
TASK_PP(16'h8CD7,4);
TASK_PP(16'h8CD8,4);
TASK_PP(16'h8CD9,4);
TASK_PP(16'h8CDA,4);
TASK_PP(16'h8CDB,4);
TASK_PP(16'h8CDC,4);
TASK_PP(16'h8CDD,4);
TASK_PP(16'h8CDE,4);
TASK_PP(16'h8CDF,4);
TASK_PP(16'h8CE0,4);
TASK_PP(16'h8CE1,4);
TASK_PP(16'h8CE2,4);
TASK_PP(16'h8CE3,4);
TASK_PP(16'h8CE4,4);
TASK_PP(16'h8CE5,4);
TASK_PP(16'h8CE6,4);
TASK_PP(16'h8CE7,4);
TASK_PP(16'h8CE8,4);
TASK_PP(16'h8CE9,4);
TASK_PP(16'h8CEA,4);
TASK_PP(16'h8CEB,4);
TASK_PP(16'h8CEC,4);
TASK_PP(16'h8CED,4);
TASK_PP(16'h8CEE,4);
TASK_PP(16'h8CEF,4);
TASK_PP(16'h8CF0,4);
TASK_PP(16'h8CF1,4);
TASK_PP(16'h8CF2,4);
TASK_PP(16'h8CF3,4);
TASK_PP(16'h8CF4,4);
TASK_PP(16'h8CF5,4);
TASK_PP(16'h8CF6,4);
TASK_PP(16'h8CF7,4);
TASK_PP(16'h8CF8,4);
TASK_PP(16'h8CF9,4);
TASK_PP(16'h8CFA,4);
TASK_PP(16'h8CFB,4);
TASK_PP(16'h8CFC,4);
TASK_PP(16'h8CFD,4);
TASK_PP(16'h8CFE,4);
TASK_PP(16'h8CFF,4);
TASK_PP(16'h8D00,4);
TASK_PP(16'h8D01,4);
TASK_PP(16'h8D02,4);
TASK_PP(16'h8D03,4);
TASK_PP(16'h8D04,4);
TASK_PP(16'h8D05,4);
TASK_PP(16'h8D06,4);
TASK_PP(16'h8D07,4);
TASK_PP(16'h8D08,4);
TASK_PP(16'h8D09,4);
TASK_PP(16'h8D0A,4);
TASK_PP(16'h8D0B,4);
TASK_PP(16'h8D0C,4);
TASK_PP(16'h8D0D,4);
TASK_PP(16'h8D0E,4);
TASK_PP(16'h8D0F,4);
TASK_PP(16'h8D10,4);
TASK_PP(16'h8D11,4);
TASK_PP(16'h8D12,4);
TASK_PP(16'h8D13,4);
TASK_PP(16'h8D14,4);
TASK_PP(16'h8D15,4);
TASK_PP(16'h8D16,4);
TASK_PP(16'h8D17,4);
TASK_PP(16'h8D18,4);
TASK_PP(16'h8D19,4);
TASK_PP(16'h8D1A,4);
TASK_PP(16'h8D1B,4);
TASK_PP(16'h8D1C,4);
TASK_PP(16'h8D1D,4);
TASK_PP(16'h8D1E,4);
TASK_PP(16'h8D1F,4);
TASK_PP(16'h8D20,4);
TASK_PP(16'h8D21,4);
TASK_PP(16'h8D22,4);
TASK_PP(16'h8D23,4);
TASK_PP(16'h8D24,4);
TASK_PP(16'h8D25,4);
TASK_PP(16'h8D26,4);
TASK_PP(16'h8D27,4);
TASK_PP(16'h8D28,4);
TASK_PP(16'h8D29,4);
TASK_PP(16'h8D2A,4);
TASK_PP(16'h8D2B,4);
TASK_PP(16'h8D2C,4);
TASK_PP(16'h8D2D,4);
TASK_PP(16'h8D2E,4);
TASK_PP(16'h8D2F,4);
TASK_PP(16'h8D30,4);
TASK_PP(16'h8D31,4);
TASK_PP(16'h8D32,4);
TASK_PP(16'h8D33,4);
TASK_PP(16'h8D34,4);
TASK_PP(16'h8D35,4);
TASK_PP(16'h8D36,4);
TASK_PP(16'h8D37,4);
TASK_PP(16'h8D38,4);
TASK_PP(16'h8D39,4);
TASK_PP(16'h8D3A,4);
TASK_PP(16'h8D3B,4);
TASK_PP(16'h8D3C,4);
TASK_PP(16'h8D3D,4);
TASK_PP(16'h8D3E,4);
TASK_PP(16'h8D3F,4);
TASK_PP(16'h8D40,4);
TASK_PP(16'h8D41,4);
TASK_PP(16'h8D42,4);
TASK_PP(16'h8D43,4);
TASK_PP(16'h8D44,4);
TASK_PP(16'h8D45,4);
TASK_PP(16'h8D46,4);
TASK_PP(16'h8D47,4);
TASK_PP(16'h8D48,4);
TASK_PP(16'h8D49,4);
TASK_PP(16'h8D4A,4);
TASK_PP(16'h8D4B,4);
TASK_PP(16'h8D4C,4);
TASK_PP(16'h8D4D,4);
TASK_PP(16'h8D4E,4);
TASK_PP(16'h8D4F,4);
TASK_PP(16'h8D50,4);
TASK_PP(16'h8D51,4);
TASK_PP(16'h8D52,4);
TASK_PP(16'h8D53,4);
TASK_PP(16'h8D54,4);
TASK_PP(16'h8D55,4);
TASK_PP(16'h8D56,4);
TASK_PP(16'h8D57,4);
TASK_PP(16'h8D58,4);
TASK_PP(16'h8D59,4);
TASK_PP(16'h8D5A,4);
TASK_PP(16'h8D5B,4);
TASK_PP(16'h8D5C,4);
TASK_PP(16'h8D5D,4);
TASK_PP(16'h8D5E,4);
TASK_PP(16'h8D5F,4);
TASK_PP(16'h8D60,4);
TASK_PP(16'h8D61,4);
TASK_PP(16'h8D62,4);
TASK_PP(16'h8D63,4);
TASK_PP(16'h8D64,4);
TASK_PP(16'h8D65,4);
TASK_PP(16'h8D66,4);
TASK_PP(16'h8D67,4);
TASK_PP(16'h8D68,4);
TASK_PP(16'h8D69,4);
TASK_PP(16'h8D6A,4);
TASK_PP(16'h8D6B,4);
TASK_PP(16'h8D6C,4);
TASK_PP(16'h8D6D,4);
TASK_PP(16'h8D6E,4);
TASK_PP(16'h8D6F,4);
TASK_PP(16'h8D70,4);
TASK_PP(16'h8D71,4);
TASK_PP(16'h8D72,4);
TASK_PP(16'h8D73,4);
TASK_PP(16'h8D74,4);
TASK_PP(16'h8D75,4);
TASK_PP(16'h8D76,4);
TASK_PP(16'h8D77,4);
TASK_PP(16'h8D78,4);
TASK_PP(16'h8D79,4);
TASK_PP(16'h8D7A,4);
TASK_PP(16'h8D7B,4);
TASK_PP(16'h8D7C,4);
TASK_PP(16'h8D7D,4);
TASK_PP(16'h8D7E,4);
TASK_PP(16'h8D7F,4);
TASK_PP(16'h8D80,4);
TASK_PP(16'h8D81,4);
TASK_PP(16'h8D82,4);
TASK_PP(16'h8D83,4);
TASK_PP(16'h8D84,4);
TASK_PP(16'h8D85,4);
TASK_PP(16'h8D86,4);
TASK_PP(16'h8D87,4);
TASK_PP(16'h8D88,4);
TASK_PP(16'h8D89,4);
TASK_PP(16'h8D8A,4);
TASK_PP(16'h8D8B,4);
TASK_PP(16'h8D8C,4);
TASK_PP(16'h8D8D,4);
TASK_PP(16'h8D8E,4);
TASK_PP(16'h8D8F,4);
TASK_PP(16'h8D90,4);
TASK_PP(16'h8D91,4);
TASK_PP(16'h8D92,4);
TASK_PP(16'h8D93,4);
TASK_PP(16'h8D94,4);
TASK_PP(16'h8D95,4);
TASK_PP(16'h8D96,4);
TASK_PP(16'h8D97,4);
TASK_PP(16'h8D98,4);
TASK_PP(16'h8D99,4);
TASK_PP(16'h8D9A,4);
TASK_PP(16'h8D9B,4);
TASK_PP(16'h8D9C,4);
TASK_PP(16'h8D9D,4);
TASK_PP(16'h8D9E,4);
TASK_PP(16'h8D9F,4);
TASK_PP(16'h8DA0,4);
TASK_PP(16'h8DA1,4);
TASK_PP(16'h8DA2,4);
TASK_PP(16'h8DA3,4);
TASK_PP(16'h8DA4,4);
TASK_PP(16'h8DA5,4);
TASK_PP(16'h8DA6,4);
TASK_PP(16'h8DA7,4);
TASK_PP(16'h8DA8,4);
TASK_PP(16'h8DA9,4);
TASK_PP(16'h8DAA,4);
TASK_PP(16'h8DAB,4);
TASK_PP(16'h8DAC,4);
TASK_PP(16'h8DAD,4);
TASK_PP(16'h8DAE,4);
TASK_PP(16'h8DAF,4);
TASK_PP(16'h8DB0,4);
TASK_PP(16'h8DB1,4);
TASK_PP(16'h8DB2,4);
TASK_PP(16'h8DB3,4);
TASK_PP(16'h8DB4,4);
TASK_PP(16'h8DB5,4);
TASK_PP(16'h8DB6,4);
TASK_PP(16'h8DB7,4);
TASK_PP(16'h8DB8,4);
TASK_PP(16'h8DB9,4);
TASK_PP(16'h8DBA,4);
TASK_PP(16'h8DBB,4);
TASK_PP(16'h8DBC,4);
TASK_PP(16'h8DBD,4);
TASK_PP(16'h8DBE,4);
TASK_PP(16'h8DBF,4);
TASK_PP(16'h8DC0,4);
TASK_PP(16'h8DC1,4);
TASK_PP(16'h8DC2,4);
TASK_PP(16'h8DC3,4);
TASK_PP(16'h8DC4,4);
TASK_PP(16'h8DC5,4);
TASK_PP(16'h8DC6,4);
TASK_PP(16'h8DC7,4);
TASK_PP(16'h8DC8,4);
TASK_PP(16'h8DC9,4);
TASK_PP(16'h8DCA,4);
TASK_PP(16'h8DCB,4);
TASK_PP(16'h8DCC,4);
TASK_PP(16'h8DCD,4);
TASK_PP(16'h8DCE,4);
TASK_PP(16'h8DCF,4);
TASK_PP(16'h8DD0,4);
TASK_PP(16'h8DD1,4);
TASK_PP(16'h8DD2,4);
TASK_PP(16'h8DD3,4);
TASK_PP(16'h8DD4,4);
TASK_PP(16'h8DD5,4);
TASK_PP(16'h8DD6,4);
TASK_PP(16'h8DD7,4);
TASK_PP(16'h8DD8,4);
TASK_PP(16'h8DD9,4);
TASK_PP(16'h8DDA,4);
TASK_PP(16'h8DDB,4);
TASK_PP(16'h8DDC,4);
TASK_PP(16'h8DDD,4);
TASK_PP(16'h8DDE,4);
TASK_PP(16'h8DDF,4);
TASK_PP(16'h8DE0,4);
TASK_PP(16'h8DE1,4);
TASK_PP(16'h8DE2,4);
TASK_PP(16'h8DE3,4);
TASK_PP(16'h8DE4,4);
TASK_PP(16'h8DE5,4);
TASK_PP(16'h8DE6,4);
TASK_PP(16'h8DE7,4);
TASK_PP(16'h8DE8,4);
TASK_PP(16'h8DE9,4);
TASK_PP(16'h8DEA,4);
TASK_PP(16'h8DEB,4);
TASK_PP(16'h8DEC,4);
TASK_PP(16'h8DED,4);
TASK_PP(16'h8DEE,4);
TASK_PP(16'h8DEF,4);
TASK_PP(16'h8DF0,4);
TASK_PP(16'h8DF1,4);
TASK_PP(16'h8DF2,4);
TASK_PP(16'h8DF3,4);
TASK_PP(16'h8DF4,4);
TASK_PP(16'h8DF5,4);
TASK_PP(16'h8DF6,4);
TASK_PP(16'h8DF7,4);
TASK_PP(16'h8DF8,4);
TASK_PP(16'h8DF9,4);
TASK_PP(16'h8DFA,4);
TASK_PP(16'h8DFB,4);
TASK_PP(16'h8DFC,4);
TASK_PP(16'h8DFD,4);
TASK_PP(16'h8DFE,4);
TASK_PP(16'h8DFF,4);
TASK_PP(16'h8E00,4);
TASK_PP(16'h8E01,4);
TASK_PP(16'h8E02,4);
TASK_PP(16'h8E03,4);
TASK_PP(16'h8E04,4);
TASK_PP(16'h8E05,4);
TASK_PP(16'h8E06,4);
TASK_PP(16'h8E07,4);
TASK_PP(16'h8E08,4);
TASK_PP(16'h8E09,4);
TASK_PP(16'h8E0A,4);
TASK_PP(16'h8E0B,4);
TASK_PP(16'h8E0C,4);
TASK_PP(16'h8E0D,4);
TASK_PP(16'h8E0E,4);
TASK_PP(16'h8E0F,4);
TASK_PP(16'h8E10,4);
TASK_PP(16'h8E11,4);
TASK_PP(16'h8E12,4);
TASK_PP(16'h8E13,4);
TASK_PP(16'h8E14,4);
TASK_PP(16'h8E15,4);
TASK_PP(16'h8E16,4);
TASK_PP(16'h8E17,4);
TASK_PP(16'h8E18,4);
TASK_PP(16'h8E19,4);
TASK_PP(16'h8E1A,4);
TASK_PP(16'h8E1B,4);
TASK_PP(16'h8E1C,4);
TASK_PP(16'h8E1D,4);
TASK_PP(16'h8E1E,4);
TASK_PP(16'h8E1F,4);
TASK_PP(16'h8E20,4);
TASK_PP(16'h8E21,4);
TASK_PP(16'h8E22,4);
TASK_PP(16'h8E23,4);
TASK_PP(16'h8E24,4);
TASK_PP(16'h8E25,4);
TASK_PP(16'h8E26,4);
TASK_PP(16'h8E27,4);
TASK_PP(16'h8E28,4);
TASK_PP(16'h8E29,4);
TASK_PP(16'h8E2A,4);
TASK_PP(16'h8E2B,4);
TASK_PP(16'h8E2C,4);
TASK_PP(16'h8E2D,4);
TASK_PP(16'h8E2E,4);
TASK_PP(16'h8E2F,4);
TASK_PP(16'h8E30,4);
TASK_PP(16'h8E31,4);
TASK_PP(16'h8E32,4);
TASK_PP(16'h8E33,4);
TASK_PP(16'h8E34,4);
TASK_PP(16'h8E35,4);
TASK_PP(16'h8E36,4);
TASK_PP(16'h8E37,4);
TASK_PP(16'h8E38,4);
TASK_PP(16'h8E39,4);
TASK_PP(16'h8E3A,4);
TASK_PP(16'h8E3B,4);
TASK_PP(16'h8E3C,4);
TASK_PP(16'h8E3D,4);
TASK_PP(16'h8E3E,4);
TASK_PP(16'h8E3F,4);
TASK_PP(16'h8E40,4);
TASK_PP(16'h8E41,4);
TASK_PP(16'h8E42,4);
TASK_PP(16'h8E43,4);
TASK_PP(16'h8E44,4);
TASK_PP(16'h8E45,4);
TASK_PP(16'h8E46,4);
TASK_PP(16'h8E47,4);
TASK_PP(16'h8E48,4);
TASK_PP(16'h8E49,4);
TASK_PP(16'h8E4A,4);
TASK_PP(16'h8E4B,4);
TASK_PP(16'h8E4C,4);
TASK_PP(16'h8E4D,4);
TASK_PP(16'h8E4E,4);
TASK_PP(16'h8E4F,4);
TASK_PP(16'h8E50,4);
TASK_PP(16'h8E51,4);
TASK_PP(16'h8E52,4);
TASK_PP(16'h8E53,4);
TASK_PP(16'h8E54,4);
TASK_PP(16'h8E55,4);
TASK_PP(16'h8E56,4);
TASK_PP(16'h8E57,4);
TASK_PP(16'h8E58,4);
TASK_PP(16'h8E59,4);
TASK_PP(16'h8E5A,4);
TASK_PP(16'h8E5B,4);
TASK_PP(16'h8E5C,4);
TASK_PP(16'h8E5D,4);
TASK_PP(16'h8E5E,4);
TASK_PP(16'h8E5F,4);
TASK_PP(16'h8E60,4);
TASK_PP(16'h8E61,4);
TASK_PP(16'h8E62,4);
TASK_PP(16'h8E63,4);
TASK_PP(16'h8E64,4);
TASK_PP(16'h8E65,4);
TASK_PP(16'h8E66,4);
TASK_PP(16'h8E67,4);
TASK_PP(16'h8E68,4);
TASK_PP(16'h8E69,4);
TASK_PP(16'h8E6A,4);
TASK_PP(16'h8E6B,4);
TASK_PP(16'h8E6C,4);
TASK_PP(16'h8E6D,4);
TASK_PP(16'h8E6E,4);
TASK_PP(16'h8E6F,4);
TASK_PP(16'h8E70,4);
TASK_PP(16'h8E71,4);
TASK_PP(16'h8E72,4);
TASK_PP(16'h8E73,4);
TASK_PP(16'h8E74,4);
TASK_PP(16'h8E75,4);
TASK_PP(16'h8E76,4);
TASK_PP(16'h8E77,4);
TASK_PP(16'h8E78,4);
TASK_PP(16'h8E79,4);
TASK_PP(16'h8E7A,4);
TASK_PP(16'h8E7B,4);
TASK_PP(16'h8E7C,4);
TASK_PP(16'h8E7D,4);
TASK_PP(16'h8E7E,4);
TASK_PP(16'h8E7F,4);
TASK_PP(16'h8E80,4);
TASK_PP(16'h8E81,4);
TASK_PP(16'h8E82,4);
TASK_PP(16'h8E83,4);
TASK_PP(16'h8E84,4);
TASK_PP(16'h8E85,4);
TASK_PP(16'h8E86,4);
TASK_PP(16'h8E87,4);
TASK_PP(16'h8E88,4);
TASK_PP(16'h8E89,4);
TASK_PP(16'h8E8A,4);
TASK_PP(16'h8E8B,4);
TASK_PP(16'h8E8C,4);
TASK_PP(16'h8E8D,4);
TASK_PP(16'h8E8E,4);
TASK_PP(16'h8E8F,4);
TASK_PP(16'h8E90,4);
TASK_PP(16'h8E91,4);
TASK_PP(16'h8E92,4);
TASK_PP(16'h8E93,4);
TASK_PP(16'h8E94,4);
TASK_PP(16'h8E95,4);
TASK_PP(16'h8E96,4);
TASK_PP(16'h8E97,4);
TASK_PP(16'h8E98,4);
TASK_PP(16'h8E99,4);
TASK_PP(16'h8E9A,4);
TASK_PP(16'h8E9B,4);
TASK_PP(16'h8E9C,4);
TASK_PP(16'h8E9D,4);
TASK_PP(16'h8E9E,4);
TASK_PP(16'h8E9F,4);
TASK_PP(16'h8EA0,4);
TASK_PP(16'h8EA1,4);
TASK_PP(16'h8EA2,4);
TASK_PP(16'h8EA3,4);
TASK_PP(16'h8EA4,4);
TASK_PP(16'h8EA5,4);
TASK_PP(16'h8EA6,4);
TASK_PP(16'h8EA7,4);
TASK_PP(16'h8EA8,4);
TASK_PP(16'h8EA9,4);
TASK_PP(16'h8EAA,4);
TASK_PP(16'h8EAB,4);
TASK_PP(16'h8EAC,4);
TASK_PP(16'h8EAD,4);
TASK_PP(16'h8EAE,4);
TASK_PP(16'h8EAF,4);
TASK_PP(16'h8EB0,4);
TASK_PP(16'h8EB1,4);
TASK_PP(16'h8EB2,4);
TASK_PP(16'h8EB3,4);
TASK_PP(16'h8EB4,4);
TASK_PP(16'h8EB5,4);
TASK_PP(16'h8EB6,4);
TASK_PP(16'h8EB7,4);
TASK_PP(16'h8EB8,4);
TASK_PP(16'h8EB9,4);
TASK_PP(16'h8EBA,4);
TASK_PP(16'h8EBB,4);
TASK_PP(16'h8EBC,4);
TASK_PP(16'h8EBD,4);
TASK_PP(16'h8EBE,4);
TASK_PP(16'h8EBF,4);
TASK_PP(16'h8EC0,4);
TASK_PP(16'h8EC1,4);
TASK_PP(16'h8EC2,4);
TASK_PP(16'h8EC3,4);
TASK_PP(16'h8EC4,4);
TASK_PP(16'h8EC5,4);
TASK_PP(16'h8EC6,4);
TASK_PP(16'h8EC7,4);
TASK_PP(16'h8EC8,4);
TASK_PP(16'h8EC9,4);
TASK_PP(16'h8ECA,4);
TASK_PP(16'h8ECB,4);
TASK_PP(16'h8ECC,4);
TASK_PP(16'h8ECD,4);
TASK_PP(16'h8ECE,4);
TASK_PP(16'h8ECF,4);
TASK_PP(16'h8ED0,4);
TASK_PP(16'h8ED1,4);
TASK_PP(16'h8ED2,4);
TASK_PP(16'h8ED3,4);
TASK_PP(16'h8ED4,4);
TASK_PP(16'h8ED5,4);
TASK_PP(16'h8ED6,4);
TASK_PP(16'h8ED7,4);
TASK_PP(16'h8ED8,4);
TASK_PP(16'h8ED9,4);
TASK_PP(16'h8EDA,4);
TASK_PP(16'h8EDB,4);
TASK_PP(16'h8EDC,4);
TASK_PP(16'h8EDD,4);
TASK_PP(16'h8EDE,4);
TASK_PP(16'h8EDF,4);
TASK_PP(16'h8EE0,4);
TASK_PP(16'h8EE1,4);
TASK_PP(16'h8EE2,4);
TASK_PP(16'h8EE3,4);
TASK_PP(16'h8EE4,4);
TASK_PP(16'h8EE5,4);
TASK_PP(16'h8EE6,4);
TASK_PP(16'h8EE7,4);
TASK_PP(16'h8EE8,4);
TASK_PP(16'h8EE9,4);
TASK_PP(16'h8EEA,4);
TASK_PP(16'h8EEB,4);
TASK_PP(16'h8EEC,4);
TASK_PP(16'h8EED,4);
TASK_PP(16'h8EEE,4);
TASK_PP(16'h8EEF,4);
TASK_PP(16'h8EF0,4);
TASK_PP(16'h8EF1,4);
TASK_PP(16'h8EF2,4);
TASK_PP(16'h8EF3,4);
TASK_PP(16'h8EF4,4);
TASK_PP(16'h8EF5,4);
TASK_PP(16'h8EF6,4);
TASK_PP(16'h8EF7,4);
TASK_PP(16'h8EF8,4);
TASK_PP(16'h8EF9,4);
TASK_PP(16'h8EFA,4);
TASK_PP(16'h8EFB,4);
TASK_PP(16'h8EFC,4);
TASK_PP(16'h8EFD,4);
TASK_PP(16'h8EFE,4);
TASK_PP(16'h8EFF,4);
TASK_PP(16'h8F00,4);
TASK_PP(16'h8F01,4);
TASK_PP(16'h8F02,4);
TASK_PP(16'h8F03,4);
TASK_PP(16'h8F04,4);
TASK_PP(16'h8F05,4);
TASK_PP(16'h8F06,4);
TASK_PP(16'h8F07,4);
TASK_PP(16'h8F08,4);
TASK_PP(16'h8F09,4);
TASK_PP(16'h8F0A,4);
TASK_PP(16'h8F0B,4);
TASK_PP(16'h8F0C,4);
TASK_PP(16'h8F0D,4);
TASK_PP(16'h8F0E,4);
TASK_PP(16'h8F0F,4);
TASK_PP(16'h8F10,4);
TASK_PP(16'h8F11,4);
TASK_PP(16'h8F12,4);
TASK_PP(16'h8F13,4);
TASK_PP(16'h8F14,4);
TASK_PP(16'h8F15,4);
TASK_PP(16'h8F16,4);
TASK_PP(16'h8F17,4);
TASK_PP(16'h8F18,4);
TASK_PP(16'h8F19,4);
TASK_PP(16'h8F1A,4);
TASK_PP(16'h8F1B,4);
TASK_PP(16'h8F1C,4);
TASK_PP(16'h8F1D,4);
TASK_PP(16'h8F1E,4);
TASK_PP(16'h8F1F,4);
TASK_PP(16'h8F20,4);
TASK_PP(16'h8F21,4);
TASK_PP(16'h8F22,4);
TASK_PP(16'h8F23,4);
TASK_PP(16'h8F24,4);
TASK_PP(16'h8F25,4);
TASK_PP(16'h8F26,4);
TASK_PP(16'h8F27,4);
TASK_PP(16'h8F28,4);
TASK_PP(16'h8F29,4);
TASK_PP(16'h8F2A,4);
TASK_PP(16'h8F2B,4);
TASK_PP(16'h8F2C,4);
TASK_PP(16'h8F2D,4);
TASK_PP(16'h8F2E,4);
TASK_PP(16'h8F2F,4);
TASK_PP(16'h8F30,4);
TASK_PP(16'h8F31,4);
TASK_PP(16'h8F32,4);
TASK_PP(16'h8F33,4);
TASK_PP(16'h8F34,4);
TASK_PP(16'h8F35,4);
TASK_PP(16'h8F36,4);
TASK_PP(16'h8F37,4);
TASK_PP(16'h8F38,4);
TASK_PP(16'h8F39,4);
TASK_PP(16'h8F3A,4);
TASK_PP(16'h8F3B,4);
TASK_PP(16'h8F3C,4);
TASK_PP(16'h8F3D,4);
TASK_PP(16'h8F3E,4);
TASK_PP(16'h8F3F,4);
TASK_PP(16'h8F40,4);
TASK_PP(16'h8F41,4);
TASK_PP(16'h8F42,4);
TASK_PP(16'h8F43,4);
TASK_PP(16'h8F44,4);
TASK_PP(16'h8F45,4);
TASK_PP(16'h8F46,4);
TASK_PP(16'h8F47,4);
TASK_PP(16'h8F48,4);
TASK_PP(16'h8F49,4);
TASK_PP(16'h8F4A,4);
TASK_PP(16'h8F4B,4);
TASK_PP(16'h8F4C,4);
TASK_PP(16'h8F4D,4);
TASK_PP(16'h8F4E,4);
TASK_PP(16'h8F4F,4);
TASK_PP(16'h8F50,4);
TASK_PP(16'h8F51,4);
TASK_PP(16'h8F52,4);
TASK_PP(16'h8F53,4);
TASK_PP(16'h8F54,4);
TASK_PP(16'h8F55,4);
TASK_PP(16'h8F56,4);
TASK_PP(16'h8F57,4);
TASK_PP(16'h8F58,4);
TASK_PP(16'h8F59,4);
TASK_PP(16'h8F5A,4);
TASK_PP(16'h8F5B,4);
TASK_PP(16'h8F5C,4);
TASK_PP(16'h8F5D,4);
TASK_PP(16'h8F5E,4);
TASK_PP(16'h8F5F,4);
TASK_PP(16'h8F60,4);
TASK_PP(16'h8F61,4);
TASK_PP(16'h8F62,4);
TASK_PP(16'h8F63,4);
TASK_PP(16'h8F64,4);
TASK_PP(16'h8F65,4);
TASK_PP(16'h8F66,4);
TASK_PP(16'h8F67,4);
TASK_PP(16'h8F68,4);
TASK_PP(16'h8F69,4);
TASK_PP(16'h8F6A,4);
TASK_PP(16'h8F6B,4);
TASK_PP(16'h8F6C,4);
TASK_PP(16'h8F6D,4);
TASK_PP(16'h8F6E,4);
TASK_PP(16'h8F6F,4);
TASK_PP(16'h8F70,4);
TASK_PP(16'h8F71,4);
TASK_PP(16'h8F72,4);
TASK_PP(16'h8F73,4);
TASK_PP(16'h8F74,4);
TASK_PP(16'h8F75,4);
TASK_PP(16'h8F76,4);
TASK_PP(16'h8F77,4);
TASK_PP(16'h8F78,4);
TASK_PP(16'h8F79,4);
TASK_PP(16'h8F7A,4);
TASK_PP(16'h8F7B,4);
TASK_PP(16'h8F7C,4);
TASK_PP(16'h8F7D,4);
TASK_PP(16'h8F7E,4);
TASK_PP(16'h8F7F,4);
TASK_PP(16'h8F80,4);
TASK_PP(16'h8F81,4);
TASK_PP(16'h8F82,4);
TASK_PP(16'h8F83,4);
TASK_PP(16'h8F84,4);
TASK_PP(16'h8F85,4);
TASK_PP(16'h8F86,4);
TASK_PP(16'h8F87,4);
TASK_PP(16'h8F88,4);
TASK_PP(16'h8F89,4);
TASK_PP(16'h8F8A,4);
TASK_PP(16'h8F8B,4);
TASK_PP(16'h8F8C,4);
TASK_PP(16'h8F8D,4);
TASK_PP(16'h8F8E,4);
TASK_PP(16'h8F8F,4);
TASK_PP(16'h8F90,4);
TASK_PP(16'h8F91,4);
TASK_PP(16'h8F92,4);
TASK_PP(16'h8F93,4);
TASK_PP(16'h8F94,4);
TASK_PP(16'h8F95,4);
TASK_PP(16'h8F96,4);
TASK_PP(16'h8F97,4);
TASK_PP(16'h8F98,4);
TASK_PP(16'h8F99,4);
TASK_PP(16'h8F9A,4);
TASK_PP(16'h8F9B,4);
TASK_PP(16'h8F9C,4);
TASK_PP(16'h8F9D,4);
TASK_PP(16'h8F9E,4);
TASK_PP(16'h8F9F,4);
TASK_PP(16'h8FA0,4);
TASK_PP(16'h8FA1,4);
TASK_PP(16'h8FA2,4);
TASK_PP(16'h8FA3,4);
TASK_PP(16'h8FA4,4);
TASK_PP(16'h8FA5,4);
TASK_PP(16'h8FA6,4);
TASK_PP(16'h8FA7,4);
TASK_PP(16'h8FA8,4);
TASK_PP(16'h8FA9,4);
TASK_PP(16'h8FAA,4);
TASK_PP(16'h8FAB,4);
TASK_PP(16'h8FAC,4);
TASK_PP(16'h8FAD,4);
TASK_PP(16'h8FAE,4);
TASK_PP(16'h8FAF,4);
TASK_PP(16'h8FB0,4);
TASK_PP(16'h8FB1,4);
TASK_PP(16'h8FB2,4);
TASK_PP(16'h8FB3,4);
TASK_PP(16'h8FB4,4);
TASK_PP(16'h8FB5,4);
TASK_PP(16'h8FB6,4);
TASK_PP(16'h8FB7,4);
TASK_PP(16'h8FB8,4);
TASK_PP(16'h8FB9,4);
TASK_PP(16'h8FBA,4);
TASK_PP(16'h8FBB,4);
TASK_PP(16'h8FBC,4);
TASK_PP(16'h8FBD,4);
TASK_PP(16'h8FBE,4);
TASK_PP(16'h8FBF,4);
TASK_PP(16'h8FC0,4);
TASK_PP(16'h8FC1,4);
TASK_PP(16'h8FC2,4);
TASK_PP(16'h8FC3,4);
TASK_PP(16'h8FC4,4);
TASK_PP(16'h8FC5,4);
TASK_PP(16'h8FC6,4);
TASK_PP(16'h8FC7,4);
TASK_PP(16'h8FC8,4);
TASK_PP(16'h8FC9,4);
TASK_PP(16'h8FCA,4);
TASK_PP(16'h8FCB,4);
TASK_PP(16'h8FCC,4);
TASK_PP(16'h8FCD,4);
TASK_PP(16'h8FCE,4);
TASK_PP(16'h8FCF,4);
TASK_PP(16'h8FD0,4);
TASK_PP(16'h8FD1,4);
TASK_PP(16'h8FD2,4);
TASK_PP(16'h8FD3,4);
TASK_PP(16'h8FD4,4);
TASK_PP(16'h8FD5,4);
TASK_PP(16'h8FD6,4);
TASK_PP(16'h8FD7,4);
TASK_PP(16'h8FD8,4);
TASK_PP(16'h8FD9,4);
TASK_PP(16'h8FDA,4);
TASK_PP(16'h8FDB,4);
TASK_PP(16'h8FDC,4);
TASK_PP(16'h8FDD,4);
TASK_PP(16'h8FDE,4);
TASK_PP(16'h8FDF,4);
TASK_PP(16'h8FE0,4);
TASK_PP(16'h8FE1,4);
TASK_PP(16'h8FE2,4);
TASK_PP(16'h8FE3,4);
TASK_PP(16'h8FE4,4);
TASK_PP(16'h8FE5,4);
TASK_PP(16'h8FE6,4);
TASK_PP(16'h8FE7,4);
TASK_PP(16'h8FE8,4);
TASK_PP(16'h8FE9,4);
TASK_PP(16'h8FEA,4);
TASK_PP(16'h8FEB,4);
TASK_PP(16'h8FEC,4);
TASK_PP(16'h8FED,4);
TASK_PP(16'h8FEE,4);
TASK_PP(16'h8FEF,4);
TASK_PP(16'h8FF0,4);
TASK_PP(16'h8FF1,4);
TASK_PP(16'h8FF2,4);
TASK_PP(16'h8FF3,4);
TASK_PP(16'h8FF4,4);
TASK_PP(16'h8FF5,4);
TASK_PP(16'h8FF6,4);
TASK_PP(16'h8FF7,4);
TASK_PP(16'h8FF8,4);
TASK_PP(16'h8FF9,4);
TASK_PP(16'h8FFA,4);
TASK_PP(16'h8FFB,4);
TASK_PP(16'h8FFC,4);
TASK_PP(16'h8FFD,4);
TASK_PP(16'h8FFE,4);
TASK_PP(16'h8FFF,4);
TASK_PP(16'h9000,4);
TASK_PP(16'h9001,4);
TASK_PP(16'h9002,4);
TASK_PP(16'h9003,4);
TASK_PP(16'h9004,4);
TASK_PP(16'h9005,4);
TASK_PP(16'h9006,4);
TASK_PP(16'h9007,4);
TASK_PP(16'h9008,4);
TASK_PP(16'h9009,4);
TASK_PP(16'h900A,4);
TASK_PP(16'h900B,4);
TASK_PP(16'h900C,4);
TASK_PP(16'h900D,4);
TASK_PP(16'h900E,4);
TASK_PP(16'h900F,4);
TASK_PP(16'h9010,4);
TASK_PP(16'h9011,4);
TASK_PP(16'h9012,4);
TASK_PP(16'h9013,4);
TASK_PP(16'h9014,4);
TASK_PP(16'h9015,4);
TASK_PP(16'h9016,4);
TASK_PP(16'h9017,4);
TASK_PP(16'h9018,4);
TASK_PP(16'h9019,4);
TASK_PP(16'h901A,4);
TASK_PP(16'h901B,4);
TASK_PP(16'h901C,4);
TASK_PP(16'h901D,4);
TASK_PP(16'h901E,4);
TASK_PP(16'h901F,4);
TASK_PP(16'h9020,4);
TASK_PP(16'h9021,4);
TASK_PP(16'h9022,4);
TASK_PP(16'h9023,4);
TASK_PP(16'h9024,4);
TASK_PP(16'h9025,4);
TASK_PP(16'h9026,4);
TASK_PP(16'h9027,4);
TASK_PP(16'h9028,4);
TASK_PP(16'h9029,4);
TASK_PP(16'h902A,4);
TASK_PP(16'h902B,4);
TASK_PP(16'h902C,4);
TASK_PP(16'h902D,4);
TASK_PP(16'h902E,4);
TASK_PP(16'h902F,4);
TASK_PP(16'h9030,4);
TASK_PP(16'h9031,4);
TASK_PP(16'h9032,4);
TASK_PP(16'h9033,4);
TASK_PP(16'h9034,4);
TASK_PP(16'h9035,4);
TASK_PP(16'h9036,4);
TASK_PP(16'h9037,4);
TASK_PP(16'h9038,4);
TASK_PP(16'h9039,4);
TASK_PP(16'h903A,4);
TASK_PP(16'h903B,4);
TASK_PP(16'h903C,4);
TASK_PP(16'h903D,4);
TASK_PP(16'h903E,4);
TASK_PP(16'h903F,4);
TASK_PP(16'h9040,4);
TASK_PP(16'h9041,4);
TASK_PP(16'h9042,4);
TASK_PP(16'h9043,4);
TASK_PP(16'h9044,4);
TASK_PP(16'h9045,4);
TASK_PP(16'h9046,4);
TASK_PP(16'h9047,4);
TASK_PP(16'h9048,4);
TASK_PP(16'h9049,4);
TASK_PP(16'h904A,4);
TASK_PP(16'h904B,4);
TASK_PP(16'h904C,4);
TASK_PP(16'h904D,4);
TASK_PP(16'h904E,4);
TASK_PP(16'h904F,4);
TASK_PP(16'h9050,4);
TASK_PP(16'h9051,4);
TASK_PP(16'h9052,4);
TASK_PP(16'h9053,4);
TASK_PP(16'h9054,4);
TASK_PP(16'h9055,4);
TASK_PP(16'h9056,4);
TASK_PP(16'h9057,4);
TASK_PP(16'h9058,4);
TASK_PP(16'h9059,4);
TASK_PP(16'h905A,4);
TASK_PP(16'h905B,4);
TASK_PP(16'h905C,4);
TASK_PP(16'h905D,4);
TASK_PP(16'h905E,4);
TASK_PP(16'h905F,4);
TASK_PP(16'h9060,4);
TASK_PP(16'h9061,4);
TASK_PP(16'h9062,4);
TASK_PP(16'h9063,4);
TASK_PP(16'h9064,4);
TASK_PP(16'h9065,4);
TASK_PP(16'h9066,4);
TASK_PP(16'h9067,4);
TASK_PP(16'h9068,4);
TASK_PP(16'h9069,4);
TASK_PP(16'h906A,4);
TASK_PP(16'h906B,4);
TASK_PP(16'h906C,4);
TASK_PP(16'h906D,4);
TASK_PP(16'h906E,4);
TASK_PP(16'h906F,4);
TASK_PP(16'h9070,4);
TASK_PP(16'h9071,4);
TASK_PP(16'h9072,4);
TASK_PP(16'h9073,4);
TASK_PP(16'h9074,4);
TASK_PP(16'h9075,4);
TASK_PP(16'h9076,4);
TASK_PP(16'h9077,4);
TASK_PP(16'h9078,4);
TASK_PP(16'h9079,4);
TASK_PP(16'h907A,4);
TASK_PP(16'h907B,4);
TASK_PP(16'h907C,4);
TASK_PP(16'h907D,4);
TASK_PP(16'h907E,4);
TASK_PP(16'h907F,4);
TASK_PP(16'h9080,4);
TASK_PP(16'h9081,4);
TASK_PP(16'h9082,4);
TASK_PP(16'h9083,4);
TASK_PP(16'h9084,4);
TASK_PP(16'h9085,4);
TASK_PP(16'h9086,4);
TASK_PP(16'h9087,4);
TASK_PP(16'h9088,4);
TASK_PP(16'h9089,4);
TASK_PP(16'h908A,4);
TASK_PP(16'h908B,4);
TASK_PP(16'h908C,4);
TASK_PP(16'h908D,4);
TASK_PP(16'h908E,4);
TASK_PP(16'h908F,4);
TASK_PP(16'h9090,4);
TASK_PP(16'h9091,4);
TASK_PP(16'h9092,4);
TASK_PP(16'h9093,4);
TASK_PP(16'h9094,4);
TASK_PP(16'h9095,4);
TASK_PP(16'h9096,4);
TASK_PP(16'h9097,4);
TASK_PP(16'h9098,4);
TASK_PP(16'h9099,4);
TASK_PP(16'h909A,4);
TASK_PP(16'h909B,4);
TASK_PP(16'h909C,4);
TASK_PP(16'h909D,4);
TASK_PP(16'h909E,4);
TASK_PP(16'h909F,4);
TASK_PP(16'h90A0,4);
TASK_PP(16'h90A1,4);
TASK_PP(16'h90A2,4);
TASK_PP(16'h90A3,4);
TASK_PP(16'h90A4,4);
TASK_PP(16'h90A5,4);
TASK_PP(16'h90A6,4);
TASK_PP(16'h90A7,4);
TASK_PP(16'h90A8,4);
TASK_PP(16'h90A9,4);
TASK_PP(16'h90AA,4);
TASK_PP(16'h90AB,4);
TASK_PP(16'h90AC,4);
TASK_PP(16'h90AD,4);
TASK_PP(16'h90AE,4);
TASK_PP(16'h90AF,4);
TASK_PP(16'h90B0,4);
TASK_PP(16'h90B1,4);
TASK_PP(16'h90B2,4);
TASK_PP(16'h90B3,4);
TASK_PP(16'h90B4,4);
TASK_PP(16'h90B5,4);
TASK_PP(16'h90B6,4);
TASK_PP(16'h90B7,4);
TASK_PP(16'h90B8,4);
TASK_PP(16'h90B9,4);
TASK_PP(16'h90BA,4);
TASK_PP(16'h90BB,4);
TASK_PP(16'h90BC,4);
TASK_PP(16'h90BD,4);
TASK_PP(16'h90BE,4);
TASK_PP(16'h90BF,4);
TASK_PP(16'h90C0,4);
TASK_PP(16'h90C1,4);
TASK_PP(16'h90C2,4);
TASK_PP(16'h90C3,4);
TASK_PP(16'h90C4,4);
TASK_PP(16'h90C5,4);
TASK_PP(16'h90C6,4);
TASK_PP(16'h90C7,4);
TASK_PP(16'h90C8,4);
TASK_PP(16'h90C9,4);
TASK_PP(16'h90CA,4);
TASK_PP(16'h90CB,4);
TASK_PP(16'h90CC,4);
TASK_PP(16'h90CD,4);
TASK_PP(16'h90CE,4);
TASK_PP(16'h90CF,4);
TASK_PP(16'h90D0,4);
TASK_PP(16'h90D1,4);
TASK_PP(16'h90D2,4);
TASK_PP(16'h90D3,4);
TASK_PP(16'h90D4,4);
TASK_PP(16'h90D5,4);
TASK_PP(16'h90D6,4);
TASK_PP(16'h90D7,4);
TASK_PP(16'h90D8,4);
TASK_PP(16'h90D9,4);
TASK_PP(16'h90DA,4);
TASK_PP(16'h90DB,4);
TASK_PP(16'h90DC,4);
TASK_PP(16'h90DD,4);
TASK_PP(16'h90DE,4);
TASK_PP(16'h90DF,4);
TASK_PP(16'h90E0,4);
TASK_PP(16'h90E1,4);
TASK_PP(16'h90E2,4);
TASK_PP(16'h90E3,4);
TASK_PP(16'h90E4,4);
TASK_PP(16'h90E5,4);
TASK_PP(16'h90E6,4);
TASK_PP(16'h90E7,4);
TASK_PP(16'h90E8,4);
TASK_PP(16'h90E9,4);
TASK_PP(16'h90EA,4);
TASK_PP(16'h90EB,4);
TASK_PP(16'h90EC,4);
TASK_PP(16'h90ED,4);
TASK_PP(16'h90EE,4);
TASK_PP(16'h90EF,4);
TASK_PP(16'h90F0,4);
TASK_PP(16'h90F1,4);
TASK_PP(16'h90F2,4);
TASK_PP(16'h90F3,4);
TASK_PP(16'h90F4,4);
TASK_PP(16'h90F5,4);
TASK_PP(16'h90F6,4);
TASK_PP(16'h90F7,4);
TASK_PP(16'h90F8,4);
TASK_PP(16'h90F9,4);
TASK_PP(16'h90FA,4);
TASK_PP(16'h90FB,4);
TASK_PP(16'h90FC,4);
TASK_PP(16'h90FD,4);
TASK_PP(16'h90FE,4);
TASK_PP(16'h90FF,4);
TASK_PP(16'h9100,4);
TASK_PP(16'h9101,4);
TASK_PP(16'h9102,4);
TASK_PP(16'h9103,4);
TASK_PP(16'h9104,4);
TASK_PP(16'h9105,4);
TASK_PP(16'h9106,4);
TASK_PP(16'h9107,4);
TASK_PP(16'h9108,4);
TASK_PP(16'h9109,4);
TASK_PP(16'h910A,4);
TASK_PP(16'h910B,4);
TASK_PP(16'h910C,4);
TASK_PP(16'h910D,4);
TASK_PP(16'h910E,4);
TASK_PP(16'h910F,4);
TASK_PP(16'h9110,4);
TASK_PP(16'h9111,4);
TASK_PP(16'h9112,4);
TASK_PP(16'h9113,4);
TASK_PP(16'h9114,4);
TASK_PP(16'h9115,4);
TASK_PP(16'h9116,4);
TASK_PP(16'h9117,4);
TASK_PP(16'h9118,4);
TASK_PP(16'h9119,4);
TASK_PP(16'h911A,4);
TASK_PP(16'h911B,4);
TASK_PP(16'h911C,4);
TASK_PP(16'h911D,4);
TASK_PP(16'h911E,4);
TASK_PP(16'h911F,4);
TASK_PP(16'h9120,4);
TASK_PP(16'h9121,4);
TASK_PP(16'h9122,4);
TASK_PP(16'h9123,4);
TASK_PP(16'h9124,4);
TASK_PP(16'h9125,4);
TASK_PP(16'h9126,4);
TASK_PP(16'h9127,4);
TASK_PP(16'h9128,4);
TASK_PP(16'h9129,4);
TASK_PP(16'h912A,4);
TASK_PP(16'h912B,4);
TASK_PP(16'h912C,4);
TASK_PP(16'h912D,4);
TASK_PP(16'h912E,4);
TASK_PP(16'h912F,4);
TASK_PP(16'h9130,4);
TASK_PP(16'h9131,4);
TASK_PP(16'h9132,4);
TASK_PP(16'h9133,4);
TASK_PP(16'h9134,4);
TASK_PP(16'h9135,4);
TASK_PP(16'h9136,4);
TASK_PP(16'h9137,4);
TASK_PP(16'h9138,4);
TASK_PP(16'h9139,4);
TASK_PP(16'h913A,4);
TASK_PP(16'h913B,4);
TASK_PP(16'h913C,4);
TASK_PP(16'h913D,4);
TASK_PP(16'h913E,4);
TASK_PP(16'h913F,4);
TASK_PP(16'h9140,4);
TASK_PP(16'h9141,4);
TASK_PP(16'h9142,4);
TASK_PP(16'h9143,4);
TASK_PP(16'h9144,4);
TASK_PP(16'h9145,4);
TASK_PP(16'h9146,4);
TASK_PP(16'h9147,4);
TASK_PP(16'h9148,4);
TASK_PP(16'h9149,4);
TASK_PP(16'h914A,4);
TASK_PP(16'h914B,4);
TASK_PP(16'h914C,4);
TASK_PP(16'h914D,4);
TASK_PP(16'h914E,4);
TASK_PP(16'h914F,4);
TASK_PP(16'h9150,4);
TASK_PP(16'h9151,4);
TASK_PP(16'h9152,4);
TASK_PP(16'h9153,4);
TASK_PP(16'h9154,4);
TASK_PP(16'h9155,4);
TASK_PP(16'h9156,4);
TASK_PP(16'h9157,4);
TASK_PP(16'h9158,4);
TASK_PP(16'h9159,4);
TASK_PP(16'h915A,4);
TASK_PP(16'h915B,4);
TASK_PP(16'h915C,4);
TASK_PP(16'h915D,4);
TASK_PP(16'h915E,4);
TASK_PP(16'h915F,4);
TASK_PP(16'h9160,4);
TASK_PP(16'h9161,4);
TASK_PP(16'h9162,4);
TASK_PP(16'h9163,4);
TASK_PP(16'h9164,4);
TASK_PP(16'h9165,4);
TASK_PP(16'h9166,4);
TASK_PP(16'h9167,4);
TASK_PP(16'h9168,4);
TASK_PP(16'h9169,4);
TASK_PP(16'h916A,4);
TASK_PP(16'h916B,4);
TASK_PP(16'h916C,4);
TASK_PP(16'h916D,4);
TASK_PP(16'h916E,4);
TASK_PP(16'h916F,4);
TASK_PP(16'h9170,4);
TASK_PP(16'h9171,4);
TASK_PP(16'h9172,4);
TASK_PP(16'h9173,4);
TASK_PP(16'h9174,4);
TASK_PP(16'h9175,4);
TASK_PP(16'h9176,4);
TASK_PP(16'h9177,4);
TASK_PP(16'h9178,4);
TASK_PP(16'h9179,4);
TASK_PP(16'h917A,4);
TASK_PP(16'h917B,4);
TASK_PP(16'h917C,4);
TASK_PP(16'h917D,4);
TASK_PP(16'h917E,4);
TASK_PP(16'h917F,4);
TASK_PP(16'h9180,4);
TASK_PP(16'h9181,4);
TASK_PP(16'h9182,4);
TASK_PP(16'h9183,4);
TASK_PP(16'h9184,4);
TASK_PP(16'h9185,4);
TASK_PP(16'h9186,4);
TASK_PP(16'h9187,4);
TASK_PP(16'h9188,4);
TASK_PP(16'h9189,4);
TASK_PP(16'h918A,4);
TASK_PP(16'h918B,4);
TASK_PP(16'h918C,4);
TASK_PP(16'h918D,4);
TASK_PP(16'h918E,4);
TASK_PP(16'h918F,4);
TASK_PP(16'h9190,4);
TASK_PP(16'h9191,4);
TASK_PP(16'h9192,4);
TASK_PP(16'h9193,4);
TASK_PP(16'h9194,4);
TASK_PP(16'h9195,4);
TASK_PP(16'h9196,4);
TASK_PP(16'h9197,4);
TASK_PP(16'h9198,4);
TASK_PP(16'h9199,4);
TASK_PP(16'h919A,4);
TASK_PP(16'h919B,4);
TASK_PP(16'h919C,4);
TASK_PP(16'h919D,4);
TASK_PP(16'h919E,4);
TASK_PP(16'h919F,4);
TASK_PP(16'h91A0,4);
TASK_PP(16'h91A1,4);
TASK_PP(16'h91A2,4);
TASK_PP(16'h91A3,4);
TASK_PP(16'h91A4,4);
TASK_PP(16'h91A5,4);
TASK_PP(16'h91A6,4);
TASK_PP(16'h91A7,4);
TASK_PP(16'h91A8,4);
TASK_PP(16'h91A9,4);
TASK_PP(16'h91AA,4);
TASK_PP(16'h91AB,4);
TASK_PP(16'h91AC,4);
TASK_PP(16'h91AD,4);
TASK_PP(16'h91AE,4);
TASK_PP(16'h91AF,4);
TASK_PP(16'h91B0,4);
TASK_PP(16'h91B1,4);
TASK_PP(16'h91B2,4);
TASK_PP(16'h91B3,4);
TASK_PP(16'h91B4,4);
TASK_PP(16'h91B5,4);
TASK_PP(16'h91B6,4);
TASK_PP(16'h91B7,4);
TASK_PP(16'h91B8,4);
TASK_PP(16'h91B9,4);
TASK_PP(16'h91BA,4);
TASK_PP(16'h91BB,4);
TASK_PP(16'h91BC,4);
TASK_PP(16'h91BD,4);
TASK_PP(16'h91BE,4);
TASK_PP(16'h91BF,4);
TASK_PP(16'h91C0,4);
TASK_PP(16'h91C1,4);
TASK_PP(16'h91C2,4);
TASK_PP(16'h91C3,4);
TASK_PP(16'h91C4,4);
TASK_PP(16'h91C5,4);
TASK_PP(16'h91C6,4);
TASK_PP(16'h91C7,4);
TASK_PP(16'h91C8,4);
TASK_PP(16'h91C9,4);
TASK_PP(16'h91CA,4);
TASK_PP(16'h91CB,4);
TASK_PP(16'h91CC,4);
TASK_PP(16'h91CD,4);
TASK_PP(16'h91CE,4);
TASK_PP(16'h91CF,4);
TASK_PP(16'h91D0,4);
TASK_PP(16'h91D1,4);
TASK_PP(16'h91D2,4);
TASK_PP(16'h91D3,4);
TASK_PP(16'h91D4,4);
TASK_PP(16'h91D5,4);
TASK_PP(16'h91D6,4);
TASK_PP(16'h91D7,4);
TASK_PP(16'h91D8,4);
TASK_PP(16'h91D9,4);
TASK_PP(16'h91DA,4);
TASK_PP(16'h91DB,4);
TASK_PP(16'h91DC,4);
TASK_PP(16'h91DD,4);
TASK_PP(16'h91DE,4);
TASK_PP(16'h91DF,4);
TASK_PP(16'h91E0,4);
TASK_PP(16'h91E1,4);
TASK_PP(16'h91E2,4);
TASK_PP(16'h91E3,4);
TASK_PP(16'h91E4,4);
TASK_PP(16'h91E5,4);
TASK_PP(16'h91E6,4);
TASK_PP(16'h91E7,4);
TASK_PP(16'h91E8,4);
TASK_PP(16'h91E9,4);
TASK_PP(16'h91EA,4);
TASK_PP(16'h91EB,4);
TASK_PP(16'h91EC,4);
TASK_PP(16'h91ED,4);
TASK_PP(16'h91EE,4);
TASK_PP(16'h91EF,4);
TASK_PP(16'h91F0,4);
TASK_PP(16'h91F1,4);
TASK_PP(16'h91F2,4);
TASK_PP(16'h91F3,4);
TASK_PP(16'h91F4,4);
TASK_PP(16'h91F5,4);
TASK_PP(16'h91F6,4);
TASK_PP(16'h91F7,4);
TASK_PP(16'h91F8,4);
TASK_PP(16'h91F9,4);
TASK_PP(16'h91FA,4);
TASK_PP(16'h91FB,4);
TASK_PP(16'h91FC,4);
TASK_PP(16'h91FD,4);
TASK_PP(16'h91FE,4);
TASK_PP(16'h91FF,4);
TASK_PP(16'h9200,4);
TASK_PP(16'h9201,4);
TASK_PP(16'h9202,4);
TASK_PP(16'h9203,4);
TASK_PP(16'h9204,4);
TASK_PP(16'h9205,4);
TASK_PP(16'h9206,4);
TASK_PP(16'h9207,4);
TASK_PP(16'h9208,4);
TASK_PP(16'h9209,4);
TASK_PP(16'h920A,4);
TASK_PP(16'h920B,4);
TASK_PP(16'h920C,4);
TASK_PP(16'h920D,4);
TASK_PP(16'h920E,4);
TASK_PP(16'h920F,4);
TASK_PP(16'h9210,4);
TASK_PP(16'h9211,4);
TASK_PP(16'h9212,4);
TASK_PP(16'h9213,4);
TASK_PP(16'h9214,4);
TASK_PP(16'h9215,4);
TASK_PP(16'h9216,4);
TASK_PP(16'h9217,4);
TASK_PP(16'h9218,4);
TASK_PP(16'h9219,4);
TASK_PP(16'h921A,4);
TASK_PP(16'h921B,4);
TASK_PP(16'h921C,4);
TASK_PP(16'h921D,4);
TASK_PP(16'h921E,4);
TASK_PP(16'h921F,4);
TASK_PP(16'h9220,4);
TASK_PP(16'h9221,4);
TASK_PP(16'h9222,4);
TASK_PP(16'h9223,4);
TASK_PP(16'h9224,4);
TASK_PP(16'h9225,4);
TASK_PP(16'h9226,4);
TASK_PP(16'h9227,4);
TASK_PP(16'h9228,4);
TASK_PP(16'h9229,4);
TASK_PP(16'h922A,4);
TASK_PP(16'h922B,4);
TASK_PP(16'h922C,4);
TASK_PP(16'h922D,4);
TASK_PP(16'h922E,4);
TASK_PP(16'h922F,4);
TASK_PP(16'h9230,4);
TASK_PP(16'h9231,4);
TASK_PP(16'h9232,4);
TASK_PP(16'h9233,4);
TASK_PP(16'h9234,4);
TASK_PP(16'h9235,4);
TASK_PP(16'h9236,4);
TASK_PP(16'h9237,4);
TASK_PP(16'h9238,4);
TASK_PP(16'h9239,4);
TASK_PP(16'h923A,4);
TASK_PP(16'h923B,4);
TASK_PP(16'h923C,4);
TASK_PP(16'h923D,4);
TASK_PP(16'h923E,4);
TASK_PP(16'h923F,4);
TASK_PP(16'h9240,4);
TASK_PP(16'h9241,4);
TASK_PP(16'h9242,4);
TASK_PP(16'h9243,4);
TASK_PP(16'h9244,4);
TASK_PP(16'h9245,4);
TASK_PP(16'h9246,4);
TASK_PP(16'h9247,4);
TASK_PP(16'h9248,4);
TASK_PP(16'h9249,4);
TASK_PP(16'h924A,4);
TASK_PP(16'h924B,4);
TASK_PP(16'h924C,4);
TASK_PP(16'h924D,4);
TASK_PP(16'h924E,4);
TASK_PP(16'h924F,4);
TASK_PP(16'h9250,4);
TASK_PP(16'h9251,4);
TASK_PP(16'h9252,4);
TASK_PP(16'h9253,4);
TASK_PP(16'h9254,4);
TASK_PP(16'h9255,4);
TASK_PP(16'h9256,4);
TASK_PP(16'h9257,4);
TASK_PP(16'h9258,4);
TASK_PP(16'h9259,4);
TASK_PP(16'h925A,4);
TASK_PP(16'h925B,4);
TASK_PP(16'h925C,4);
TASK_PP(16'h925D,4);
TASK_PP(16'h925E,4);
TASK_PP(16'h925F,4);
TASK_PP(16'h9260,4);
TASK_PP(16'h9261,4);
TASK_PP(16'h9262,4);
TASK_PP(16'h9263,4);
TASK_PP(16'h9264,4);
TASK_PP(16'h9265,4);
TASK_PP(16'h9266,4);
TASK_PP(16'h9267,4);
TASK_PP(16'h9268,4);
TASK_PP(16'h9269,4);
TASK_PP(16'h926A,4);
TASK_PP(16'h926B,4);
TASK_PP(16'h926C,4);
TASK_PP(16'h926D,4);
TASK_PP(16'h926E,4);
TASK_PP(16'h926F,4);
TASK_PP(16'h9270,4);
TASK_PP(16'h9271,4);
TASK_PP(16'h9272,4);
TASK_PP(16'h9273,4);
TASK_PP(16'h9274,4);
TASK_PP(16'h9275,4);
TASK_PP(16'h9276,4);
TASK_PP(16'h9277,4);
TASK_PP(16'h9278,4);
TASK_PP(16'h9279,4);
TASK_PP(16'h927A,4);
TASK_PP(16'h927B,4);
TASK_PP(16'h927C,4);
TASK_PP(16'h927D,4);
TASK_PP(16'h927E,4);
TASK_PP(16'h927F,4);
TASK_PP(16'h9280,4);
TASK_PP(16'h9281,4);
TASK_PP(16'h9282,4);
TASK_PP(16'h9283,4);
TASK_PP(16'h9284,4);
TASK_PP(16'h9285,4);
TASK_PP(16'h9286,4);
TASK_PP(16'h9287,4);
TASK_PP(16'h9288,4);
TASK_PP(16'h9289,4);
TASK_PP(16'h928A,4);
TASK_PP(16'h928B,4);
TASK_PP(16'h928C,4);
TASK_PP(16'h928D,4);
TASK_PP(16'h928E,4);
TASK_PP(16'h928F,4);
TASK_PP(16'h9290,4);
TASK_PP(16'h9291,4);
TASK_PP(16'h9292,4);
TASK_PP(16'h9293,4);
TASK_PP(16'h9294,4);
TASK_PP(16'h9295,4);
TASK_PP(16'h9296,4);
TASK_PP(16'h9297,4);
TASK_PP(16'h9298,4);
TASK_PP(16'h9299,4);
TASK_PP(16'h929A,4);
TASK_PP(16'h929B,4);
TASK_PP(16'h929C,4);
TASK_PP(16'h929D,4);
TASK_PP(16'h929E,4);
TASK_PP(16'h929F,4);
TASK_PP(16'h92A0,4);
TASK_PP(16'h92A1,4);
TASK_PP(16'h92A2,4);
TASK_PP(16'h92A3,4);
TASK_PP(16'h92A4,4);
TASK_PP(16'h92A5,4);
TASK_PP(16'h92A6,4);
TASK_PP(16'h92A7,4);
TASK_PP(16'h92A8,4);
TASK_PP(16'h92A9,4);
TASK_PP(16'h92AA,4);
TASK_PP(16'h92AB,4);
TASK_PP(16'h92AC,4);
TASK_PP(16'h92AD,4);
TASK_PP(16'h92AE,4);
TASK_PP(16'h92AF,4);
TASK_PP(16'h92B0,4);
TASK_PP(16'h92B1,4);
TASK_PP(16'h92B2,4);
TASK_PP(16'h92B3,4);
TASK_PP(16'h92B4,4);
TASK_PP(16'h92B5,4);
TASK_PP(16'h92B6,4);
TASK_PP(16'h92B7,4);
TASK_PP(16'h92B8,4);
TASK_PP(16'h92B9,4);
TASK_PP(16'h92BA,4);
TASK_PP(16'h92BB,4);
TASK_PP(16'h92BC,4);
TASK_PP(16'h92BD,4);
TASK_PP(16'h92BE,4);
TASK_PP(16'h92BF,4);
TASK_PP(16'h92C0,4);
TASK_PP(16'h92C1,4);
TASK_PP(16'h92C2,4);
TASK_PP(16'h92C3,4);
TASK_PP(16'h92C4,4);
TASK_PP(16'h92C5,4);
TASK_PP(16'h92C6,4);
TASK_PP(16'h92C7,4);
TASK_PP(16'h92C8,4);
TASK_PP(16'h92C9,4);
TASK_PP(16'h92CA,4);
TASK_PP(16'h92CB,4);
TASK_PP(16'h92CC,4);
TASK_PP(16'h92CD,4);
TASK_PP(16'h92CE,4);
TASK_PP(16'h92CF,4);
TASK_PP(16'h92D0,4);
TASK_PP(16'h92D1,4);
TASK_PP(16'h92D2,4);
TASK_PP(16'h92D3,4);
TASK_PP(16'h92D4,4);
TASK_PP(16'h92D5,4);
TASK_PP(16'h92D6,4);
TASK_PP(16'h92D7,4);
TASK_PP(16'h92D8,4);
TASK_PP(16'h92D9,4);
TASK_PP(16'h92DA,4);
TASK_PP(16'h92DB,4);
TASK_PP(16'h92DC,4);
TASK_PP(16'h92DD,4);
TASK_PP(16'h92DE,4);
TASK_PP(16'h92DF,4);
TASK_PP(16'h92E0,4);
TASK_PP(16'h92E1,4);
TASK_PP(16'h92E2,4);
TASK_PP(16'h92E3,4);
TASK_PP(16'h92E4,4);
TASK_PP(16'h92E5,4);
TASK_PP(16'h92E6,4);
TASK_PP(16'h92E7,4);
TASK_PP(16'h92E8,4);
TASK_PP(16'h92E9,4);
TASK_PP(16'h92EA,4);
TASK_PP(16'h92EB,4);
TASK_PP(16'h92EC,4);
TASK_PP(16'h92ED,4);
TASK_PP(16'h92EE,4);
TASK_PP(16'h92EF,4);
TASK_PP(16'h92F0,4);
TASK_PP(16'h92F1,4);
TASK_PP(16'h92F2,4);
TASK_PP(16'h92F3,4);
TASK_PP(16'h92F4,4);
TASK_PP(16'h92F5,4);
TASK_PP(16'h92F6,4);
TASK_PP(16'h92F7,4);
TASK_PP(16'h92F8,4);
TASK_PP(16'h92F9,4);
TASK_PP(16'h92FA,4);
TASK_PP(16'h92FB,4);
TASK_PP(16'h92FC,4);
TASK_PP(16'h92FD,4);
TASK_PP(16'h92FE,4);
TASK_PP(16'h92FF,4);
TASK_PP(16'h9300,4);
TASK_PP(16'h9301,4);
TASK_PP(16'h9302,4);
TASK_PP(16'h9303,4);
TASK_PP(16'h9304,4);
TASK_PP(16'h9305,4);
TASK_PP(16'h9306,4);
TASK_PP(16'h9307,4);
TASK_PP(16'h9308,4);
TASK_PP(16'h9309,4);
TASK_PP(16'h930A,4);
TASK_PP(16'h930B,4);
TASK_PP(16'h930C,4);
TASK_PP(16'h930D,4);
TASK_PP(16'h930E,4);
TASK_PP(16'h930F,4);
TASK_PP(16'h9310,4);
TASK_PP(16'h9311,4);
TASK_PP(16'h9312,4);
TASK_PP(16'h9313,4);
TASK_PP(16'h9314,4);
TASK_PP(16'h9315,4);
TASK_PP(16'h9316,4);
TASK_PP(16'h9317,4);
TASK_PP(16'h9318,4);
TASK_PP(16'h9319,4);
TASK_PP(16'h931A,4);
TASK_PP(16'h931B,4);
TASK_PP(16'h931C,4);
TASK_PP(16'h931D,4);
TASK_PP(16'h931E,4);
TASK_PP(16'h931F,4);
TASK_PP(16'h9320,4);
TASK_PP(16'h9321,4);
TASK_PP(16'h9322,4);
TASK_PP(16'h9323,4);
TASK_PP(16'h9324,4);
TASK_PP(16'h9325,4);
TASK_PP(16'h9326,4);
TASK_PP(16'h9327,4);
TASK_PP(16'h9328,4);
TASK_PP(16'h9329,4);
TASK_PP(16'h932A,4);
TASK_PP(16'h932B,4);
TASK_PP(16'h932C,4);
TASK_PP(16'h932D,4);
TASK_PP(16'h932E,4);
TASK_PP(16'h932F,4);
TASK_PP(16'h9330,4);
TASK_PP(16'h9331,4);
TASK_PP(16'h9332,4);
TASK_PP(16'h9333,4);
TASK_PP(16'h9334,4);
TASK_PP(16'h9335,4);
TASK_PP(16'h9336,4);
TASK_PP(16'h9337,4);
TASK_PP(16'h9338,4);
TASK_PP(16'h9339,4);
TASK_PP(16'h933A,4);
TASK_PP(16'h933B,4);
TASK_PP(16'h933C,4);
TASK_PP(16'h933D,4);
TASK_PP(16'h933E,4);
TASK_PP(16'h933F,4);
TASK_PP(16'h9340,4);
TASK_PP(16'h9341,4);
TASK_PP(16'h9342,4);
TASK_PP(16'h9343,4);
TASK_PP(16'h9344,4);
TASK_PP(16'h9345,4);
TASK_PP(16'h9346,4);
TASK_PP(16'h9347,4);
TASK_PP(16'h9348,4);
TASK_PP(16'h9349,4);
TASK_PP(16'h934A,4);
TASK_PP(16'h934B,4);
TASK_PP(16'h934C,4);
TASK_PP(16'h934D,4);
TASK_PP(16'h934E,4);
TASK_PP(16'h934F,4);
TASK_PP(16'h9350,4);
TASK_PP(16'h9351,4);
TASK_PP(16'h9352,4);
TASK_PP(16'h9353,4);
TASK_PP(16'h9354,4);
TASK_PP(16'h9355,4);
TASK_PP(16'h9356,4);
TASK_PP(16'h9357,4);
TASK_PP(16'h9358,4);
TASK_PP(16'h9359,4);
TASK_PP(16'h935A,4);
TASK_PP(16'h935B,4);
TASK_PP(16'h935C,4);
TASK_PP(16'h935D,4);
TASK_PP(16'h935E,4);
TASK_PP(16'h935F,4);
TASK_PP(16'h9360,4);
TASK_PP(16'h9361,4);
TASK_PP(16'h9362,4);
TASK_PP(16'h9363,4);
TASK_PP(16'h9364,4);
TASK_PP(16'h9365,4);
TASK_PP(16'h9366,4);
TASK_PP(16'h9367,4);
TASK_PP(16'h9368,4);
TASK_PP(16'h9369,4);
TASK_PP(16'h936A,4);
TASK_PP(16'h936B,4);
TASK_PP(16'h936C,4);
TASK_PP(16'h936D,4);
TASK_PP(16'h936E,4);
TASK_PP(16'h936F,4);
TASK_PP(16'h9370,4);
TASK_PP(16'h9371,4);
TASK_PP(16'h9372,4);
TASK_PP(16'h9373,4);
TASK_PP(16'h9374,4);
TASK_PP(16'h9375,4);
TASK_PP(16'h9376,4);
TASK_PP(16'h9377,4);
TASK_PP(16'h9378,4);
TASK_PP(16'h9379,4);
TASK_PP(16'h937A,4);
TASK_PP(16'h937B,4);
TASK_PP(16'h937C,4);
TASK_PP(16'h937D,4);
TASK_PP(16'h937E,4);
TASK_PP(16'h937F,4);
TASK_PP(16'h9380,4);
TASK_PP(16'h9381,4);
TASK_PP(16'h9382,4);
TASK_PP(16'h9383,4);
TASK_PP(16'h9384,4);
TASK_PP(16'h9385,4);
TASK_PP(16'h9386,4);
TASK_PP(16'h9387,4);
TASK_PP(16'h9388,4);
TASK_PP(16'h9389,4);
TASK_PP(16'h938A,4);
TASK_PP(16'h938B,4);
TASK_PP(16'h938C,4);
TASK_PP(16'h938D,4);
TASK_PP(16'h938E,4);
TASK_PP(16'h938F,4);
TASK_PP(16'h9390,4);
TASK_PP(16'h9391,4);
TASK_PP(16'h9392,4);
TASK_PP(16'h9393,4);
TASK_PP(16'h9394,4);
TASK_PP(16'h9395,4);
TASK_PP(16'h9396,4);
TASK_PP(16'h9397,4);
TASK_PP(16'h9398,4);
TASK_PP(16'h9399,4);
TASK_PP(16'h939A,4);
TASK_PP(16'h939B,4);
TASK_PP(16'h939C,4);
TASK_PP(16'h939D,4);
TASK_PP(16'h939E,4);
TASK_PP(16'h939F,4);
TASK_PP(16'h93A0,4);
TASK_PP(16'h93A1,4);
TASK_PP(16'h93A2,4);
TASK_PP(16'h93A3,4);
TASK_PP(16'h93A4,4);
TASK_PP(16'h93A5,4);
TASK_PP(16'h93A6,4);
TASK_PP(16'h93A7,4);
TASK_PP(16'h93A8,4);
TASK_PP(16'h93A9,4);
TASK_PP(16'h93AA,4);
TASK_PP(16'h93AB,4);
TASK_PP(16'h93AC,4);
TASK_PP(16'h93AD,4);
TASK_PP(16'h93AE,4);
TASK_PP(16'h93AF,4);
TASK_PP(16'h93B0,4);
TASK_PP(16'h93B1,4);
TASK_PP(16'h93B2,4);
TASK_PP(16'h93B3,4);
TASK_PP(16'h93B4,4);
TASK_PP(16'h93B5,4);
TASK_PP(16'h93B6,4);
TASK_PP(16'h93B7,4);
TASK_PP(16'h93B8,4);
TASK_PP(16'h93B9,4);
TASK_PP(16'h93BA,4);
TASK_PP(16'h93BB,4);
TASK_PP(16'h93BC,4);
TASK_PP(16'h93BD,4);
TASK_PP(16'h93BE,4);
TASK_PP(16'h93BF,4);
TASK_PP(16'h93C0,4);
TASK_PP(16'h93C1,4);
TASK_PP(16'h93C2,4);
TASK_PP(16'h93C3,4);
TASK_PP(16'h93C4,4);
TASK_PP(16'h93C5,4);
TASK_PP(16'h93C6,4);
TASK_PP(16'h93C7,4);
TASK_PP(16'h93C8,4);
TASK_PP(16'h93C9,4);
TASK_PP(16'h93CA,4);
TASK_PP(16'h93CB,4);
TASK_PP(16'h93CC,4);
TASK_PP(16'h93CD,4);
TASK_PP(16'h93CE,4);
TASK_PP(16'h93CF,4);
TASK_PP(16'h93D0,4);
TASK_PP(16'h93D1,4);
TASK_PP(16'h93D2,4);
TASK_PP(16'h93D3,4);
TASK_PP(16'h93D4,4);
TASK_PP(16'h93D5,4);
TASK_PP(16'h93D6,4);
TASK_PP(16'h93D7,4);
TASK_PP(16'h93D8,4);
TASK_PP(16'h93D9,4);
TASK_PP(16'h93DA,4);
TASK_PP(16'h93DB,4);
TASK_PP(16'h93DC,4);
TASK_PP(16'h93DD,4);
TASK_PP(16'h93DE,4);
TASK_PP(16'h93DF,4);
TASK_PP(16'h93E0,4);
TASK_PP(16'h93E1,4);
TASK_PP(16'h93E2,4);
TASK_PP(16'h93E3,4);
TASK_PP(16'h93E4,4);
TASK_PP(16'h93E5,4);
TASK_PP(16'h93E6,4);
TASK_PP(16'h93E7,4);
TASK_PP(16'h93E8,4);
TASK_PP(16'h93E9,4);
TASK_PP(16'h93EA,4);
TASK_PP(16'h93EB,4);
TASK_PP(16'h93EC,4);
TASK_PP(16'h93ED,4);
TASK_PP(16'h93EE,4);
TASK_PP(16'h93EF,4);
TASK_PP(16'h93F0,4);
TASK_PP(16'h93F1,4);
TASK_PP(16'h93F2,4);
TASK_PP(16'h93F3,4);
TASK_PP(16'h93F4,4);
TASK_PP(16'h93F5,4);
TASK_PP(16'h93F6,4);
TASK_PP(16'h93F7,4);
TASK_PP(16'h93F8,4);
TASK_PP(16'h93F9,4);
TASK_PP(16'h93FA,4);
TASK_PP(16'h93FB,4);
TASK_PP(16'h93FC,4);
TASK_PP(16'h93FD,4);
TASK_PP(16'h93FE,4);
TASK_PP(16'h93FF,4);
TASK_PP(16'h9400,4);
TASK_PP(16'h9401,4);
TASK_PP(16'h9402,4);
TASK_PP(16'h9403,4);
TASK_PP(16'h9404,4);
TASK_PP(16'h9405,4);
TASK_PP(16'h9406,4);
TASK_PP(16'h9407,4);
TASK_PP(16'h9408,4);
TASK_PP(16'h9409,4);
TASK_PP(16'h940A,4);
TASK_PP(16'h940B,4);
TASK_PP(16'h940C,4);
TASK_PP(16'h940D,4);
TASK_PP(16'h940E,4);
TASK_PP(16'h940F,4);
TASK_PP(16'h9410,4);
TASK_PP(16'h9411,4);
TASK_PP(16'h9412,4);
TASK_PP(16'h9413,4);
TASK_PP(16'h9414,4);
TASK_PP(16'h9415,4);
TASK_PP(16'h9416,4);
TASK_PP(16'h9417,4);
TASK_PP(16'h9418,4);
TASK_PP(16'h9419,4);
TASK_PP(16'h941A,4);
TASK_PP(16'h941B,4);
TASK_PP(16'h941C,4);
TASK_PP(16'h941D,4);
TASK_PP(16'h941E,4);
TASK_PP(16'h941F,4);
TASK_PP(16'h9420,4);
TASK_PP(16'h9421,4);
TASK_PP(16'h9422,4);
TASK_PP(16'h9423,4);
TASK_PP(16'h9424,4);
TASK_PP(16'h9425,4);
TASK_PP(16'h9426,4);
TASK_PP(16'h9427,4);
TASK_PP(16'h9428,4);
TASK_PP(16'h9429,4);
TASK_PP(16'h942A,4);
TASK_PP(16'h942B,4);
TASK_PP(16'h942C,4);
TASK_PP(16'h942D,4);
TASK_PP(16'h942E,4);
TASK_PP(16'h942F,4);
TASK_PP(16'h9430,4);
TASK_PP(16'h9431,4);
TASK_PP(16'h9432,4);
TASK_PP(16'h9433,4);
TASK_PP(16'h9434,4);
TASK_PP(16'h9435,4);
TASK_PP(16'h9436,4);
TASK_PP(16'h9437,4);
TASK_PP(16'h9438,4);
TASK_PP(16'h9439,4);
TASK_PP(16'h943A,4);
TASK_PP(16'h943B,4);
TASK_PP(16'h943C,4);
TASK_PP(16'h943D,4);
TASK_PP(16'h943E,4);
TASK_PP(16'h943F,4);
TASK_PP(16'h9440,4);
TASK_PP(16'h9441,4);
TASK_PP(16'h9442,4);
TASK_PP(16'h9443,4);
TASK_PP(16'h9444,4);
TASK_PP(16'h9445,4);
TASK_PP(16'h9446,4);
TASK_PP(16'h9447,4);
TASK_PP(16'h9448,4);
TASK_PP(16'h9449,4);
TASK_PP(16'h944A,4);
TASK_PP(16'h944B,4);
TASK_PP(16'h944C,4);
TASK_PP(16'h944D,4);
TASK_PP(16'h944E,4);
TASK_PP(16'h944F,4);
TASK_PP(16'h9450,4);
TASK_PP(16'h9451,4);
TASK_PP(16'h9452,4);
TASK_PP(16'h9453,4);
TASK_PP(16'h9454,4);
TASK_PP(16'h9455,4);
TASK_PP(16'h9456,4);
TASK_PP(16'h9457,4);
TASK_PP(16'h9458,4);
TASK_PP(16'h9459,4);
TASK_PP(16'h945A,4);
TASK_PP(16'h945B,4);
TASK_PP(16'h945C,4);
TASK_PP(16'h945D,4);
TASK_PP(16'h945E,4);
TASK_PP(16'h945F,4);
TASK_PP(16'h9460,4);
TASK_PP(16'h9461,4);
TASK_PP(16'h9462,4);
TASK_PP(16'h9463,4);
TASK_PP(16'h9464,4);
TASK_PP(16'h9465,4);
TASK_PP(16'h9466,4);
TASK_PP(16'h9467,4);
TASK_PP(16'h9468,4);
TASK_PP(16'h9469,4);
TASK_PP(16'h946A,4);
TASK_PP(16'h946B,4);
TASK_PP(16'h946C,4);
TASK_PP(16'h946D,4);
TASK_PP(16'h946E,4);
TASK_PP(16'h946F,4);
TASK_PP(16'h9470,4);
TASK_PP(16'h9471,4);
TASK_PP(16'h9472,4);
TASK_PP(16'h9473,4);
TASK_PP(16'h9474,4);
TASK_PP(16'h9475,4);
TASK_PP(16'h9476,4);
TASK_PP(16'h9477,4);
TASK_PP(16'h9478,4);
TASK_PP(16'h9479,4);
TASK_PP(16'h947A,4);
TASK_PP(16'h947B,4);
TASK_PP(16'h947C,4);
TASK_PP(16'h947D,4);
TASK_PP(16'h947E,4);
TASK_PP(16'h947F,4);
TASK_PP(16'h9480,4);
TASK_PP(16'h9481,4);
TASK_PP(16'h9482,4);
TASK_PP(16'h9483,4);
TASK_PP(16'h9484,4);
TASK_PP(16'h9485,4);
TASK_PP(16'h9486,4);
TASK_PP(16'h9487,4);
TASK_PP(16'h9488,4);
TASK_PP(16'h9489,4);
TASK_PP(16'h948A,4);
TASK_PP(16'h948B,4);
TASK_PP(16'h948C,4);
TASK_PP(16'h948D,4);
TASK_PP(16'h948E,4);
TASK_PP(16'h948F,4);
TASK_PP(16'h9490,4);
TASK_PP(16'h9491,4);
TASK_PP(16'h9492,4);
TASK_PP(16'h9493,4);
TASK_PP(16'h9494,4);
TASK_PP(16'h9495,4);
TASK_PP(16'h9496,4);
TASK_PP(16'h9497,4);
TASK_PP(16'h9498,4);
TASK_PP(16'h9499,4);
TASK_PP(16'h949A,4);
TASK_PP(16'h949B,4);
TASK_PP(16'h949C,4);
TASK_PP(16'h949D,4);
TASK_PP(16'h949E,4);
TASK_PP(16'h949F,4);
TASK_PP(16'h94A0,4);
TASK_PP(16'h94A1,4);
TASK_PP(16'h94A2,4);
TASK_PP(16'h94A3,4);
TASK_PP(16'h94A4,4);
TASK_PP(16'h94A5,4);
TASK_PP(16'h94A6,4);
TASK_PP(16'h94A7,4);
TASK_PP(16'h94A8,4);
TASK_PP(16'h94A9,4);
TASK_PP(16'h94AA,4);
TASK_PP(16'h94AB,4);
TASK_PP(16'h94AC,4);
TASK_PP(16'h94AD,4);
TASK_PP(16'h94AE,4);
TASK_PP(16'h94AF,4);
TASK_PP(16'h94B0,4);
TASK_PP(16'h94B1,4);
TASK_PP(16'h94B2,4);
TASK_PP(16'h94B3,4);
TASK_PP(16'h94B4,4);
TASK_PP(16'h94B5,4);
TASK_PP(16'h94B6,4);
TASK_PP(16'h94B7,4);
TASK_PP(16'h94B8,4);
TASK_PP(16'h94B9,4);
TASK_PP(16'h94BA,4);
TASK_PP(16'h94BB,4);
TASK_PP(16'h94BC,4);
TASK_PP(16'h94BD,4);
TASK_PP(16'h94BE,4);
TASK_PP(16'h94BF,4);
TASK_PP(16'h94C0,4);
TASK_PP(16'h94C1,4);
TASK_PP(16'h94C2,4);
TASK_PP(16'h94C3,4);
TASK_PP(16'h94C4,4);
TASK_PP(16'h94C5,4);
TASK_PP(16'h94C6,4);
TASK_PP(16'h94C7,4);
TASK_PP(16'h94C8,4);
TASK_PP(16'h94C9,4);
TASK_PP(16'h94CA,4);
TASK_PP(16'h94CB,4);
TASK_PP(16'h94CC,4);
TASK_PP(16'h94CD,4);
TASK_PP(16'h94CE,4);
TASK_PP(16'h94CF,4);
TASK_PP(16'h94D0,4);
TASK_PP(16'h94D1,4);
TASK_PP(16'h94D2,4);
TASK_PP(16'h94D3,4);
TASK_PP(16'h94D4,4);
TASK_PP(16'h94D5,4);
TASK_PP(16'h94D6,4);
TASK_PP(16'h94D7,4);
TASK_PP(16'h94D8,4);
TASK_PP(16'h94D9,4);
TASK_PP(16'h94DA,4);
TASK_PP(16'h94DB,4);
TASK_PP(16'h94DC,4);
TASK_PP(16'h94DD,4);
TASK_PP(16'h94DE,4);
TASK_PP(16'h94DF,4);
TASK_PP(16'h94E0,4);
TASK_PP(16'h94E1,4);
TASK_PP(16'h94E2,4);
TASK_PP(16'h94E3,4);
TASK_PP(16'h94E4,4);
TASK_PP(16'h94E5,4);
TASK_PP(16'h94E6,4);
TASK_PP(16'h94E7,4);
TASK_PP(16'h94E8,4);
TASK_PP(16'h94E9,4);
TASK_PP(16'h94EA,4);
TASK_PP(16'h94EB,4);
TASK_PP(16'h94EC,4);
TASK_PP(16'h94ED,4);
TASK_PP(16'h94EE,4);
TASK_PP(16'h94EF,4);
TASK_PP(16'h94F0,4);
TASK_PP(16'h94F1,4);
TASK_PP(16'h94F2,4);
TASK_PP(16'h94F3,4);
TASK_PP(16'h94F4,4);
TASK_PP(16'h94F5,4);
TASK_PP(16'h94F6,4);
TASK_PP(16'h94F7,4);
TASK_PP(16'h94F8,4);
TASK_PP(16'h94F9,4);
TASK_PP(16'h94FA,4);
TASK_PP(16'h94FB,4);
TASK_PP(16'h94FC,4);
TASK_PP(16'h94FD,4);
TASK_PP(16'h94FE,4);
TASK_PP(16'h94FF,4);
TASK_PP(16'h9500,4);
TASK_PP(16'h9501,4);
TASK_PP(16'h9502,4);
TASK_PP(16'h9503,4);
TASK_PP(16'h9504,4);
TASK_PP(16'h9505,4);
TASK_PP(16'h9506,4);
TASK_PP(16'h9507,4);
TASK_PP(16'h9508,4);
TASK_PP(16'h9509,4);
TASK_PP(16'h950A,4);
TASK_PP(16'h950B,4);
TASK_PP(16'h950C,4);
TASK_PP(16'h950D,4);
TASK_PP(16'h950E,4);
TASK_PP(16'h950F,4);
TASK_PP(16'h9510,4);
TASK_PP(16'h9511,4);
TASK_PP(16'h9512,4);
TASK_PP(16'h9513,4);
TASK_PP(16'h9514,4);
TASK_PP(16'h9515,4);
TASK_PP(16'h9516,4);
TASK_PP(16'h9517,4);
TASK_PP(16'h9518,4);
TASK_PP(16'h9519,4);
TASK_PP(16'h951A,4);
TASK_PP(16'h951B,4);
TASK_PP(16'h951C,4);
TASK_PP(16'h951D,4);
TASK_PP(16'h951E,4);
TASK_PP(16'h951F,4);
TASK_PP(16'h9520,4);
TASK_PP(16'h9521,4);
TASK_PP(16'h9522,4);
TASK_PP(16'h9523,4);
TASK_PP(16'h9524,4);
TASK_PP(16'h9525,4);
TASK_PP(16'h9526,4);
TASK_PP(16'h9527,4);
TASK_PP(16'h9528,4);
TASK_PP(16'h9529,4);
TASK_PP(16'h952A,4);
TASK_PP(16'h952B,4);
TASK_PP(16'h952C,4);
TASK_PP(16'h952D,4);
TASK_PP(16'h952E,4);
TASK_PP(16'h952F,4);
TASK_PP(16'h9530,4);
TASK_PP(16'h9531,4);
TASK_PP(16'h9532,4);
TASK_PP(16'h9533,4);
TASK_PP(16'h9534,4);
TASK_PP(16'h9535,4);
TASK_PP(16'h9536,4);
TASK_PP(16'h9537,4);
TASK_PP(16'h9538,4);
TASK_PP(16'h9539,4);
TASK_PP(16'h953A,4);
TASK_PP(16'h953B,4);
TASK_PP(16'h953C,4);
TASK_PP(16'h953D,4);
TASK_PP(16'h953E,4);
TASK_PP(16'h953F,4);
TASK_PP(16'h9540,4);
TASK_PP(16'h9541,4);
TASK_PP(16'h9542,4);
TASK_PP(16'h9543,4);
TASK_PP(16'h9544,4);
TASK_PP(16'h9545,4);
TASK_PP(16'h9546,4);
TASK_PP(16'h9547,4);
TASK_PP(16'h9548,4);
TASK_PP(16'h9549,4);
TASK_PP(16'h954A,4);
TASK_PP(16'h954B,4);
TASK_PP(16'h954C,4);
TASK_PP(16'h954D,4);
TASK_PP(16'h954E,4);
TASK_PP(16'h954F,4);
TASK_PP(16'h9550,4);
TASK_PP(16'h9551,4);
TASK_PP(16'h9552,4);
TASK_PP(16'h9553,4);
TASK_PP(16'h9554,4);
TASK_PP(16'h9555,4);
TASK_PP(16'h9556,4);
TASK_PP(16'h9557,4);
TASK_PP(16'h9558,4);
TASK_PP(16'h9559,4);
TASK_PP(16'h955A,4);
TASK_PP(16'h955B,4);
TASK_PP(16'h955C,4);
TASK_PP(16'h955D,4);
TASK_PP(16'h955E,4);
TASK_PP(16'h955F,4);
TASK_PP(16'h9560,4);
TASK_PP(16'h9561,4);
TASK_PP(16'h9562,4);
TASK_PP(16'h9563,4);
TASK_PP(16'h9564,4);
TASK_PP(16'h9565,4);
TASK_PP(16'h9566,4);
TASK_PP(16'h9567,4);
TASK_PP(16'h9568,4);
TASK_PP(16'h9569,4);
TASK_PP(16'h956A,4);
TASK_PP(16'h956B,4);
TASK_PP(16'h956C,4);
TASK_PP(16'h956D,4);
TASK_PP(16'h956E,4);
TASK_PP(16'h956F,4);
TASK_PP(16'h9570,4);
TASK_PP(16'h9571,4);
TASK_PP(16'h9572,4);
TASK_PP(16'h9573,4);
TASK_PP(16'h9574,4);
TASK_PP(16'h9575,4);
TASK_PP(16'h9576,4);
TASK_PP(16'h9577,4);
TASK_PP(16'h9578,4);
TASK_PP(16'h9579,4);
TASK_PP(16'h957A,4);
TASK_PP(16'h957B,4);
TASK_PP(16'h957C,4);
TASK_PP(16'h957D,4);
TASK_PP(16'h957E,4);
TASK_PP(16'h957F,4);
TASK_PP(16'h9580,4);
TASK_PP(16'h9581,4);
TASK_PP(16'h9582,4);
TASK_PP(16'h9583,4);
TASK_PP(16'h9584,4);
TASK_PP(16'h9585,4);
TASK_PP(16'h9586,4);
TASK_PP(16'h9587,4);
TASK_PP(16'h9588,4);
TASK_PP(16'h9589,4);
TASK_PP(16'h958A,4);
TASK_PP(16'h958B,4);
TASK_PP(16'h958C,4);
TASK_PP(16'h958D,4);
TASK_PP(16'h958E,4);
TASK_PP(16'h958F,4);
TASK_PP(16'h9590,4);
TASK_PP(16'h9591,4);
TASK_PP(16'h9592,4);
TASK_PP(16'h9593,4);
TASK_PP(16'h9594,4);
TASK_PP(16'h9595,4);
TASK_PP(16'h9596,4);
TASK_PP(16'h9597,4);
TASK_PP(16'h9598,4);
TASK_PP(16'h9599,4);
TASK_PP(16'h959A,4);
TASK_PP(16'h959B,4);
TASK_PP(16'h959C,4);
TASK_PP(16'h959D,4);
TASK_PP(16'h959E,4);
TASK_PP(16'h959F,4);
TASK_PP(16'h95A0,4);
TASK_PP(16'h95A1,4);
TASK_PP(16'h95A2,4);
TASK_PP(16'h95A3,4);
TASK_PP(16'h95A4,4);
TASK_PP(16'h95A5,4);
TASK_PP(16'h95A6,4);
TASK_PP(16'h95A7,4);
TASK_PP(16'h95A8,4);
TASK_PP(16'h95A9,4);
TASK_PP(16'h95AA,4);
TASK_PP(16'h95AB,4);
TASK_PP(16'h95AC,4);
TASK_PP(16'h95AD,4);
TASK_PP(16'h95AE,4);
TASK_PP(16'h95AF,4);
TASK_PP(16'h95B0,4);
TASK_PP(16'h95B1,4);
TASK_PP(16'h95B2,4);
TASK_PP(16'h95B3,4);
TASK_PP(16'h95B4,4);
TASK_PP(16'h95B5,4);
TASK_PP(16'h95B6,4);
TASK_PP(16'h95B7,4);
TASK_PP(16'h95B8,4);
TASK_PP(16'h95B9,4);
TASK_PP(16'h95BA,4);
TASK_PP(16'h95BB,4);
TASK_PP(16'h95BC,4);
TASK_PP(16'h95BD,4);
TASK_PP(16'h95BE,4);
TASK_PP(16'h95BF,4);
TASK_PP(16'h95C0,4);
TASK_PP(16'h95C1,4);
TASK_PP(16'h95C2,4);
TASK_PP(16'h95C3,4);
TASK_PP(16'h95C4,4);
TASK_PP(16'h95C5,4);
TASK_PP(16'h95C6,4);
TASK_PP(16'h95C7,4);
TASK_PP(16'h95C8,4);
TASK_PP(16'h95C9,4);
TASK_PP(16'h95CA,4);
TASK_PP(16'h95CB,4);
TASK_PP(16'h95CC,4);
TASK_PP(16'h95CD,4);
TASK_PP(16'h95CE,4);
TASK_PP(16'h95CF,4);
TASK_PP(16'h95D0,4);
TASK_PP(16'h95D1,4);
TASK_PP(16'h95D2,4);
TASK_PP(16'h95D3,4);
TASK_PP(16'h95D4,4);
TASK_PP(16'h95D5,4);
TASK_PP(16'h95D6,4);
TASK_PP(16'h95D7,4);
TASK_PP(16'h95D8,4);
TASK_PP(16'h95D9,4);
TASK_PP(16'h95DA,4);
TASK_PP(16'h95DB,4);
TASK_PP(16'h95DC,4);
TASK_PP(16'h95DD,4);
TASK_PP(16'h95DE,4);
TASK_PP(16'h95DF,4);
TASK_PP(16'h95E0,4);
TASK_PP(16'h95E1,4);
TASK_PP(16'h95E2,4);
TASK_PP(16'h95E3,4);
TASK_PP(16'h95E4,4);
TASK_PP(16'h95E5,4);
TASK_PP(16'h95E6,4);
TASK_PP(16'h95E7,4);
TASK_PP(16'h95E8,4);
TASK_PP(16'h95E9,4);
TASK_PP(16'h95EA,4);
TASK_PP(16'h95EB,4);
TASK_PP(16'h95EC,4);
TASK_PP(16'h95ED,4);
TASK_PP(16'h95EE,4);
TASK_PP(16'h95EF,4);
TASK_PP(16'h95F0,4);
TASK_PP(16'h95F1,4);
TASK_PP(16'h95F2,4);
TASK_PP(16'h95F3,4);
TASK_PP(16'h95F4,4);
TASK_PP(16'h95F5,4);
TASK_PP(16'h95F6,4);
TASK_PP(16'h95F7,4);
TASK_PP(16'h95F8,4);
TASK_PP(16'h95F9,4);
TASK_PP(16'h95FA,4);
TASK_PP(16'h95FB,4);
TASK_PP(16'h95FC,4);
TASK_PP(16'h95FD,4);
TASK_PP(16'h95FE,4);
TASK_PP(16'h95FF,4);
TASK_PP(16'h9600,4);
TASK_PP(16'h9601,4);
TASK_PP(16'h9602,4);
TASK_PP(16'h9603,4);
TASK_PP(16'h9604,4);
TASK_PP(16'h9605,4);
TASK_PP(16'h9606,4);
TASK_PP(16'h9607,4);
TASK_PP(16'h9608,4);
TASK_PP(16'h9609,4);
TASK_PP(16'h960A,4);
TASK_PP(16'h960B,4);
TASK_PP(16'h960C,4);
TASK_PP(16'h960D,4);
TASK_PP(16'h960E,4);
TASK_PP(16'h960F,4);
TASK_PP(16'h9610,4);
TASK_PP(16'h9611,4);
TASK_PP(16'h9612,4);
TASK_PP(16'h9613,4);
TASK_PP(16'h9614,4);
TASK_PP(16'h9615,4);
TASK_PP(16'h9616,4);
TASK_PP(16'h9617,4);
TASK_PP(16'h9618,4);
TASK_PP(16'h9619,4);
TASK_PP(16'h961A,4);
TASK_PP(16'h961B,4);
TASK_PP(16'h961C,4);
TASK_PP(16'h961D,4);
TASK_PP(16'h961E,4);
TASK_PP(16'h961F,4);
TASK_PP(16'h9620,4);
TASK_PP(16'h9621,4);
TASK_PP(16'h9622,4);
TASK_PP(16'h9623,4);
TASK_PP(16'h9624,4);
TASK_PP(16'h9625,4);
TASK_PP(16'h9626,4);
TASK_PP(16'h9627,4);
TASK_PP(16'h9628,4);
TASK_PP(16'h9629,4);
TASK_PP(16'h962A,4);
TASK_PP(16'h962B,4);
TASK_PP(16'h962C,4);
TASK_PP(16'h962D,4);
TASK_PP(16'h962E,4);
TASK_PP(16'h962F,4);
TASK_PP(16'h9630,4);
TASK_PP(16'h9631,4);
TASK_PP(16'h9632,4);
TASK_PP(16'h9633,4);
TASK_PP(16'h9634,4);
TASK_PP(16'h9635,4);
TASK_PP(16'h9636,4);
TASK_PP(16'h9637,4);
TASK_PP(16'h9638,4);
TASK_PP(16'h9639,4);
TASK_PP(16'h963A,4);
TASK_PP(16'h963B,4);
TASK_PP(16'h963C,4);
TASK_PP(16'h963D,4);
TASK_PP(16'h963E,4);
TASK_PP(16'h963F,4);
TASK_PP(16'h9640,4);
TASK_PP(16'h9641,4);
TASK_PP(16'h9642,4);
TASK_PP(16'h9643,4);
TASK_PP(16'h9644,4);
TASK_PP(16'h9645,4);
TASK_PP(16'h9646,4);
TASK_PP(16'h9647,4);
TASK_PP(16'h9648,4);
TASK_PP(16'h9649,4);
TASK_PP(16'h964A,4);
TASK_PP(16'h964B,4);
TASK_PP(16'h964C,4);
TASK_PP(16'h964D,4);
TASK_PP(16'h964E,4);
TASK_PP(16'h964F,4);
TASK_PP(16'h9650,4);
TASK_PP(16'h9651,4);
TASK_PP(16'h9652,4);
TASK_PP(16'h9653,4);
TASK_PP(16'h9654,4);
TASK_PP(16'h9655,4);
TASK_PP(16'h9656,4);
TASK_PP(16'h9657,4);
TASK_PP(16'h9658,4);
TASK_PP(16'h9659,4);
TASK_PP(16'h965A,4);
TASK_PP(16'h965B,4);
TASK_PP(16'h965C,4);
TASK_PP(16'h965D,4);
TASK_PP(16'h965E,4);
TASK_PP(16'h965F,4);
TASK_PP(16'h9660,4);
TASK_PP(16'h9661,4);
TASK_PP(16'h9662,4);
TASK_PP(16'h9663,4);
TASK_PP(16'h9664,4);
TASK_PP(16'h9665,4);
TASK_PP(16'h9666,4);
TASK_PP(16'h9667,4);
TASK_PP(16'h9668,4);
TASK_PP(16'h9669,4);
TASK_PP(16'h966A,4);
TASK_PP(16'h966B,4);
TASK_PP(16'h966C,4);
TASK_PP(16'h966D,4);
TASK_PP(16'h966E,4);
TASK_PP(16'h966F,4);
TASK_PP(16'h9670,4);
TASK_PP(16'h9671,4);
TASK_PP(16'h9672,4);
TASK_PP(16'h9673,4);
TASK_PP(16'h9674,4);
TASK_PP(16'h9675,4);
TASK_PP(16'h9676,4);
TASK_PP(16'h9677,4);
TASK_PP(16'h9678,4);
TASK_PP(16'h9679,4);
TASK_PP(16'h967A,4);
TASK_PP(16'h967B,4);
TASK_PP(16'h967C,4);
TASK_PP(16'h967D,4);
TASK_PP(16'h967E,4);
TASK_PP(16'h967F,4);
TASK_PP(16'h9680,4);
TASK_PP(16'h9681,4);
TASK_PP(16'h9682,4);
TASK_PP(16'h9683,4);
TASK_PP(16'h9684,4);
TASK_PP(16'h9685,4);
TASK_PP(16'h9686,4);
TASK_PP(16'h9687,4);
TASK_PP(16'h9688,4);
TASK_PP(16'h9689,4);
TASK_PP(16'h968A,4);
TASK_PP(16'h968B,4);
TASK_PP(16'h968C,4);
TASK_PP(16'h968D,4);
TASK_PP(16'h968E,4);
TASK_PP(16'h968F,4);
TASK_PP(16'h9690,4);
TASK_PP(16'h9691,4);
TASK_PP(16'h9692,4);
TASK_PP(16'h9693,4);
TASK_PP(16'h9694,4);
TASK_PP(16'h9695,4);
TASK_PP(16'h9696,4);
TASK_PP(16'h9697,4);
TASK_PP(16'h9698,4);
TASK_PP(16'h9699,4);
TASK_PP(16'h969A,4);
TASK_PP(16'h969B,4);
TASK_PP(16'h969C,4);
TASK_PP(16'h969D,4);
TASK_PP(16'h969E,4);
TASK_PP(16'h969F,4);
TASK_PP(16'h96A0,4);
TASK_PP(16'h96A1,4);
TASK_PP(16'h96A2,4);
TASK_PP(16'h96A3,4);
TASK_PP(16'h96A4,4);
TASK_PP(16'h96A5,4);
TASK_PP(16'h96A6,4);
TASK_PP(16'h96A7,4);
TASK_PP(16'h96A8,4);
TASK_PP(16'h96A9,4);
TASK_PP(16'h96AA,4);
TASK_PP(16'h96AB,4);
TASK_PP(16'h96AC,4);
TASK_PP(16'h96AD,4);
TASK_PP(16'h96AE,4);
TASK_PP(16'h96AF,4);
TASK_PP(16'h96B0,4);
TASK_PP(16'h96B1,4);
TASK_PP(16'h96B2,4);
TASK_PP(16'h96B3,4);
TASK_PP(16'h96B4,4);
TASK_PP(16'h96B5,4);
TASK_PP(16'h96B6,4);
TASK_PP(16'h96B7,4);
TASK_PP(16'h96B8,4);
TASK_PP(16'h96B9,4);
TASK_PP(16'h96BA,4);
TASK_PP(16'h96BB,4);
TASK_PP(16'h96BC,4);
TASK_PP(16'h96BD,4);
TASK_PP(16'h96BE,4);
TASK_PP(16'h96BF,4);
TASK_PP(16'h96C0,4);
TASK_PP(16'h96C1,4);
TASK_PP(16'h96C2,4);
TASK_PP(16'h96C3,4);
TASK_PP(16'h96C4,4);
TASK_PP(16'h96C5,4);
TASK_PP(16'h96C6,4);
TASK_PP(16'h96C7,4);
TASK_PP(16'h96C8,4);
TASK_PP(16'h96C9,4);
TASK_PP(16'h96CA,4);
TASK_PP(16'h96CB,4);
TASK_PP(16'h96CC,4);
TASK_PP(16'h96CD,4);
TASK_PP(16'h96CE,4);
TASK_PP(16'h96CF,4);
TASK_PP(16'h96D0,4);
TASK_PP(16'h96D1,4);
TASK_PP(16'h96D2,4);
TASK_PP(16'h96D3,4);
TASK_PP(16'h96D4,4);
TASK_PP(16'h96D5,4);
TASK_PP(16'h96D6,4);
TASK_PP(16'h96D7,4);
TASK_PP(16'h96D8,4);
TASK_PP(16'h96D9,4);
TASK_PP(16'h96DA,4);
TASK_PP(16'h96DB,4);
TASK_PP(16'h96DC,4);
TASK_PP(16'h96DD,4);
TASK_PP(16'h96DE,4);
TASK_PP(16'h96DF,4);
TASK_PP(16'h96E0,4);
TASK_PP(16'h96E1,4);
TASK_PP(16'h96E2,4);
TASK_PP(16'h96E3,4);
TASK_PP(16'h96E4,4);
TASK_PP(16'h96E5,4);
TASK_PP(16'h96E6,4);
TASK_PP(16'h96E7,4);
TASK_PP(16'h96E8,4);
TASK_PP(16'h96E9,4);
TASK_PP(16'h96EA,4);
TASK_PP(16'h96EB,4);
TASK_PP(16'h96EC,4);
TASK_PP(16'h96ED,4);
TASK_PP(16'h96EE,4);
TASK_PP(16'h96EF,4);
TASK_PP(16'h96F0,4);
TASK_PP(16'h96F1,4);
TASK_PP(16'h96F2,4);
TASK_PP(16'h96F3,4);
TASK_PP(16'h96F4,4);
TASK_PP(16'h96F5,4);
TASK_PP(16'h96F6,4);
TASK_PP(16'h96F7,4);
TASK_PP(16'h96F8,4);
TASK_PP(16'h96F9,4);
TASK_PP(16'h96FA,4);
TASK_PP(16'h96FB,4);
TASK_PP(16'h96FC,4);
TASK_PP(16'h96FD,4);
TASK_PP(16'h96FE,4);
TASK_PP(16'h96FF,4);
TASK_PP(16'h9700,4);
TASK_PP(16'h9701,4);
TASK_PP(16'h9702,4);
TASK_PP(16'h9703,4);
TASK_PP(16'h9704,4);
TASK_PP(16'h9705,4);
TASK_PP(16'h9706,4);
TASK_PP(16'h9707,4);
TASK_PP(16'h9708,4);
TASK_PP(16'h9709,4);
TASK_PP(16'h970A,4);
TASK_PP(16'h970B,4);
TASK_PP(16'h970C,4);
TASK_PP(16'h970D,4);
TASK_PP(16'h970E,4);
TASK_PP(16'h970F,4);
TASK_PP(16'h9710,4);
TASK_PP(16'h9711,4);
TASK_PP(16'h9712,4);
TASK_PP(16'h9713,4);
TASK_PP(16'h9714,4);
TASK_PP(16'h9715,4);
TASK_PP(16'h9716,4);
TASK_PP(16'h9717,4);
TASK_PP(16'h9718,4);
TASK_PP(16'h9719,4);
TASK_PP(16'h971A,4);
TASK_PP(16'h971B,4);
TASK_PP(16'h971C,4);
TASK_PP(16'h971D,4);
TASK_PP(16'h971E,4);
TASK_PP(16'h971F,4);
TASK_PP(16'h9720,4);
TASK_PP(16'h9721,4);
TASK_PP(16'h9722,4);
TASK_PP(16'h9723,4);
TASK_PP(16'h9724,4);
TASK_PP(16'h9725,4);
TASK_PP(16'h9726,4);
TASK_PP(16'h9727,4);
TASK_PP(16'h9728,4);
TASK_PP(16'h9729,4);
TASK_PP(16'h972A,4);
TASK_PP(16'h972B,4);
TASK_PP(16'h972C,4);
TASK_PP(16'h972D,4);
TASK_PP(16'h972E,4);
TASK_PP(16'h972F,4);
TASK_PP(16'h9730,4);
TASK_PP(16'h9731,4);
TASK_PP(16'h9732,4);
TASK_PP(16'h9733,4);
TASK_PP(16'h9734,4);
TASK_PP(16'h9735,4);
TASK_PP(16'h9736,4);
TASK_PP(16'h9737,4);
TASK_PP(16'h9738,4);
TASK_PP(16'h9739,4);
TASK_PP(16'h973A,4);
TASK_PP(16'h973B,4);
TASK_PP(16'h973C,4);
TASK_PP(16'h973D,4);
TASK_PP(16'h973E,4);
TASK_PP(16'h973F,4);
TASK_PP(16'h9740,4);
TASK_PP(16'h9741,4);
TASK_PP(16'h9742,4);
TASK_PP(16'h9743,4);
TASK_PP(16'h9744,4);
TASK_PP(16'h9745,4);
TASK_PP(16'h9746,4);
TASK_PP(16'h9747,4);
TASK_PP(16'h9748,4);
TASK_PP(16'h9749,4);
TASK_PP(16'h974A,4);
TASK_PP(16'h974B,4);
TASK_PP(16'h974C,4);
TASK_PP(16'h974D,4);
TASK_PP(16'h974E,4);
TASK_PP(16'h974F,4);
TASK_PP(16'h9750,4);
TASK_PP(16'h9751,4);
TASK_PP(16'h9752,4);
TASK_PP(16'h9753,4);
TASK_PP(16'h9754,4);
TASK_PP(16'h9755,4);
TASK_PP(16'h9756,4);
TASK_PP(16'h9757,4);
TASK_PP(16'h9758,4);
TASK_PP(16'h9759,4);
TASK_PP(16'h975A,4);
TASK_PP(16'h975B,4);
TASK_PP(16'h975C,4);
TASK_PP(16'h975D,4);
TASK_PP(16'h975E,4);
TASK_PP(16'h975F,4);
TASK_PP(16'h9760,4);
TASK_PP(16'h9761,4);
TASK_PP(16'h9762,4);
TASK_PP(16'h9763,4);
TASK_PP(16'h9764,4);
TASK_PP(16'h9765,4);
TASK_PP(16'h9766,4);
TASK_PP(16'h9767,4);
TASK_PP(16'h9768,4);
TASK_PP(16'h9769,4);
TASK_PP(16'h976A,4);
TASK_PP(16'h976B,4);
TASK_PP(16'h976C,4);
TASK_PP(16'h976D,4);
TASK_PP(16'h976E,4);
TASK_PP(16'h976F,4);
TASK_PP(16'h9770,4);
TASK_PP(16'h9771,4);
TASK_PP(16'h9772,4);
TASK_PP(16'h9773,4);
TASK_PP(16'h9774,4);
TASK_PP(16'h9775,4);
TASK_PP(16'h9776,4);
TASK_PP(16'h9777,4);
TASK_PP(16'h9778,4);
TASK_PP(16'h9779,4);
TASK_PP(16'h977A,4);
TASK_PP(16'h977B,4);
TASK_PP(16'h977C,4);
TASK_PP(16'h977D,4);
TASK_PP(16'h977E,4);
TASK_PP(16'h977F,4);
TASK_PP(16'h9780,4);
TASK_PP(16'h9781,4);
TASK_PP(16'h9782,4);
TASK_PP(16'h9783,4);
TASK_PP(16'h9784,4);
TASK_PP(16'h9785,4);
TASK_PP(16'h9786,4);
TASK_PP(16'h9787,4);
TASK_PP(16'h9788,4);
TASK_PP(16'h9789,4);
TASK_PP(16'h978A,4);
TASK_PP(16'h978B,4);
TASK_PP(16'h978C,4);
TASK_PP(16'h978D,4);
TASK_PP(16'h978E,4);
TASK_PP(16'h978F,4);
TASK_PP(16'h9790,4);
TASK_PP(16'h9791,4);
TASK_PP(16'h9792,4);
TASK_PP(16'h9793,4);
TASK_PP(16'h9794,4);
TASK_PP(16'h9795,4);
TASK_PP(16'h9796,4);
TASK_PP(16'h9797,4);
TASK_PP(16'h9798,4);
TASK_PP(16'h9799,4);
TASK_PP(16'h979A,4);
TASK_PP(16'h979B,4);
TASK_PP(16'h979C,4);
TASK_PP(16'h979D,4);
TASK_PP(16'h979E,4);
TASK_PP(16'h979F,4);
TASK_PP(16'h97A0,4);
TASK_PP(16'h97A1,4);
TASK_PP(16'h97A2,4);
TASK_PP(16'h97A3,4);
TASK_PP(16'h97A4,4);
TASK_PP(16'h97A5,4);
TASK_PP(16'h97A6,4);
TASK_PP(16'h97A7,4);
TASK_PP(16'h97A8,4);
TASK_PP(16'h97A9,4);
TASK_PP(16'h97AA,4);
TASK_PP(16'h97AB,4);
TASK_PP(16'h97AC,4);
TASK_PP(16'h97AD,4);
TASK_PP(16'h97AE,4);
TASK_PP(16'h97AF,4);
TASK_PP(16'h97B0,4);
TASK_PP(16'h97B1,4);
TASK_PP(16'h97B2,4);
TASK_PP(16'h97B3,4);
TASK_PP(16'h97B4,4);
TASK_PP(16'h97B5,4);
TASK_PP(16'h97B6,4);
TASK_PP(16'h97B7,4);
TASK_PP(16'h97B8,4);
TASK_PP(16'h97B9,4);
TASK_PP(16'h97BA,4);
TASK_PP(16'h97BB,4);
TASK_PP(16'h97BC,4);
TASK_PP(16'h97BD,4);
TASK_PP(16'h97BE,4);
TASK_PP(16'h97BF,4);
TASK_PP(16'h97C0,4);
TASK_PP(16'h97C1,4);
TASK_PP(16'h97C2,4);
TASK_PP(16'h97C3,4);
TASK_PP(16'h97C4,4);
TASK_PP(16'h97C5,4);
TASK_PP(16'h97C6,4);
TASK_PP(16'h97C7,4);
TASK_PP(16'h97C8,4);
TASK_PP(16'h97C9,4);
TASK_PP(16'h97CA,4);
TASK_PP(16'h97CB,4);
TASK_PP(16'h97CC,4);
TASK_PP(16'h97CD,4);
TASK_PP(16'h97CE,4);
TASK_PP(16'h97CF,4);
TASK_PP(16'h97D0,4);
TASK_PP(16'h97D1,4);
TASK_PP(16'h97D2,4);
TASK_PP(16'h97D3,4);
TASK_PP(16'h97D4,4);
TASK_PP(16'h97D5,4);
TASK_PP(16'h97D6,4);
TASK_PP(16'h97D7,4);
TASK_PP(16'h97D8,4);
TASK_PP(16'h97D9,4);
TASK_PP(16'h97DA,4);
TASK_PP(16'h97DB,4);
TASK_PP(16'h97DC,4);
TASK_PP(16'h97DD,4);
TASK_PP(16'h97DE,4);
TASK_PP(16'h97DF,4);
TASK_PP(16'h97E0,4);
TASK_PP(16'h97E1,4);
TASK_PP(16'h97E2,4);
TASK_PP(16'h97E3,4);
TASK_PP(16'h97E4,4);
TASK_PP(16'h97E5,4);
TASK_PP(16'h97E6,4);
TASK_PP(16'h97E7,4);
TASK_PP(16'h97E8,4);
TASK_PP(16'h97E9,4);
TASK_PP(16'h97EA,4);
TASK_PP(16'h97EB,4);
TASK_PP(16'h97EC,4);
TASK_PP(16'h97ED,4);
TASK_PP(16'h97EE,4);
TASK_PP(16'h97EF,4);
TASK_PP(16'h97F0,4);
TASK_PP(16'h97F1,4);
TASK_PP(16'h97F2,4);
TASK_PP(16'h97F3,4);
TASK_PP(16'h97F4,4);
TASK_PP(16'h97F5,4);
TASK_PP(16'h97F6,4);
TASK_PP(16'h97F7,4);
TASK_PP(16'h97F8,4);
TASK_PP(16'h97F9,4);
TASK_PP(16'h97FA,4);
TASK_PP(16'h97FB,4);
TASK_PP(16'h97FC,4);
TASK_PP(16'h97FD,4);
TASK_PP(16'h97FE,4);
TASK_PP(16'h97FF,4);
TASK_PP(16'h9800,4);
TASK_PP(16'h9801,4);
TASK_PP(16'h9802,4);
TASK_PP(16'h9803,4);
TASK_PP(16'h9804,4);
TASK_PP(16'h9805,4);
TASK_PP(16'h9806,4);
TASK_PP(16'h9807,4);
TASK_PP(16'h9808,4);
TASK_PP(16'h9809,4);
TASK_PP(16'h980A,4);
TASK_PP(16'h980B,4);
TASK_PP(16'h980C,4);
TASK_PP(16'h980D,4);
TASK_PP(16'h980E,4);
TASK_PP(16'h980F,4);
TASK_PP(16'h9810,4);
TASK_PP(16'h9811,4);
TASK_PP(16'h9812,4);
TASK_PP(16'h9813,4);
TASK_PP(16'h9814,4);
TASK_PP(16'h9815,4);
TASK_PP(16'h9816,4);
TASK_PP(16'h9817,4);
TASK_PP(16'h9818,4);
TASK_PP(16'h9819,4);
TASK_PP(16'h981A,4);
TASK_PP(16'h981B,4);
TASK_PP(16'h981C,4);
TASK_PP(16'h981D,4);
TASK_PP(16'h981E,4);
TASK_PP(16'h981F,4);
TASK_PP(16'h9820,4);
TASK_PP(16'h9821,4);
TASK_PP(16'h9822,4);
TASK_PP(16'h9823,4);
TASK_PP(16'h9824,4);
TASK_PP(16'h9825,4);
TASK_PP(16'h9826,4);
TASK_PP(16'h9827,4);
TASK_PP(16'h9828,4);
TASK_PP(16'h9829,4);
TASK_PP(16'h982A,4);
TASK_PP(16'h982B,4);
TASK_PP(16'h982C,4);
TASK_PP(16'h982D,4);
TASK_PP(16'h982E,4);
TASK_PP(16'h982F,4);
TASK_PP(16'h9830,4);
TASK_PP(16'h9831,4);
TASK_PP(16'h9832,4);
TASK_PP(16'h9833,4);
TASK_PP(16'h9834,4);
TASK_PP(16'h9835,4);
TASK_PP(16'h9836,4);
TASK_PP(16'h9837,4);
TASK_PP(16'h9838,4);
TASK_PP(16'h9839,4);
TASK_PP(16'h983A,4);
TASK_PP(16'h983B,4);
TASK_PP(16'h983C,4);
TASK_PP(16'h983D,4);
TASK_PP(16'h983E,4);
TASK_PP(16'h983F,4);
TASK_PP(16'h9840,4);
TASK_PP(16'h9841,4);
TASK_PP(16'h9842,4);
TASK_PP(16'h9843,4);
TASK_PP(16'h9844,4);
TASK_PP(16'h9845,4);
TASK_PP(16'h9846,4);
TASK_PP(16'h9847,4);
TASK_PP(16'h9848,4);
TASK_PP(16'h9849,4);
TASK_PP(16'h984A,4);
TASK_PP(16'h984B,4);
TASK_PP(16'h984C,4);
TASK_PP(16'h984D,4);
TASK_PP(16'h984E,4);
TASK_PP(16'h984F,4);
TASK_PP(16'h9850,4);
TASK_PP(16'h9851,4);
TASK_PP(16'h9852,4);
TASK_PP(16'h9853,4);
TASK_PP(16'h9854,4);
TASK_PP(16'h9855,4);
TASK_PP(16'h9856,4);
TASK_PP(16'h9857,4);
TASK_PP(16'h9858,4);
TASK_PP(16'h9859,4);
TASK_PP(16'h985A,4);
TASK_PP(16'h985B,4);
TASK_PP(16'h985C,4);
TASK_PP(16'h985D,4);
TASK_PP(16'h985E,4);
TASK_PP(16'h985F,4);
TASK_PP(16'h9860,4);
TASK_PP(16'h9861,4);
TASK_PP(16'h9862,4);
TASK_PP(16'h9863,4);
TASK_PP(16'h9864,4);
TASK_PP(16'h9865,4);
TASK_PP(16'h9866,4);
TASK_PP(16'h9867,4);
TASK_PP(16'h9868,4);
TASK_PP(16'h9869,4);
TASK_PP(16'h986A,4);
TASK_PP(16'h986B,4);
TASK_PP(16'h986C,4);
TASK_PP(16'h986D,4);
TASK_PP(16'h986E,4);
TASK_PP(16'h986F,4);
TASK_PP(16'h9870,4);
TASK_PP(16'h9871,4);
TASK_PP(16'h9872,4);
TASK_PP(16'h9873,4);
TASK_PP(16'h9874,4);
TASK_PP(16'h9875,4);
TASK_PP(16'h9876,4);
TASK_PP(16'h9877,4);
TASK_PP(16'h9878,4);
TASK_PP(16'h9879,4);
TASK_PP(16'h987A,4);
TASK_PP(16'h987B,4);
TASK_PP(16'h987C,4);
TASK_PP(16'h987D,4);
TASK_PP(16'h987E,4);
TASK_PP(16'h987F,4);
TASK_PP(16'h9880,4);
TASK_PP(16'h9881,4);
TASK_PP(16'h9882,4);
TASK_PP(16'h9883,4);
TASK_PP(16'h9884,4);
TASK_PP(16'h9885,4);
TASK_PP(16'h9886,4);
TASK_PP(16'h9887,4);
TASK_PP(16'h9888,4);
TASK_PP(16'h9889,4);
TASK_PP(16'h988A,4);
TASK_PP(16'h988B,4);
TASK_PP(16'h988C,4);
TASK_PP(16'h988D,4);
TASK_PP(16'h988E,4);
TASK_PP(16'h988F,4);
TASK_PP(16'h9890,4);
TASK_PP(16'h9891,4);
TASK_PP(16'h9892,4);
TASK_PP(16'h9893,4);
TASK_PP(16'h9894,4);
TASK_PP(16'h9895,4);
TASK_PP(16'h9896,4);
TASK_PP(16'h9897,4);
TASK_PP(16'h9898,4);
TASK_PP(16'h9899,4);
TASK_PP(16'h989A,4);
TASK_PP(16'h989B,4);
TASK_PP(16'h989C,4);
TASK_PP(16'h989D,4);
TASK_PP(16'h989E,4);
TASK_PP(16'h989F,4);
TASK_PP(16'h98A0,4);
TASK_PP(16'h98A1,4);
TASK_PP(16'h98A2,4);
TASK_PP(16'h98A3,4);
TASK_PP(16'h98A4,4);
TASK_PP(16'h98A5,4);
TASK_PP(16'h98A6,4);
TASK_PP(16'h98A7,4);
TASK_PP(16'h98A8,4);
TASK_PP(16'h98A9,4);
TASK_PP(16'h98AA,4);
TASK_PP(16'h98AB,4);
TASK_PP(16'h98AC,4);
TASK_PP(16'h98AD,4);
TASK_PP(16'h98AE,4);
TASK_PP(16'h98AF,4);
TASK_PP(16'h98B0,4);
TASK_PP(16'h98B1,4);
TASK_PP(16'h98B2,4);
TASK_PP(16'h98B3,4);
TASK_PP(16'h98B4,4);
TASK_PP(16'h98B5,4);
TASK_PP(16'h98B6,4);
TASK_PP(16'h98B7,4);
TASK_PP(16'h98B8,4);
TASK_PP(16'h98B9,4);
TASK_PP(16'h98BA,4);
TASK_PP(16'h98BB,4);
TASK_PP(16'h98BC,4);
TASK_PP(16'h98BD,4);
TASK_PP(16'h98BE,4);
TASK_PP(16'h98BF,4);
TASK_PP(16'h98C0,4);
TASK_PP(16'h98C1,4);
TASK_PP(16'h98C2,4);
TASK_PP(16'h98C3,4);
TASK_PP(16'h98C4,4);
TASK_PP(16'h98C5,4);
TASK_PP(16'h98C6,4);
TASK_PP(16'h98C7,4);
TASK_PP(16'h98C8,4);
TASK_PP(16'h98C9,4);
TASK_PP(16'h98CA,4);
TASK_PP(16'h98CB,4);
TASK_PP(16'h98CC,4);
TASK_PP(16'h98CD,4);
TASK_PP(16'h98CE,4);
TASK_PP(16'h98CF,4);
TASK_PP(16'h98D0,4);
TASK_PP(16'h98D1,4);
TASK_PP(16'h98D2,4);
TASK_PP(16'h98D3,4);
TASK_PP(16'h98D4,4);
TASK_PP(16'h98D5,4);
TASK_PP(16'h98D6,4);
TASK_PP(16'h98D7,4);
TASK_PP(16'h98D8,4);
TASK_PP(16'h98D9,4);
TASK_PP(16'h98DA,4);
TASK_PP(16'h98DB,4);
TASK_PP(16'h98DC,4);
TASK_PP(16'h98DD,4);
TASK_PP(16'h98DE,4);
TASK_PP(16'h98DF,4);
TASK_PP(16'h98E0,4);
TASK_PP(16'h98E1,4);
TASK_PP(16'h98E2,4);
TASK_PP(16'h98E3,4);
TASK_PP(16'h98E4,4);
TASK_PP(16'h98E5,4);
TASK_PP(16'h98E6,4);
TASK_PP(16'h98E7,4);
TASK_PP(16'h98E8,4);
TASK_PP(16'h98E9,4);
TASK_PP(16'h98EA,4);
TASK_PP(16'h98EB,4);
TASK_PP(16'h98EC,4);
TASK_PP(16'h98ED,4);
TASK_PP(16'h98EE,4);
TASK_PP(16'h98EF,4);
TASK_PP(16'h98F0,4);
TASK_PP(16'h98F1,4);
TASK_PP(16'h98F2,4);
TASK_PP(16'h98F3,4);
TASK_PP(16'h98F4,4);
TASK_PP(16'h98F5,4);
TASK_PP(16'h98F6,4);
TASK_PP(16'h98F7,4);
TASK_PP(16'h98F8,4);
TASK_PP(16'h98F9,4);
TASK_PP(16'h98FA,4);
TASK_PP(16'h98FB,4);
TASK_PP(16'h98FC,4);
TASK_PP(16'h98FD,4);
TASK_PP(16'h98FE,4);
TASK_PP(16'h98FF,4);
TASK_PP(16'h9900,4);
TASK_PP(16'h9901,4);
TASK_PP(16'h9902,4);
TASK_PP(16'h9903,4);
TASK_PP(16'h9904,4);
TASK_PP(16'h9905,4);
TASK_PP(16'h9906,4);
TASK_PP(16'h9907,4);
TASK_PP(16'h9908,4);
TASK_PP(16'h9909,4);
TASK_PP(16'h990A,4);
TASK_PP(16'h990B,4);
TASK_PP(16'h990C,4);
TASK_PP(16'h990D,4);
TASK_PP(16'h990E,4);
TASK_PP(16'h990F,4);
TASK_PP(16'h9910,4);
TASK_PP(16'h9911,4);
TASK_PP(16'h9912,4);
TASK_PP(16'h9913,4);
TASK_PP(16'h9914,4);
TASK_PP(16'h9915,4);
TASK_PP(16'h9916,4);
TASK_PP(16'h9917,4);
TASK_PP(16'h9918,4);
TASK_PP(16'h9919,4);
TASK_PP(16'h991A,4);
TASK_PP(16'h991B,4);
TASK_PP(16'h991C,4);
TASK_PP(16'h991D,4);
TASK_PP(16'h991E,4);
TASK_PP(16'h991F,4);
TASK_PP(16'h9920,4);
TASK_PP(16'h9921,4);
TASK_PP(16'h9922,4);
TASK_PP(16'h9923,4);
TASK_PP(16'h9924,4);
TASK_PP(16'h9925,4);
TASK_PP(16'h9926,4);
TASK_PP(16'h9927,4);
TASK_PP(16'h9928,4);
TASK_PP(16'h9929,4);
TASK_PP(16'h992A,4);
TASK_PP(16'h992B,4);
TASK_PP(16'h992C,4);
TASK_PP(16'h992D,4);
TASK_PP(16'h992E,4);
TASK_PP(16'h992F,4);
TASK_PP(16'h9930,4);
TASK_PP(16'h9931,4);
TASK_PP(16'h9932,4);
TASK_PP(16'h9933,4);
TASK_PP(16'h9934,4);
TASK_PP(16'h9935,4);
TASK_PP(16'h9936,4);
TASK_PP(16'h9937,4);
TASK_PP(16'h9938,4);
TASK_PP(16'h9939,4);
TASK_PP(16'h993A,4);
TASK_PP(16'h993B,4);
TASK_PP(16'h993C,4);
TASK_PP(16'h993D,4);
TASK_PP(16'h993E,4);
TASK_PP(16'h993F,4);
TASK_PP(16'h9940,4);
TASK_PP(16'h9941,4);
TASK_PP(16'h9942,4);
TASK_PP(16'h9943,4);
TASK_PP(16'h9944,4);
TASK_PP(16'h9945,4);
TASK_PP(16'h9946,4);
TASK_PP(16'h9947,4);
TASK_PP(16'h9948,4);
TASK_PP(16'h9949,4);
TASK_PP(16'h994A,4);
TASK_PP(16'h994B,4);
TASK_PP(16'h994C,4);
TASK_PP(16'h994D,4);
TASK_PP(16'h994E,4);
TASK_PP(16'h994F,4);
TASK_PP(16'h9950,4);
TASK_PP(16'h9951,4);
TASK_PP(16'h9952,4);
TASK_PP(16'h9953,4);
TASK_PP(16'h9954,4);
TASK_PP(16'h9955,4);
TASK_PP(16'h9956,4);
TASK_PP(16'h9957,4);
TASK_PP(16'h9958,4);
TASK_PP(16'h9959,4);
TASK_PP(16'h995A,4);
TASK_PP(16'h995B,4);
TASK_PP(16'h995C,4);
TASK_PP(16'h995D,4);
TASK_PP(16'h995E,4);
TASK_PP(16'h995F,4);
TASK_PP(16'h9960,4);
TASK_PP(16'h9961,4);
TASK_PP(16'h9962,4);
TASK_PP(16'h9963,4);
TASK_PP(16'h9964,4);
TASK_PP(16'h9965,4);
TASK_PP(16'h9966,4);
TASK_PP(16'h9967,4);
TASK_PP(16'h9968,4);
TASK_PP(16'h9969,4);
TASK_PP(16'h996A,4);
TASK_PP(16'h996B,4);
TASK_PP(16'h996C,4);
TASK_PP(16'h996D,4);
TASK_PP(16'h996E,4);
TASK_PP(16'h996F,4);
TASK_PP(16'h9970,4);
TASK_PP(16'h9971,4);
TASK_PP(16'h9972,4);
TASK_PP(16'h9973,4);
TASK_PP(16'h9974,4);
TASK_PP(16'h9975,4);
TASK_PP(16'h9976,4);
TASK_PP(16'h9977,4);
TASK_PP(16'h9978,4);
TASK_PP(16'h9979,4);
TASK_PP(16'h997A,4);
TASK_PP(16'h997B,4);
TASK_PP(16'h997C,4);
TASK_PP(16'h997D,4);
TASK_PP(16'h997E,4);
TASK_PP(16'h997F,4);
TASK_PP(16'h9980,4);
TASK_PP(16'h9981,4);
TASK_PP(16'h9982,4);
TASK_PP(16'h9983,4);
TASK_PP(16'h9984,4);
TASK_PP(16'h9985,4);
TASK_PP(16'h9986,4);
TASK_PP(16'h9987,4);
TASK_PP(16'h9988,4);
TASK_PP(16'h9989,4);
TASK_PP(16'h998A,4);
TASK_PP(16'h998B,4);
TASK_PP(16'h998C,4);
TASK_PP(16'h998D,4);
TASK_PP(16'h998E,4);
TASK_PP(16'h998F,4);
TASK_PP(16'h9990,4);
TASK_PP(16'h9991,4);
TASK_PP(16'h9992,4);
TASK_PP(16'h9993,4);
TASK_PP(16'h9994,4);
TASK_PP(16'h9995,4);
TASK_PP(16'h9996,4);
TASK_PP(16'h9997,4);
TASK_PP(16'h9998,4);
TASK_PP(16'h9999,4);
TASK_PP(16'h999A,4);
TASK_PP(16'h999B,4);
TASK_PP(16'h999C,4);
TASK_PP(16'h999D,4);
TASK_PP(16'h999E,4);
TASK_PP(16'h999F,4);
TASK_PP(16'h99A0,4);
TASK_PP(16'h99A1,4);
TASK_PP(16'h99A2,4);
TASK_PP(16'h99A3,4);
TASK_PP(16'h99A4,4);
TASK_PP(16'h99A5,4);
TASK_PP(16'h99A6,4);
TASK_PP(16'h99A7,4);
TASK_PP(16'h99A8,4);
TASK_PP(16'h99A9,4);
TASK_PP(16'h99AA,4);
TASK_PP(16'h99AB,4);
TASK_PP(16'h99AC,4);
TASK_PP(16'h99AD,4);
TASK_PP(16'h99AE,4);
TASK_PP(16'h99AF,4);
TASK_PP(16'h99B0,4);
TASK_PP(16'h99B1,4);
TASK_PP(16'h99B2,4);
TASK_PP(16'h99B3,4);
TASK_PP(16'h99B4,4);
TASK_PP(16'h99B5,4);
TASK_PP(16'h99B6,4);
TASK_PP(16'h99B7,4);
TASK_PP(16'h99B8,4);
TASK_PP(16'h99B9,4);
TASK_PP(16'h99BA,4);
TASK_PP(16'h99BB,4);
TASK_PP(16'h99BC,4);
TASK_PP(16'h99BD,4);
TASK_PP(16'h99BE,4);
TASK_PP(16'h99BF,4);
TASK_PP(16'h99C0,4);
TASK_PP(16'h99C1,4);
TASK_PP(16'h99C2,4);
TASK_PP(16'h99C3,4);
TASK_PP(16'h99C4,4);
TASK_PP(16'h99C5,4);
TASK_PP(16'h99C6,4);
TASK_PP(16'h99C7,4);
TASK_PP(16'h99C8,4);
TASK_PP(16'h99C9,4);
TASK_PP(16'h99CA,4);
TASK_PP(16'h99CB,4);
TASK_PP(16'h99CC,4);
TASK_PP(16'h99CD,4);
TASK_PP(16'h99CE,4);
TASK_PP(16'h99CF,4);
TASK_PP(16'h99D0,4);
TASK_PP(16'h99D1,4);
TASK_PP(16'h99D2,4);
TASK_PP(16'h99D3,4);
TASK_PP(16'h99D4,4);
TASK_PP(16'h99D5,4);
TASK_PP(16'h99D6,4);
TASK_PP(16'h99D7,4);
TASK_PP(16'h99D8,4);
TASK_PP(16'h99D9,4);
TASK_PP(16'h99DA,4);
TASK_PP(16'h99DB,4);
TASK_PP(16'h99DC,4);
TASK_PP(16'h99DD,4);
TASK_PP(16'h99DE,4);
TASK_PP(16'h99DF,4);
TASK_PP(16'h99E0,4);
TASK_PP(16'h99E1,4);
TASK_PP(16'h99E2,4);
TASK_PP(16'h99E3,4);
TASK_PP(16'h99E4,4);
TASK_PP(16'h99E5,4);
TASK_PP(16'h99E6,4);
TASK_PP(16'h99E7,4);
TASK_PP(16'h99E8,4);
TASK_PP(16'h99E9,4);
TASK_PP(16'h99EA,4);
TASK_PP(16'h99EB,4);
TASK_PP(16'h99EC,4);
TASK_PP(16'h99ED,4);
TASK_PP(16'h99EE,4);
TASK_PP(16'h99EF,4);
TASK_PP(16'h99F0,4);
TASK_PP(16'h99F1,4);
TASK_PP(16'h99F2,4);
TASK_PP(16'h99F3,4);
TASK_PP(16'h99F4,4);
TASK_PP(16'h99F5,4);
TASK_PP(16'h99F6,4);
TASK_PP(16'h99F7,4);
TASK_PP(16'h99F8,4);
TASK_PP(16'h99F9,4);
TASK_PP(16'h99FA,4);
TASK_PP(16'h99FB,4);
TASK_PP(16'h99FC,4);
TASK_PP(16'h99FD,4);
TASK_PP(16'h99FE,4);
TASK_PP(16'h99FF,4);
TASK_PP(16'h9A00,4);
TASK_PP(16'h9A01,4);
TASK_PP(16'h9A02,4);
TASK_PP(16'h9A03,4);
TASK_PP(16'h9A04,4);
TASK_PP(16'h9A05,4);
TASK_PP(16'h9A06,4);
TASK_PP(16'h9A07,4);
TASK_PP(16'h9A08,4);
TASK_PP(16'h9A09,4);
TASK_PP(16'h9A0A,4);
TASK_PP(16'h9A0B,4);
TASK_PP(16'h9A0C,4);
TASK_PP(16'h9A0D,4);
TASK_PP(16'h9A0E,4);
TASK_PP(16'h9A0F,4);
TASK_PP(16'h9A10,4);
TASK_PP(16'h9A11,4);
TASK_PP(16'h9A12,4);
TASK_PP(16'h9A13,4);
TASK_PP(16'h9A14,4);
TASK_PP(16'h9A15,4);
TASK_PP(16'h9A16,4);
TASK_PP(16'h9A17,4);
TASK_PP(16'h9A18,4);
TASK_PP(16'h9A19,4);
TASK_PP(16'h9A1A,4);
TASK_PP(16'h9A1B,4);
TASK_PP(16'h9A1C,4);
TASK_PP(16'h9A1D,4);
TASK_PP(16'h9A1E,4);
TASK_PP(16'h9A1F,4);
TASK_PP(16'h9A20,4);
TASK_PP(16'h9A21,4);
TASK_PP(16'h9A22,4);
TASK_PP(16'h9A23,4);
TASK_PP(16'h9A24,4);
TASK_PP(16'h9A25,4);
TASK_PP(16'h9A26,4);
TASK_PP(16'h9A27,4);
TASK_PP(16'h9A28,4);
TASK_PP(16'h9A29,4);
TASK_PP(16'h9A2A,4);
TASK_PP(16'h9A2B,4);
TASK_PP(16'h9A2C,4);
TASK_PP(16'h9A2D,4);
TASK_PP(16'h9A2E,4);
TASK_PP(16'h9A2F,4);
TASK_PP(16'h9A30,4);
TASK_PP(16'h9A31,4);
TASK_PP(16'h9A32,4);
TASK_PP(16'h9A33,4);
TASK_PP(16'h9A34,4);
TASK_PP(16'h9A35,4);
TASK_PP(16'h9A36,4);
TASK_PP(16'h9A37,4);
TASK_PP(16'h9A38,4);
TASK_PP(16'h9A39,4);
TASK_PP(16'h9A3A,4);
TASK_PP(16'h9A3B,4);
TASK_PP(16'h9A3C,4);
TASK_PP(16'h9A3D,4);
TASK_PP(16'h9A3E,4);
TASK_PP(16'h9A3F,4);
TASK_PP(16'h9A40,4);
TASK_PP(16'h9A41,4);
TASK_PP(16'h9A42,4);
TASK_PP(16'h9A43,4);
TASK_PP(16'h9A44,4);
TASK_PP(16'h9A45,4);
TASK_PP(16'h9A46,4);
TASK_PP(16'h9A47,4);
TASK_PP(16'h9A48,4);
TASK_PP(16'h9A49,4);
TASK_PP(16'h9A4A,4);
TASK_PP(16'h9A4B,4);
TASK_PP(16'h9A4C,4);
TASK_PP(16'h9A4D,4);
TASK_PP(16'h9A4E,4);
TASK_PP(16'h9A4F,4);
TASK_PP(16'h9A50,4);
TASK_PP(16'h9A51,4);
TASK_PP(16'h9A52,4);
TASK_PP(16'h9A53,4);
TASK_PP(16'h9A54,4);
TASK_PP(16'h9A55,4);
TASK_PP(16'h9A56,4);
TASK_PP(16'h9A57,4);
TASK_PP(16'h9A58,4);
TASK_PP(16'h9A59,4);
TASK_PP(16'h9A5A,4);
TASK_PP(16'h9A5B,4);
TASK_PP(16'h9A5C,4);
TASK_PP(16'h9A5D,4);
TASK_PP(16'h9A5E,4);
TASK_PP(16'h9A5F,4);
TASK_PP(16'h9A60,4);
TASK_PP(16'h9A61,4);
TASK_PP(16'h9A62,4);
TASK_PP(16'h9A63,4);
TASK_PP(16'h9A64,4);
TASK_PP(16'h9A65,4);
TASK_PP(16'h9A66,4);
TASK_PP(16'h9A67,4);
TASK_PP(16'h9A68,4);
TASK_PP(16'h9A69,4);
TASK_PP(16'h9A6A,4);
TASK_PP(16'h9A6B,4);
TASK_PP(16'h9A6C,4);
TASK_PP(16'h9A6D,4);
TASK_PP(16'h9A6E,4);
TASK_PP(16'h9A6F,4);
TASK_PP(16'h9A70,4);
TASK_PP(16'h9A71,4);
TASK_PP(16'h9A72,4);
TASK_PP(16'h9A73,4);
TASK_PP(16'h9A74,4);
TASK_PP(16'h9A75,4);
TASK_PP(16'h9A76,4);
TASK_PP(16'h9A77,4);
TASK_PP(16'h9A78,4);
TASK_PP(16'h9A79,4);
TASK_PP(16'h9A7A,4);
TASK_PP(16'h9A7B,4);
TASK_PP(16'h9A7C,4);
TASK_PP(16'h9A7D,4);
TASK_PP(16'h9A7E,4);
TASK_PP(16'h9A7F,4);
TASK_PP(16'h9A80,4);
TASK_PP(16'h9A81,4);
TASK_PP(16'h9A82,4);
TASK_PP(16'h9A83,4);
TASK_PP(16'h9A84,4);
TASK_PP(16'h9A85,4);
TASK_PP(16'h9A86,4);
TASK_PP(16'h9A87,4);
TASK_PP(16'h9A88,4);
TASK_PP(16'h9A89,4);
TASK_PP(16'h9A8A,4);
TASK_PP(16'h9A8B,4);
TASK_PP(16'h9A8C,4);
TASK_PP(16'h9A8D,4);
TASK_PP(16'h9A8E,4);
TASK_PP(16'h9A8F,4);
TASK_PP(16'h9A90,4);
TASK_PP(16'h9A91,4);
TASK_PP(16'h9A92,4);
TASK_PP(16'h9A93,4);
TASK_PP(16'h9A94,4);
TASK_PP(16'h9A95,4);
TASK_PP(16'h9A96,4);
TASK_PP(16'h9A97,4);
TASK_PP(16'h9A98,4);
TASK_PP(16'h9A99,4);
TASK_PP(16'h9A9A,4);
TASK_PP(16'h9A9B,4);
TASK_PP(16'h9A9C,4);
TASK_PP(16'h9A9D,4);
TASK_PP(16'h9A9E,4);
TASK_PP(16'h9A9F,4);
TASK_PP(16'h9AA0,4);
TASK_PP(16'h9AA1,4);
TASK_PP(16'h9AA2,4);
TASK_PP(16'h9AA3,4);
TASK_PP(16'h9AA4,4);
TASK_PP(16'h9AA5,4);
TASK_PP(16'h9AA6,4);
TASK_PP(16'h9AA7,4);
TASK_PP(16'h9AA8,4);
TASK_PP(16'h9AA9,4);
TASK_PP(16'h9AAA,4);
TASK_PP(16'h9AAB,4);
TASK_PP(16'h9AAC,4);
TASK_PP(16'h9AAD,4);
TASK_PP(16'h9AAE,4);
TASK_PP(16'h9AAF,4);
TASK_PP(16'h9AB0,4);
TASK_PP(16'h9AB1,4);
TASK_PP(16'h9AB2,4);
TASK_PP(16'h9AB3,4);
TASK_PP(16'h9AB4,4);
TASK_PP(16'h9AB5,4);
TASK_PP(16'h9AB6,4);
TASK_PP(16'h9AB7,4);
TASK_PP(16'h9AB8,4);
TASK_PP(16'h9AB9,4);
TASK_PP(16'h9ABA,4);
TASK_PP(16'h9ABB,4);
TASK_PP(16'h9ABC,4);
TASK_PP(16'h9ABD,4);
TASK_PP(16'h9ABE,4);
TASK_PP(16'h9ABF,4);
TASK_PP(16'h9AC0,4);
TASK_PP(16'h9AC1,4);
TASK_PP(16'h9AC2,4);
TASK_PP(16'h9AC3,4);
TASK_PP(16'h9AC4,4);
TASK_PP(16'h9AC5,4);
TASK_PP(16'h9AC6,4);
TASK_PP(16'h9AC7,4);
TASK_PP(16'h9AC8,4);
TASK_PP(16'h9AC9,4);
TASK_PP(16'h9ACA,4);
TASK_PP(16'h9ACB,4);
TASK_PP(16'h9ACC,4);
TASK_PP(16'h9ACD,4);
TASK_PP(16'h9ACE,4);
TASK_PP(16'h9ACF,4);
TASK_PP(16'h9AD0,4);
TASK_PP(16'h9AD1,4);
TASK_PP(16'h9AD2,4);
TASK_PP(16'h9AD3,4);
TASK_PP(16'h9AD4,4);
TASK_PP(16'h9AD5,4);
TASK_PP(16'h9AD6,4);
TASK_PP(16'h9AD7,4);
TASK_PP(16'h9AD8,4);
TASK_PP(16'h9AD9,4);
TASK_PP(16'h9ADA,4);
TASK_PP(16'h9ADB,4);
TASK_PP(16'h9ADC,4);
TASK_PP(16'h9ADD,4);
TASK_PP(16'h9ADE,4);
TASK_PP(16'h9ADF,4);
TASK_PP(16'h9AE0,4);
TASK_PP(16'h9AE1,4);
TASK_PP(16'h9AE2,4);
TASK_PP(16'h9AE3,4);
TASK_PP(16'h9AE4,4);
TASK_PP(16'h9AE5,4);
TASK_PP(16'h9AE6,4);
TASK_PP(16'h9AE7,4);
TASK_PP(16'h9AE8,4);
TASK_PP(16'h9AE9,4);
TASK_PP(16'h9AEA,4);
TASK_PP(16'h9AEB,4);
TASK_PP(16'h9AEC,4);
TASK_PP(16'h9AED,4);
TASK_PP(16'h9AEE,4);
TASK_PP(16'h9AEF,4);
TASK_PP(16'h9AF0,4);
TASK_PP(16'h9AF1,4);
TASK_PP(16'h9AF2,4);
TASK_PP(16'h9AF3,4);
TASK_PP(16'h9AF4,4);
TASK_PP(16'h9AF5,4);
TASK_PP(16'h9AF6,4);
TASK_PP(16'h9AF7,4);
TASK_PP(16'h9AF8,4);
TASK_PP(16'h9AF9,4);
TASK_PP(16'h9AFA,4);
TASK_PP(16'h9AFB,4);
TASK_PP(16'h9AFC,4);
TASK_PP(16'h9AFD,4);
TASK_PP(16'h9AFE,4);
TASK_PP(16'h9AFF,4);
TASK_PP(16'h9B00,4);
TASK_PP(16'h9B01,4);
TASK_PP(16'h9B02,4);
TASK_PP(16'h9B03,4);
TASK_PP(16'h9B04,4);
TASK_PP(16'h9B05,4);
TASK_PP(16'h9B06,4);
TASK_PP(16'h9B07,4);
TASK_PP(16'h9B08,4);
TASK_PP(16'h9B09,4);
TASK_PP(16'h9B0A,4);
TASK_PP(16'h9B0B,4);
TASK_PP(16'h9B0C,4);
TASK_PP(16'h9B0D,4);
TASK_PP(16'h9B0E,4);
TASK_PP(16'h9B0F,4);
TASK_PP(16'h9B10,4);
TASK_PP(16'h9B11,4);
TASK_PP(16'h9B12,4);
TASK_PP(16'h9B13,4);
TASK_PP(16'h9B14,4);
TASK_PP(16'h9B15,4);
TASK_PP(16'h9B16,4);
TASK_PP(16'h9B17,4);
TASK_PP(16'h9B18,4);
TASK_PP(16'h9B19,4);
TASK_PP(16'h9B1A,4);
TASK_PP(16'h9B1B,4);
TASK_PP(16'h9B1C,4);
TASK_PP(16'h9B1D,4);
TASK_PP(16'h9B1E,4);
TASK_PP(16'h9B1F,4);
TASK_PP(16'h9B20,4);
TASK_PP(16'h9B21,4);
TASK_PP(16'h9B22,4);
TASK_PP(16'h9B23,4);
TASK_PP(16'h9B24,4);
TASK_PP(16'h9B25,4);
TASK_PP(16'h9B26,4);
TASK_PP(16'h9B27,4);
TASK_PP(16'h9B28,4);
TASK_PP(16'h9B29,4);
TASK_PP(16'h9B2A,4);
TASK_PP(16'h9B2B,4);
TASK_PP(16'h9B2C,4);
TASK_PP(16'h9B2D,4);
TASK_PP(16'h9B2E,4);
TASK_PP(16'h9B2F,4);
TASK_PP(16'h9B30,4);
TASK_PP(16'h9B31,4);
TASK_PP(16'h9B32,4);
TASK_PP(16'h9B33,4);
TASK_PP(16'h9B34,4);
TASK_PP(16'h9B35,4);
TASK_PP(16'h9B36,4);
TASK_PP(16'h9B37,4);
TASK_PP(16'h9B38,4);
TASK_PP(16'h9B39,4);
TASK_PP(16'h9B3A,4);
TASK_PP(16'h9B3B,4);
TASK_PP(16'h9B3C,4);
TASK_PP(16'h9B3D,4);
TASK_PP(16'h9B3E,4);
TASK_PP(16'h9B3F,4);
TASK_PP(16'h9B40,4);
TASK_PP(16'h9B41,4);
TASK_PP(16'h9B42,4);
TASK_PP(16'h9B43,4);
TASK_PP(16'h9B44,4);
TASK_PP(16'h9B45,4);
TASK_PP(16'h9B46,4);
TASK_PP(16'h9B47,4);
TASK_PP(16'h9B48,4);
TASK_PP(16'h9B49,4);
TASK_PP(16'h9B4A,4);
TASK_PP(16'h9B4B,4);
TASK_PP(16'h9B4C,4);
TASK_PP(16'h9B4D,4);
TASK_PP(16'h9B4E,4);
TASK_PP(16'h9B4F,4);
TASK_PP(16'h9B50,4);
TASK_PP(16'h9B51,4);
TASK_PP(16'h9B52,4);
TASK_PP(16'h9B53,4);
TASK_PP(16'h9B54,4);
TASK_PP(16'h9B55,4);
TASK_PP(16'h9B56,4);
TASK_PP(16'h9B57,4);
TASK_PP(16'h9B58,4);
TASK_PP(16'h9B59,4);
TASK_PP(16'h9B5A,4);
TASK_PP(16'h9B5B,4);
TASK_PP(16'h9B5C,4);
TASK_PP(16'h9B5D,4);
TASK_PP(16'h9B5E,4);
TASK_PP(16'h9B5F,4);
TASK_PP(16'h9B60,4);
TASK_PP(16'h9B61,4);
TASK_PP(16'h9B62,4);
TASK_PP(16'h9B63,4);
TASK_PP(16'h9B64,4);
TASK_PP(16'h9B65,4);
TASK_PP(16'h9B66,4);
TASK_PP(16'h9B67,4);
TASK_PP(16'h9B68,4);
TASK_PP(16'h9B69,4);
TASK_PP(16'h9B6A,4);
TASK_PP(16'h9B6B,4);
TASK_PP(16'h9B6C,4);
TASK_PP(16'h9B6D,4);
TASK_PP(16'h9B6E,4);
TASK_PP(16'h9B6F,4);
TASK_PP(16'h9B70,4);
TASK_PP(16'h9B71,4);
TASK_PP(16'h9B72,4);
TASK_PP(16'h9B73,4);
TASK_PP(16'h9B74,4);
TASK_PP(16'h9B75,4);
TASK_PP(16'h9B76,4);
TASK_PP(16'h9B77,4);
TASK_PP(16'h9B78,4);
TASK_PP(16'h9B79,4);
TASK_PP(16'h9B7A,4);
TASK_PP(16'h9B7B,4);
TASK_PP(16'h9B7C,4);
TASK_PP(16'h9B7D,4);
TASK_PP(16'h9B7E,4);
TASK_PP(16'h9B7F,4);
TASK_PP(16'h9B80,4);
TASK_PP(16'h9B81,4);
TASK_PP(16'h9B82,4);
TASK_PP(16'h9B83,4);
TASK_PP(16'h9B84,4);
TASK_PP(16'h9B85,4);
TASK_PP(16'h9B86,4);
TASK_PP(16'h9B87,4);
TASK_PP(16'h9B88,4);
TASK_PP(16'h9B89,4);
TASK_PP(16'h9B8A,4);
TASK_PP(16'h9B8B,4);
TASK_PP(16'h9B8C,4);
TASK_PP(16'h9B8D,4);
TASK_PP(16'h9B8E,4);
TASK_PP(16'h9B8F,4);
TASK_PP(16'h9B90,4);
TASK_PP(16'h9B91,4);
TASK_PP(16'h9B92,4);
TASK_PP(16'h9B93,4);
TASK_PP(16'h9B94,4);
TASK_PP(16'h9B95,4);
TASK_PP(16'h9B96,4);
TASK_PP(16'h9B97,4);
TASK_PP(16'h9B98,4);
TASK_PP(16'h9B99,4);
TASK_PP(16'h9B9A,4);
TASK_PP(16'h9B9B,4);
TASK_PP(16'h9B9C,4);
TASK_PP(16'h9B9D,4);
TASK_PP(16'h9B9E,4);
TASK_PP(16'h9B9F,4);
TASK_PP(16'h9BA0,4);
TASK_PP(16'h9BA1,4);
TASK_PP(16'h9BA2,4);
TASK_PP(16'h9BA3,4);
TASK_PP(16'h9BA4,4);
TASK_PP(16'h9BA5,4);
TASK_PP(16'h9BA6,4);
TASK_PP(16'h9BA7,4);
TASK_PP(16'h9BA8,4);
TASK_PP(16'h9BA9,4);
TASK_PP(16'h9BAA,4);
TASK_PP(16'h9BAB,4);
TASK_PP(16'h9BAC,4);
TASK_PP(16'h9BAD,4);
TASK_PP(16'h9BAE,4);
TASK_PP(16'h9BAF,4);
TASK_PP(16'h9BB0,4);
TASK_PP(16'h9BB1,4);
TASK_PP(16'h9BB2,4);
TASK_PP(16'h9BB3,4);
TASK_PP(16'h9BB4,4);
TASK_PP(16'h9BB5,4);
TASK_PP(16'h9BB6,4);
TASK_PP(16'h9BB7,4);
TASK_PP(16'h9BB8,4);
TASK_PP(16'h9BB9,4);
TASK_PP(16'h9BBA,4);
TASK_PP(16'h9BBB,4);
TASK_PP(16'h9BBC,4);
TASK_PP(16'h9BBD,4);
TASK_PP(16'h9BBE,4);
TASK_PP(16'h9BBF,4);
TASK_PP(16'h9BC0,4);
TASK_PP(16'h9BC1,4);
TASK_PP(16'h9BC2,4);
TASK_PP(16'h9BC3,4);
TASK_PP(16'h9BC4,4);
TASK_PP(16'h9BC5,4);
TASK_PP(16'h9BC6,4);
TASK_PP(16'h9BC7,4);
TASK_PP(16'h9BC8,4);
TASK_PP(16'h9BC9,4);
TASK_PP(16'h9BCA,4);
TASK_PP(16'h9BCB,4);
TASK_PP(16'h9BCC,4);
TASK_PP(16'h9BCD,4);
TASK_PP(16'h9BCE,4);
TASK_PP(16'h9BCF,4);
TASK_PP(16'h9BD0,4);
TASK_PP(16'h9BD1,4);
TASK_PP(16'h9BD2,4);
TASK_PP(16'h9BD3,4);
TASK_PP(16'h9BD4,4);
TASK_PP(16'h9BD5,4);
TASK_PP(16'h9BD6,4);
TASK_PP(16'h9BD7,4);
TASK_PP(16'h9BD8,4);
TASK_PP(16'h9BD9,4);
TASK_PP(16'h9BDA,4);
TASK_PP(16'h9BDB,4);
TASK_PP(16'h9BDC,4);
TASK_PP(16'h9BDD,4);
TASK_PP(16'h9BDE,4);
TASK_PP(16'h9BDF,4);
TASK_PP(16'h9BE0,4);
TASK_PP(16'h9BE1,4);
TASK_PP(16'h9BE2,4);
TASK_PP(16'h9BE3,4);
TASK_PP(16'h9BE4,4);
TASK_PP(16'h9BE5,4);
TASK_PP(16'h9BE6,4);
TASK_PP(16'h9BE7,4);
TASK_PP(16'h9BE8,4);
TASK_PP(16'h9BE9,4);
TASK_PP(16'h9BEA,4);
TASK_PP(16'h9BEB,4);
TASK_PP(16'h9BEC,4);
TASK_PP(16'h9BED,4);
TASK_PP(16'h9BEE,4);
TASK_PP(16'h9BEF,4);
TASK_PP(16'h9BF0,4);
TASK_PP(16'h9BF1,4);
TASK_PP(16'h9BF2,4);
TASK_PP(16'h9BF3,4);
TASK_PP(16'h9BF4,4);
TASK_PP(16'h9BF5,4);
TASK_PP(16'h9BF6,4);
TASK_PP(16'h9BF7,4);
TASK_PP(16'h9BF8,4);
TASK_PP(16'h9BF9,4);
TASK_PP(16'h9BFA,4);
TASK_PP(16'h9BFB,4);
TASK_PP(16'h9BFC,4);
TASK_PP(16'h9BFD,4);
TASK_PP(16'h9BFE,4);
TASK_PP(16'h9BFF,4);
TASK_PP(16'h9C00,4);
TASK_PP(16'h9C01,4);
TASK_PP(16'h9C02,4);
TASK_PP(16'h9C03,4);
TASK_PP(16'h9C04,4);
TASK_PP(16'h9C05,4);
TASK_PP(16'h9C06,4);
TASK_PP(16'h9C07,4);
TASK_PP(16'h9C08,4);
TASK_PP(16'h9C09,4);
TASK_PP(16'h9C0A,4);
TASK_PP(16'h9C0B,4);
TASK_PP(16'h9C0C,4);
TASK_PP(16'h9C0D,4);
TASK_PP(16'h9C0E,4);
TASK_PP(16'h9C0F,4);
TASK_PP(16'h9C10,4);
TASK_PP(16'h9C11,4);
TASK_PP(16'h9C12,4);
TASK_PP(16'h9C13,4);
TASK_PP(16'h9C14,4);
TASK_PP(16'h9C15,4);
TASK_PP(16'h9C16,4);
TASK_PP(16'h9C17,4);
TASK_PP(16'h9C18,4);
TASK_PP(16'h9C19,4);
TASK_PP(16'h9C1A,4);
TASK_PP(16'h9C1B,4);
TASK_PP(16'h9C1C,4);
TASK_PP(16'h9C1D,4);
TASK_PP(16'h9C1E,4);
TASK_PP(16'h9C1F,4);
TASK_PP(16'h9C20,4);
TASK_PP(16'h9C21,4);
TASK_PP(16'h9C22,4);
TASK_PP(16'h9C23,4);
TASK_PP(16'h9C24,4);
TASK_PP(16'h9C25,4);
TASK_PP(16'h9C26,4);
TASK_PP(16'h9C27,4);
TASK_PP(16'h9C28,4);
TASK_PP(16'h9C29,4);
TASK_PP(16'h9C2A,4);
TASK_PP(16'h9C2B,4);
TASK_PP(16'h9C2C,4);
TASK_PP(16'h9C2D,4);
TASK_PP(16'h9C2E,4);
TASK_PP(16'h9C2F,4);
TASK_PP(16'h9C30,4);
TASK_PP(16'h9C31,4);
TASK_PP(16'h9C32,4);
TASK_PP(16'h9C33,4);
TASK_PP(16'h9C34,4);
TASK_PP(16'h9C35,4);
TASK_PP(16'h9C36,4);
TASK_PP(16'h9C37,4);
TASK_PP(16'h9C38,4);
TASK_PP(16'h9C39,4);
TASK_PP(16'h9C3A,4);
TASK_PP(16'h9C3B,4);
TASK_PP(16'h9C3C,4);
TASK_PP(16'h9C3D,4);
TASK_PP(16'h9C3E,4);
TASK_PP(16'h9C3F,4);
TASK_PP(16'h9C40,4);
TASK_PP(16'h9C41,4);
TASK_PP(16'h9C42,4);
TASK_PP(16'h9C43,4);
TASK_PP(16'h9C44,4);
TASK_PP(16'h9C45,4);
TASK_PP(16'h9C46,4);
TASK_PP(16'h9C47,4);
TASK_PP(16'h9C48,4);
TASK_PP(16'h9C49,4);
TASK_PP(16'h9C4A,4);
TASK_PP(16'h9C4B,4);
TASK_PP(16'h9C4C,4);
TASK_PP(16'h9C4D,4);
TASK_PP(16'h9C4E,4);
TASK_PP(16'h9C4F,4);
TASK_PP(16'h9C50,4);
TASK_PP(16'h9C51,4);
TASK_PP(16'h9C52,4);
TASK_PP(16'h9C53,4);
TASK_PP(16'h9C54,4);
TASK_PP(16'h9C55,4);
TASK_PP(16'h9C56,4);
TASK_PP(16'h9C57,4);
TASK_PP(16'h9C58,4);
TASK_PP(16'h9C59,4);
TASK_PP(16'h9C5A,4);
TASK_PP(16'h9C5B,4);
TASK_PP(16'h9C5C,4);
TASK_PP(16'h9C5D,4);
TASK_PP(16'h9C5E,4);
TASK_PP(16'h9C5F,4);
TASK_PP(16'h9C60,4);
TASK_PP(16'h9C61,4);
TASK_PP(16'h9C62,4);
TASK_PP(16'h9C63,4);
TASK_PP(16'h9C64,4);
TASK_PP(16'h9C65,4);
TASK_PP(16'h9C66,4);
TASK_PP(16'h9C67,4);
TASK_PP(16'h9C68,4);
TASK_PP(16'h9C69,4);
TASK_PP(16'h9C6A,4);
TASK_PP(16'h9C6B,4);
TASK_PP(16'h9C6C,4);
TASK_PP(16'h9C6D,4);
TASK_PP(16'h9C6E,4);
TASK_PP(16'h9C6F,4);
TASK_PP(16'h9C70,4);
TASK_PP(16'h9C71,4);
TASK_PP(16'h9C72,4);
TASK_PP(16'h9C73,4);
TASK_PP(16'h9C74,4);
TASK_PP(16'h9C75,4);
TASK_PP(16'h9C76,4);
TASK_PP(16'h9C77,4);
TASK_PP(16'h9C78,4);
TASK_PP(16'h9C79,4);
TASK_PP(16'h9C7A,4);
TASK_PP(16'h9C7B,4);
TASK_PP(16'h9C7C,4);
TASK_PP(16'h9C7D,4);
TASK_PP(16'h9C7E,4);
TASK_PP(16'h9C7F,4);
TASK_PP(16'h9C80,4);
TASK_PP(16'h9C81,4);
TASK_PP(16'h9C82,4);
TASK_PP(16'h9C83,4);
TASK_PP(16'h9C84,4);
TASK_PP(16'h9C85,4);
TASK_PP(16'h9C86,4);
TASK_PP(16'h9C87,4);
TASK_PP(16'h9C88,4);
TASK_PP(16'h9C89,4);
TASK_PP(16'h9C8A,4);
TASK_PP(16'h9C8B,4);
TASK_PP(16'h9C8C,4);
TASK_PP(16'h9C8D,4);
TASK_PP(16'h9C8E,4);
TASK_PP(16'h9C8F,4);
TASK_PP(16'h9C90,4);
TASK_PP(16'h9C91,4);
TASK_PP(16'h9C92,4);
TASK_PP(16'h9C93,4);
TASK_PP(16'h9C94,4);
TASK_PP(16'h9C95,4);
TASK_PP(16'h9C96,4);
TASK_PP(16'h9C97,4);
TASK_PP(16'h9C98,4);
TASK_PP(16'h9C99,4);
TASK_PP(16'h9C9A,4);
TASK_PP(16'h9C9B,4);
TASK_PP(16'h9C9C,4);
TASK_PP(16'h9C9D,4);
TASK_PP(16'h9C9E,4);
TASK_PP(16'h9C9F,4);
TASK_PP(16'h9CA0,4);
TASK_PP(16'h9CA1,4);
TASK_PP(16'h9CA2,4);
TASK_PP(16'h9CA3,4);
TASK_PP(16'h9CA4,4);
TASK_PP(16'h9CA5,4);
TASK_PP(16'h9CA6,4);
TASK_PP(16'h9CA7,4);
TASK_PP(16'h9CA8,4);
TASK_PP(16'h9CA9,4);
TASK_PP(16'h9CAA,4);
TASK_PP(16'h9CAB,4);
TASK_PP(16'h9CAC,4);
TASK_PP(16'h9CAD,4);
TASK_PP(16'h9CAE,4);
TASK_PP(16'h9CAF,4);
TASK_PP(16'h9CB0,4);
TASK_PP(16'h9CB1,4);
TASK_PP(16'h9CB2,4);
TASK_PP(16'h9CB3,4);
TASK_PP(16'h9CB4,4);
TASK_PP(16'h9CB5,4);
TASK_PP(16'h9CB6,4);
TASK_PP(16'h9CB7,4);
TASK_PP(16'h9CB8,4);
TASK_PP(16'h9CB9,4);
TASK_PP(16'h9CBA,4);
TASK_PP(16'h9CBB,4);
TASK_PP(16'h9CBC,4);
TASK_PP(16'h9CBD,4);
TASK_PP(16'h9CBE,4);
TASK_PP(16'h9CBF,4);
TASK_PP(16'h9CC0,4);
TASK_PP(16'h9CC1,4);
TASK_PP(16'h9CC2,4);
TASK_PP(16'h9CC3,4);
TASK_PP(16'h9CC4,4);
TASK_PP(16'h9CC5,4);
TASK_PP(16'h9CC6,4);
TASK_PP(16'h9CC7,4);
TASK_PP(16'h9CC8,4);
TASK_PP(16'h9CC9,4);
TASK_PP(16'h9CCA,4);
TASK_PP(16'h9CCB,4);
TASK_PP(16'h9CCC,4);
TASK_PP(16'h9CCD,4);
TASK_PP(16'h9CCE,4);
TASK_PP(16'h9CCF,4);
TASK_PP(16'h9CD0,4);
TASK_PP(16'h9CD1,4);
TASK_PP(16'h9CD2,4);
TASK_PP(16'h9CD3,4);
TASK_PP(16'h9CD4,4);
TASK_PP(16'h9CD5,4);
TASK_PP(16'h9CD6,4);
TASK_PP(16'h9CD7,4);
TASK_PP(16'h9CD8,4);
TASK_PP(16'h9CD9,4);
TASK_PP(16'h9CDA,4);
TASK_PP(16'h9CDB,4);
TASK_PP(16'h9CDC,4);
TASK_PP(16'h9CDD,4);
TASK_PP(16'h9CDE,4);
TASK_PP(16'h9CDF,4);
TASK_PP(16'h9CE0,4);
TASK_PP(16'h9CE1,4);
TASK_PP(16'h9CE2,4);
TASK_PP(16'h9CE3,4);
TASK_PP(16'h9CE4,4);
TASK_PP(16'h9CE5,4);
TASK_PP(16'h9CE6,4);
TASK_PP(16'h9CE7,4);
TASK_PP(16'h9CE8,4);
TASK_PP(16'h9CE9,4);
TASK_PP(16'h9CEA,4);
TASK_PP(16'h9CEB,4);
TASK_PP(16'h9CEC,4);
TASK_PP(16'h9CED,4);
TASK_PP(16'h9CEE,4);
TASK_PP(16'h9CEF,4);
TASK_PP(16'h9CF0,4);
TASK_PP(16'h9CF1,4);
TASK_PP(16'h9CF2,4);
TASK_PP(16'h9CF3,4);
TASK_PP(16'h9CF4,4);
TASK_PP(16'h9CF5,4);
TASK_PP(16'h9CF6,4);
TASK_PP(16'h9CF7,4);
TASK_PP(16'h9CF8,4);
TASK_PP(16'h9CF9,4);
TASK_PP(16'h9CFA,4);
TASK_PP(16'h9CFB,4);
TASK_PP(16'h9CFC,4);
TASK_PP(16'h9CFD,4);
TASK_PP(16'h9CFE,4);
TASK_PP(16'h9CFF,4);
TASK_PP(16'h9D00,4);
TASK_PP(16'h9D01,4);
TASK_PP(16'h9D02,4);
TASK_PP(16'h9D03,4);
TASK_PP(16'h9D04,4);
TASK_PP(16'h9D05,4);
TASK_PP(16'h9D06,4);
TASK_PP(16'h9D07,4);
TASK_PP(16'h9D08,4);
TASK_PP(16'h9D09,4);
TASK_PP(16'h9D0A,4);
TASK_PP(16'h9D0B,4);
TASK_PP(16'h9D0C,4);
TASK_PP(16'h9D0D,4);
TASK_PP(16'h9D0E,4);
TASK_PP(16'h9D0F,4);
TASK_PP(16'h9D10,4);
TASK_PP(16'h9D11,4);
TASK_PP(16'h9D12,4);
TASK_PP(16'h9D13,4);
TASK_PP(16'h9D14,4);
TASK_PP(16'h9D15,4);
TASK_PP(16'h9D16,4);
TASK_PP(16'h9D17,4);
TASK_PP(16'h9D18,4);
TASK_PP(16'h9D19,4);
TASK_PP(16'h9D1A,4);
TASK_PP(16'h9D1B,4);
TASK_PP(16'h9D1C,4);
TASK_PP(16'h9D1D,4);
TASK_PP(16'h9D1E,4);
TASK_PP(16'h9D1F,4);
TASK_PP(16'h9D20,4);
TASK_PP(16'h9D21,4);
TASK_PP(16'h9D22,4);
TASK_PP(16'h9D23,4);
TASK_PP(16'h9D24,4);
TASK_PP(16'h9D25,4);
TASK_PP(16'h9D26,4);
TASK_PP(16'h9D27,4);
TASK_PP(16'h9D28,4);
TASK_PP(16'h9D29,4);
TASK_PP(16'h9D2A,4);
TASK_PP(16'h9D2B,4);
TASK_PP(16'h9D2C,4);
TASK_PP(16'h9D2D,4);
TASK_PP(16'h9D2E,4);
TASK_PP(16'h9D2F,4);
TASK_PP(16'h9D30,4);
TASK_PP(16'h9D31,4);
TASK_PP(16'h9D32,4);
TASK_PP(16'h9D33,4);
TASK_PP(16'h9D34,4);
TASK_PP(16'h9D35,4);
TASK_PP(16'h9D36,4);
TASK_PP(16'h9D37,4);
TASK_PP(16'h9D38,4);
TASK_PP(16'h9D39,4);
TASK_PP(16'h9D3A,4);
TASK_PP(16'h9D3B,4);
TASK_PP(16'h9D3C,4);
TASK_PP(16'h9D3D,4);
TASK_PP(16'h9D3E,4);
TASK_PP(16'h9D3F,4);
TASK_PP(16'h9D40,4);
TASK_PP(16'h9D41,4);
TASK_PP(16'h9D42,4);
TASK_PP(16'h9D43,4);
TASK_PP(16'h9D44,4);
TASK_PP(16'h9D45,4);
TASK_PP(16'h9D46,4);
TASK_PP(16'h9D47,4);
TASK_PP(16'h9D48,4);
TASK_PP(16'h9D49,4);
TASK_PP(16'h9D4A,4);
TASK_PP(16'h9D4B,4);
TASK_PP(16'h9D4C,4);
TASK_PP(16'h9D4D,4);
TASK_PP(16'h9D4E,4);
TASK_PP(16'h9D4F,4);
TASK_PP(16'h9D50,4);
TASK_PP(16'h9D51,4);
TASK_PP(16'h9D52,4);
TASK_PP(16'h9D53,4);
TASK_PP(16'h9D54,4);
TASK_PP(16'h9D55,4);
TASK_PP(16'h9D56,4);
TASK_PP(16'h9D57,4);
TASK_PP(16'h9D58,4);
TASK_PP(16'h9D59,4);
TASK_PP(16'h9D5A,4);
TASK_PP(16'h9D5B,4);
TASK_PP(16'h9D5C,4);
TASK_PP(16'h9D5D,4);
TASK_PP(16'h9D5E,4);
TASK_PP(16'h9D5F,4);
TASK_PP(16'h9D60,4);
TASK_PP(16'h9D61,4);
TASK_PP(16'h9D62,4);
TASK_PP(16'h9D63,4);
TASK_PP(16'h9D64,4);
TASK_PP(16'h9D65,4);
TASK_PP(16'h9D66,4);
TASK_PP(16'h9D67,4);
TASK_PP(16'h9D68,4);
TASK_PP(16'h9D69,4);
TASK_PP(16'h9D6A,4);
TASK_PP(16'h9D6B,4);
TASK_PP(16'h9D6C,4);
TASK_PP(16'h9D6D,4);
TASK_PP(16'h9D6E,4);
TASK_PP(16'h9D6F,4);
TASK_PP(16'h9D70,4);
TASK_PP(16'h9D71,4);
TASK_PP(16'h9D72,4);
TASK_PP(16'h9D73,4);
TASK_PP(16'h9D74,4);
TASK_PP(16'h9D75,4);
TASK_PP(16'h9D76,4);
TASK_PP(16'h9D77,4);
TASK_PP(16'h9D78,4);
TASK_PP(16'h9D79,4);
TASK_PP(16'h9D7A,4);
TASK_PP(16'h9D7B,4);
TASK_PP(16'h9D7C,4);
TASK_PP(16'h9D7D,4);
TASK_PP(16'h9D7E,4);
TASK_PP(16'h9D7F,4);
TASK_PP(16'h9D80,4);
TASK_PP(16'h9D81,4);
TASK_PP(16'h9D82,4);
TASK_PP(16'h9D83,4);
TASK_PP(16'h9D84,4);
TASK_PP(16'h9D85,4);
TASK_PP(16'h9D86,4);
TASK_PP(16'h9D87,4);
TASK_PP(16'h9D88,4);
TASK_PP(16'h9D89,4);
TASK_PP(16'h9D8A,4);
TASK_PP(16'h9D8B,4);
TASK_PP(16'h9D8C,4);
TASK_PP(16'h9D8D,4);
TASK_PP(16'h9D8E,4);
TASK_PP(16'h9D8F,4);
TASK_PP(16'h9D90,4);
TASK_PP(16'h9D91,4);
TASK_PP(16'h9D92,4);
TASK_PP(16'h9D93,4);
TASK_PP(16'h9D94,4);
TASK_PP(16'h9D95,4);
TASK_PP(16'h9D96,4);
TASK_PP(16'h9D97,4);
TASK_PP(16'h9D98,4);
TASK_PP(16'h9D99,4);
TASK_PP(16'h9D9A,4);
TASK_PP(16'h9D9B,4);
TASK_PP(16'h9D9C,4);
TASK_PP(16'h9D9D,4);
TASK_PP(16'h9D9E,4);
TASK_PP(16'h9D9F,4);
TASK_PP(16'h9DA0,4);
TASK_PP(16'h9DA1,4);
TASK_PP(16'h9DA2,4);
TASK_PP(16'h9DA3,4);
TASK_PP(16'h9DA4,4);
TASK_PP(16'h9DA5,4);
TASK_PP(16'h9DA6,4);
TASK_PP(16'h9DA7,4);
TASK_PP(16'h9DA8,4);
TASK_PP(16'h9DA9,4);
TASK_PP(16'h9DAA,4);
TASK_PP(16'h9DAB,4);
TASK_PP(16'h9DAC,4);
TASK_PP(16'h9DAD,4);
TASK_PP(16'h9DAE,4);
TASK_PP(16'h9DAF,4);
TASK_PP(16'h9DB0,4);
TASK_PP(16'h9DB1,4);
TASK_PP(16'h9DB2,4);
TASK_PP(16'h9DB3,4);
TASK_PP(16'h9DB4,4);
TASK_PP(16'h9DB5,4);
TASK_PP(16'h9DB6,4);
TASK_PP(16'h9DB7,4);
TASK_PP(16'h9DB8,4);
TASK_PP(16'h9DB9,4);
TASK_PP(16'h9DBA,4);
TASK_PP(16'h9DBB,4);
TASK_PP(16'h9DBC,4);
TASK_PP(16'h9DBD,4);
TASK_PP(16'h9DBE,4);
TASK_PP(16'h9DBF,4);
TASK_PP(16'h9DC0,4);
TASK_PP(16'h9DC1,4);
TASK_PP(16'h9DC2,4);
TASK_PP(16'h9DC3,4);
TASK_PP(16'h9DC4,4);
TASK_PP(16'h9DC5,4);
TASK_PP(16'h9DC6,4);
TASK_PP(16'h9DC7,4);
TASK_PP(16'h9DC8,4);
TASK_PP(16'h9DC9,4);
TASK_PP(16'h9DCA,4);
TASK_PP(16'h9DCB,4);
TASK_PP(16'h9DCC,4);
TASK_PP(16'h9DCD,4);
TASK_PP(16'h9DCE,4);
TASK_PP(16'h9DCF,4);
TASK_PP(16'h9DD0,4);
TASK_PP(16'h9DD1,4);
TASK_PP(16'h9DD2,4);
TASK_PP(16'h9DD3,4);
TASK_PP(16'h9DD4,4);
TASK_PP(16'h9DD5,4);
TASK_PP(16'h9DD6,4);
TASK_PP(16'h9DD7,4);
TASK_PP(16'h9DD8,4);
TASK_PP(16'h9DD9,4);
TASK_PP(16'h9DDA,4);
TASK_PP(16'h9DDB,4);
TASK_PP(16'h9DDC,4);
TASK_PP(16'h9DDD,4);
TASK_PP(16'h9DDE,4);
TASK_PP(16'h9DDF,4);
TASK_PP(16'h9DE0,4);
TASK_PP(16'h9DE1,4);
TASK_PP(16'h9DE2,4);
TASK_PP(16'h9DE3,4);
TASK_PP(16'h9DE4,4);
TASK_PP(16'h9DE5,4);
TASK_PP(16'h9DE6,4);
TASK_PP(16'h9DE7,4);
TASK_PP(16'h9DE8,4);
TASK_PP(16'h9DE9,4);
TASK_PP(16'h9DEA,4);
TASK_PP(16'h9DEB,4);
TASK_PP(16'h9DEC,4);
TASK_PP(16'h9DED,4);
TASK_PP(16'h9DEE,4);
TASK_PP(16'h9DEF,4);
TASK_PP(16'h9DF0,4);
TASK_PP(16'h9DF1,4);
TASK_PP(16'h9DF2,4);
TASK_PP(16'h9DF3,4);
TASK_PP(16'h9DF4,4);
TASK_PP(16'h9DF5,4);
TASK_PP(16'h9DF6,4);
TASK_PP(16'h9DF7,4);
TASK_PP(16'h9DF8,4);
TASK_PP(16'h9DF9,4);
TASK_PP(16'h9DFA,4);
TASK_PP(16'h9DFB,4);
TASK_PP(16'h9DFC,4);
TASK_PP(16'h9DFD,4);
TASK_PP(16'h9DFE,4);
TASK_PP(16'h9DFF,4);
TASK_PP(16'h9E00,4);
TASK_PP(16'h9E01,4);
TASK_PP(16'h9E02,4);
TASK_PP(16'h9E03,4);
TASK_PP(16'h9E04,4);
TASK_PP(16'h9E05,4);
TASK_PP(16'h9E06,4);
TASK_PP(16'h9E07,4);
TASK_PP(16'h9E08,4);
TASK_PP(16'h9E09,4);
TASK_PP(16'h9E0A,4);
TASK_PP(16'h9E0B,4);
TASK_PP(16'h9E0C,4);
TASK_PP(16'h9E0D,4);
TASK_PP(16'h9E0E,4);
TASK_PP(16'h9E0F,4);
TASK_PP(16'h9E10,4);
TASK_PP(16'h9E11,4);
TASK_PP(16'h9E12,4);
TASK_PP(16'h9E13,4);
TASK_PP(16'h9E14,4);
TASK_PP(16'h9E15,4);
TASK_PP(16'h9E16,4);
TASK_PP(16'h9E17,4);
TASK_PP(16'h9E18,4);
TASK_PP(16'h9E19,4);
TASK_PP(16'h9E1A,4);
TASK_PP(16'h9E1B,4);
TASK_PP(16'h9E1C,4);
TASK_PP(16'h9E1D,4);
TASK_PP(16'h9E1E,4);
TASK_PP(16'h9E1F,4);
TASK_PP(16'h9E20,4);
TASK_PP(16'h9E21,4);
TASK_PP(16'h9E22,4);
TASK_PP(16'h9E23,4);
TASK_PP(16'h9E24,4);
TASK_PP(16'h9E25,4);
TASK_PP(16'h9E26,4);
TASK_PP(16'h9E27,4);
TASK_PP(16'h9E28,4);
TASK_PP(16'h9E29,4);
TASK_PP(16'h9E2A,4);
TASK_PP(16'h9E2B,4);
TASK_PP(16'h9E2C,4);
TASK_PP(16'h9E2D,4);
TASK_PP(16'h9E2E,4);
TASK_PP(16'h9E2F,4);
TASK_PP(16'h9E30,4);
TASK_PP(16'h9E31,4);
TASK_PP(16'h9E32,4);
TASK_PP(16'h9E33,4);
TASK_PP(16'h9E34,4);
TASK_PP(16'h9E35,4);
TASK_PP(16'h9E36,4);
TASK_PP(16'h9E37,4);
TASK_PP(16'h9E38,4);
TASK_PP(16'h9E39,4);
TASK_PP(16'h9E3A,4);
TASK_PP(16'h9E3B,4);
TASK_PP(16'h9E3C,4);
TASK_PP(16'h9E3D,4);
TASK_PP(16'h9E3E,4);
TASK_PP(16'h9E3F,4);
TASK_PP(16'h9E40,4);
TASK_PP(16'h9E41,4);
TASK_PP(16'h9E42,4);
TASK_PP(16'h9E43,4);
TASK_PP(16'h9E44,4);
TASK_PP(16'h9E45,4);
TASK_PP(16'h9E46,4);
TASK_PP(16'h9E47,4);
TASK_PP(16'h9E48,4);
TASK_PP(16'h9E49,4);
TASK_PP(16'h9E4A,4);
TASK_PP(16'h9E4B,4);
TASK_PP(16'h9E4C,4);
TASK_PP(16'h9E4D,4);
TASK_PP(16'h9E4E,4);
TASK_PP(16'h9E4F,4);
TASK_PP(16'h9E50,4);
TASK_PP(16'h9E51,4);
TASK_PP(16'h9E52,4);
TASK_PP(16'h9E53,4);
TASK_PP(16'h9E54,4);
TASK_PP(16'h9E55,4);
TASK_PP(16'h9E56,4);
TASK_PP(16'h9E57,4);
TASK_PP(16'h9E58,4);
TASK_PP(16'h9E59,4);
TASK_PP(16'h9E5A,4);
TASK_PP(16'h9E5B,4);
TASK_PP(16'h9E5C,4);
TASK_PP(16'h9E5D,4);
TASK_PP(16'h9E5E,4);
TASK_PP(16'h9E5F,4);
TASK_PP(16'h9E60,4);
TASK_PP(16'h9E61,4);
TASK_PP(16'h9E62,4);
TASK_PP(16'h9E63,4);
TASK_PP(16'h9E64,4);
TASK_PP(16'h9E65,4);
TASK_PP(16'h9E66,4);
TASK_PP(16'h9E67,4);
TASK_PP(16'h9E68,4);
TASK_PP(16'h9E69,4);
TASK_PP(16'h9E6A,4);
TASK_PP(16'h9E6B,4);
TASK_PP(16'h9E6C,4);
TASK_PP(16'h9E6D,4);
TASK_PP(16'h9E6E,4);
TASK_PP(16'h9E6F,4);
TASK_PP(16'h9E70,4);
TASK_PP(16'h9E71,4);
TASK_PP(16'h9E72,4);
TASK_PP(16'h9E73,4);
TASK_PP(16'h9E74,4);
TASK_PP(16'h9E75,4);
TASK_PP(16'h9E76,4);
TASK_PP(16'h9E77,4);
TASK_PP(16'h9E78,4);
TASK_PP(16'h9E79,4);
TASK_PP(16'h9E7A,4);
TASK_PP(16'h9E7B,4);
TASK_PP(16'h9E7C,4);
TASK_PP(16'h9E7D,4);
TASK_PP(16'h9E7E,4);
TASK_PP(16'h9E7F,4);
TASK_PP(16'h9E80,4);
TASK_PP(16'h9E81,4);
TASK_PP(16'h9E82,4);
TASK_PP(16'h9E83,4);
TASK_PP(16'h9E84,4);
TASK_PP(16'h9E85,4);
TASK_PP(16'h9E86,4);
TASK_PP(16'h9E87,4);
TASK_PP(16'h9E88,4);
TASK_PP(16'h9E89,4);
TASK_PP(16'h9E8A,4);
TASK_PP(16'h9E8B,4);
TASK_PP(16'h9E8C,4);
TASK_PP(16'h9E8D,4);
TASK_PP(16'h9E8E,4);
TASK_PP(16'h9E8F,4);
TASK_PP(16'h9E90,4);
TASK_PP(16'h9E91,4);
TASK_PP(16'h9E92,4);
TASK_PP(16'h9E93,4);
TASK_PP(16'h9E94,4);
TASK_PP(16'h9E95,4);
TASK_PP(16'h9E96,4);
TASK_PP(16'h9E97,4);
TASK_PP(16'h9E98,4);
TASK_PP(16'h9E99,4);
TASK_PP(16'h9E9A,4);
TASK_PP(16'h9E9B,4);
TASK_PP(16'h9E9C,4);
TASK_PP(16'h9E9D,4);
TASK_PP(16'h9E9E,4);
TASK_PP(16'h9E9F,4);
TASK_PP(16'h9EA0,4);
TASK_PP(16'h9EA1,4);
TASK_PP(16'h9EA2,4);
TASK_PP(16'h9EA3,4);
TASK_PP(16'h9EA4,4);
TASK_PP(16'h9EA5,4);
TASK_PP(16'h9EA6,4);
TASK_PP(16'h9EA7,4);
TASK_PP(16'h9EA8,4);
TASK_PP(16'h9EA9,4);
TASK_PP(16'h9EAA,4);
TASK_PP(16'h9EAB,4);
TASK_PP(16'h9EAC,4);
TASK_PP(16'h9EAD,4);
TASK_PP(16'h9EAE,4);
TASK_PP(16'h9EAF,4);
TASK_PP(16'h9EB0,4);
TASK_PP(16'h9EB1,4);
TASK_PP(16'h9EB2,4);
TASK_PP(16'h9EB3,4);
TASK_PP(16'h9EB4,4);
TASK_PP(16'h9EB5,4);
TASK_PP(16'h9EB6,4);
TASK_PP(16'h9EB7,4);
TASK_PP(16'h9EB8,4);
TASK_PP(16'h9EB9,4);
TASK_PP(16'h9EBA,4);
TASK_PP(16'h9EBB,4);
TASK_PP(16'h9EBC,4);
TASK_PP(16'h9EBD,4);
TASK_PP(16'h9EBE,4);
TASK_PP(16'h9EBF,4);
TASK_PP(16'h9EC0,4);
TASK_PP(16'h9EC1,4);
TASK_PP(16'h9EC2,4);
TASK_PP(16'h9EC3,4);
TASK_PP(16'h9EC4,4);
TASK_PP(16'h9EC5,4);
TASK_PP(16'h9EC6,4);
TASK_PP(16'h9EC7,4);
TASK_PP(16'h9EC8,4);
TASK_PP(16'h9EC9,4);
TASK_PP(16'h9ECA,4);
TASK_PP(16'h9ECB,4);
TASK_PP(16'h9ECC,4);
TASK_PP(16'h9ECD,4);
TASK_PP(16'h9ECE,4);
TASK_PP(16'h9ECF,4);
TASK_PP(16'h9ED0,4);
TASK_PP(16'h9ED1,4);
TASK_PP(16'h9ED2,4);
TASK_PP(16'h9ED3,4);
TASK_PP(16'h9ED4,4);
TASK_PP(16'h9ED5,4);
TASK_PP(16'h9ED6,4);
TASK_PP(16'h9ED7,4);
TASK_PP(16'h9ED8,4);
TASK_PP(16'h9ED9,4);
TASK_PP(16'h9EDA,4);
TASK_PP(16'h9EDB,4);
TASK_PP(16'h9EDC,4);
TASK_PP(16'h9EDD,4);
TASK_PP(16'h9EDE,4);
TASK_PP(16'h9EDF,4);
TASK_PP(16'h9EE0,4);
TASK_PP(16'h9EE1,4);
TASK_PP(16'h9EE2,4);
TASK_PP(16'h9EE3,4);
TASK_PP(16'h9EE4,4);
TASK_PP(16'h9EE5,4);
TASK_PP(16'h9EE6,4);
TASK_PP(16'h9EE7,4);
TASK_PP(16'h9EE8,4);
TASK_PP(16'h9EE9,4);
TASK_PP(16'h9EEA,4);
TASK_PP(16'h9EEB,4);
TASK_PP(16'h9EEC,4);
TASK_PP(16'h9EED,4);
TASK_PP(16'h9EEE,4);
TASK_PP(16'h9EEF,4);
TASK_PP(16'h9EF0,4);
TASK_PP(16'h9EF1,4);
TASK_PP(16'h9EF2,4);
TASK_PP(16'h9EF3,4);
TASK_PP(16'h9EF4,4);
TASK_PP(16'h9EF5,4);
TASK_PP(16'h9EF6,4);
TASK_PP(16'h9EF7,4);
TASK_PP(16'h9EF8,4);
TASK_PP(16'h9EF9,4);
TASK_PP(16'h9EFA,4);
TASK_PP(16'h9EFB,4);
TASK_PP(16'h9EFC,4);
TASK_PP(16'h9EFD,4);
TASK_PP(16'h9EFE,4);
TASK_PP(16'h9EFF,4);
TASK_PP(16'h9F00,4);
TASK_PP(16'h9F01,4);
TASK_PP(16'h9F02,4);
TASK_PP(16'h9F03,4);
TASK_PP(16'h9F04,4);
TASK_PP(16'h9F05,4);
TASK_PP(16'h9F06,4);
TASK_PP(16'h9F07,4);
TASK_PP(16'h9F08,4);
TASK_PP(16'h9F09,4);
TASK_PP(16'h9F0A,4);
TASK_PP(16'h9F0B,4);
TASK_PP(16'h9F0C,4);
TASK_PP(16'h9F0D,4);
TASK_PP(16'h9F0E,4);
TASK_PP(16'h9F0F,4);
TASK_PP(16'h9F10,4);
TASK_PP(16'h9F11,4);
TASK_PP(16'h9F12,4);
TASK_PP(16'h9F13,4);
TASK_PP(16'h9F14,4);
TASK_PP(16'h9F15,4);
TASK_PP(16'h9F16,4);
TASK_PP(16'h9F17,4);
TASK_PP(16'h9F18,4);
TASK_PP(16'h9F19,4);
TASK_PP(16'h9F1A,4);
TASK_PP(16'h9F1B,4);
TASK_PP(16'h9F1C,4);
TASK_PP(16'h9F1D,4);
TASK_PP(16'h9F1E,4);
TASK_PP(16'h9F1F,4);
TASK_PP(16'h9F20,4);
TASK_PP(16'h9F21,4);
TASK_PP(16'h9F22,4);
TASK_PP(16'h9F23,4);
TASK_PP(16'h9F24,4);
TASK_PP(16'h9F25,4);
TASK_PP(16'h9F26,4);
TASK_PP(16'h9F27,4);
TASK_PP(16'h9F28,4);
TASK_PP(16'h9F29,4);
TASK_PP(16'h9F2A,4);
TASK_PP(16'h9F2B,4);
TASK_PP(16'h9F2C,4);
TASK_PP(16'h9F2D,4);
TASK_PP(16'h9F2E,4);
TASK_PP(16'h9F2F,4);
TASK_PP(16'h9F30,4);
TASK_PP(16'h9F31,4);
TASK_PP(16'h9F32,4);
TASK_PP(16'h9F33,4);
TASK_PP(16'h9F34,4);
TASK_PP(16'h9F35,4);
TASK_PP(16'h9F36,4);
TASK_PP(16'h9F37,4);
TASK_PP(16'h9F38,4);
TASK_PP(16'h9F39,4);
TASK_PP(16'h9F3A,4);
TASK_PP(16'h9F3B,4);
TASK_PP(16'h9F3C,4);
TASK_PP(16'h9F3D,4);
TASK_PP(16'h9F3E,4);
TASK_PP(16'h9F3F,4);
TASK_PP(16'h9F40,4);
TASK_PP(16'h9F41,4);
TASK_PP(16'h9F42,4);
TASK_PP(16'h9F43,4);
TASK_PP(16'h9F44,4);
TASK_PP(16'h9F45,4);
TASK_PP(16'h9F46,4);
TASK_PP(16'h9F47,4);
TASK_PP(16'h9F48,4);
TASK_PP(16'h9F49,4);
TASK_PP(16'h9F4A,4);
TASK_PP(16'h9F4B,4);
TASK_PP(16'h9F4C,4);
TASK_PP(16'h9F4D,4);
TASK_PP(16'h9F4E,4);
TASK_PP(16'h9F4F,4);
TASK_PP(16'h9F50,4);
TASK_PP(16'h9F51,4);
TASK_PP(16'h9F52,4);
TASK_PP(16'h9F53,4);
TASK_PP(16'h9F54,4);
TASK_PP(16'h9F55,4);
TASK_PP(16'h9F56,4);
TASK_PP(16'h9F57,4);
TASK_PP(16'h9F58,4);
TASK_PP(16'h9F59,4);
TASK_PP(16'h9F5A,4);
TASK_PP(16'h9F5B,4);
TASK_PP(16'h9F5C,4);
TASK_PP(16'h9F5D,4);
TASK_PP(16'h9F5E,4);
TASK_PP(16'h9F5F,4);
TASK_PP(16'h9F60,4);
TASK_PP(16'h9F61,4);
TASK_PP(16'h9F62,4);
TASK_PP(16'h9F63,4);
TASK_PP(16'h9F64,4);
TASK_PP(16'h9F65,4);
TASK_PP(16'h9F66,4);
TASK_PP(16'h9F67,4);
TASK_PP(16'h9F68,4);
TASK_PP(16'h9F69,4);
TASK_PP(16'h9F6A,4);
TASK_PP(16'h9F6B,4);
TASK_PP(16'h9F6C,4);
TASK_PP(16'h9F6D,4);
TASK_PP(16'h9F6E,4);
TASK_PP(16'h9F6F,4);
TASK_PP(16'h9F70,4);
TASK_PP(16'h9F71,4);
TASK_PP(16'h9F72,4);
TASK_PP(16'h9F73,4);
TASK_PP(16'h9F74,4);
TASK_PP(16'h9F75,4);
TASK_PP(16'h9F76,4);
TASK_PP(16'h9F77,4);
TASK_PP(16'h9F78,4);
TASK_PP(16'h9F79,4);
TASK_PP(16'h9F7A,4);
TASK_PP(16'h9F7B,4);
TASK_PP(16'h9F7C,4);
TASK_PP(16'h9F7D,4);
TASK_PP(16'h9F7E,4);
TASK_PP(16'h9F7F,4);
TASK_PP(16'h9F80,4);
TASK_PP(16'h9F81,4);
TASK_PP(16'h9F82,4);
TASK_PP(16'h9F83,4);
TASK_PP(16'h9F84,4);
TASK_PP(16'h9F85,4);
TASK_PP(16'h9F86,4);
TASK_PP(16'h9F87,4);
TASK_PP(16'h9F88,4);
TASK_PP(16'h9F89,4);
TASK_PP(16'h9F8A,4);
TASK_PP(16'h9F8B,4);
TASK_PP(16'h9F8C,4);
TASK_PP(16'h9F8D,4);
TASK_PP(16'h9F8E,4);
TASK_PP(16'h9F8F,4);
TASK_PP(16'h9F90,4);
TASK_PP(16'h9F91,4);
TASK_PP(16'h9F92,4);
TASK_PP(16'h9F93,4);
TASK_PP(16'h9F94,4);
TASK_PP(16'h9F95,4);
TASK_PP(16'h9F96,4);
TASK_PP(16'h9F97,4);
TASK_PP(16'h9F98,4);
TASK_PP(16'h9F99,4);
TASK_PP(16'h9F9A,4);
TASK_PP(16'h9F9B,4);
TASK_PP(16'h9F9C,4);
TASK_PP(16'h9F9D,4);
TASK_PP(16'h9F9E,4);
TASK_PP(16'h9F9F,4);
TASK_PP(16'h9FA0,4);
TASK_PP(16'h9FA1,4);
TASK_PP(16'h9FA2,4);
TASK_PP(16'h9FA3,4);
TASK_PP(16'h9FA4,4);
TASK_PP(16'h9FA5,4);
TASK_PP(16'h9FA6,4);
TASK_PP(16'h9FA7,4);
TASK_PP(16'h9FA8,4);
TASK_PP(16'h9FA9,4);
TASK_PP(16'h9FAA,4);
TASK_PP(16'h9FAB,4);
TASK_PP(16'h9FAC,4);
TASK_PP(16'h9FAD,4);
TASK_PP(16'h9FAE,4);
TASK_PP(16'h9FAF,4);
TASK_PP(16'h9FB0,4);
TASK_PP(16'h9FB1,4);
TASK_PP(16'h9FB2,4);
TASK_PP(16'h9FB3,4);
TASK_PP(16'h9FB4,4);
TASK_PP(16'h9FB5,4);
TASK_PP(16'h9FB6,4);
TASK_PP(16'h9FB7,4);
TASK_PP(16'h9FB8,4);
TASK_PP(16'h9FB9,4);
TASK_PP(16'h9FBA,4);
TASK_PP(16'h9FBB,4);
TASK_PP(16'h9FBC,4);
TASK_PP(16'h9FBD,4);
TASK_PP(16'h9FBE,4);
TASK_PP(16'h9FBF,4);
TASK_PP(16'h9FC0,4);
TASK_PP(16'h9FC1,4);
TASK_PP(16'h9FC2,4);
TASK_PP(16'h9FC3,4);
TASK_PP(16'h9FC4,4);
TASK_PP(16'h9FC5,4);
TASK_PP(16'h9FC6,4);
TASK_PP(16'h9FC7,4);
TASK_PP(16'h9FC8,4);
TASK_PP(16'h9FC9,4);
TASK_PP(16'h9FCA,4);
TASK_PP(16'h9FCB,4);
TASK_PP(16'h9FCC,4);
TASK_PP(16'h9FCD,4);
TASK_PP(16'h9FCE,4);
TASK_PP(16'h9FCF,4);
TASK_PP(16'h9FD0,4);
TASK_PP(16'h9FD1,4);
TASK_PP(16'h9FD2,4);
TASK_PP(16'h9FD3,4);
TASK_PP(16'h9FD4,4);
TASK_PP(16'h9FD5,4);
TASK_PP(16'h9FD6,4);
TASK_PP(16'h9FD7,4);
TASK_PP(16'h9FD8,4);
TASK_PP(16'h9FD9,4);
TASK_PP(16'h9FDA,4);
TASK_PP(16'h9FDB,4);
TASK_PP(16'h9FDC,4);
TASK_PP(16'h9FDD,4);
TASK_PP(16'h9FDE,4);
TASK_PP(16'h9FDF,4);
TASK_PP(16'h9FE0,4);
TASK_PP(16'h9FE1,4);
TASK_PP(16'h9FE2,4);
TASK_PP(16'h9FE3,4);
TASK_PP(16'h9FE4,4);
TASK_PP(16'h9FE5,4);
TASK_PP(16'h9FE6,4);
TASK_PP(16'h9FE7,4);
TASK_PP(16'h9FE8,4);
TASK_PP(16'h9FE9,4);
TASK_PP(16'h9FEA,4);
TASK_PP(16'h9FEB,4);
TASK_PP(16'h9FEC,4);
TASK_PP(16'h9FED,4);
TASK_PP(16'h9FEE,4);
TASK_PP(16'h9FEF,4);
TASK_PP(16'h9FF0,4);
TASK_PP(16'h9FF1,4);
TASK_PP(16'h9FF2,4);
TASK_PP(16'h9FF3,4);
TASK_PP(16'h9FF4,4);
TASK_PP(16'h9FF5,4);
TASK_PP(16'h9FF6,4);
TASK_PP(16'h9FF7,4);
TASK_PP(16'h9FF8,4);
TASK_PP(16'h9FF9,4);
TASK_PP(16'h9FFA,4);
TASK_PP(16'h9FFB,4);
TASK_PP(16'h9FFC,4);
TASK_PP(16'h9FFD,4);
TASK_PP(16'h9FFE,4);
TASK_PP(16'h9FFF,4);
TASK_PP(16'hA000,4);
TASK_PP(16'hA001,4);
TASK_PP(16'hA002,4);
TASK_PP(16'hA003,4);
TASK_PP(16'hA004,4);
TASK_PP(16'hA005,4);
TASK_PP(16'hA006,4);
TASK_PP(16'hA007,4);
TASK_PP(16'hA008,4);
TASK_PP(16'hA009,4);
TASK_PP(16'hA00A,4);
TASK_PP(16'hA00B,4);
TASK_PP(16'hA00C,4);
TASK_PP(16'hA00D,4);
TASK_PP(16'hA00E,4);
TASK_PP(16'hA00F,4);
TASK_PP(16'hA010,4);
TASK_PP(16'hA011,4);
TASK_PP(16'hA012,4);
TASK_PP(16'hA013,4);
TASK_PP(16'hA014,4);
TASK_PP(16'hA015,4);
TASK_PP(16'hA016,4);
TASK_PP(16'hA017,4);
TASK_PP(16'hA018,4);
TASK_PP(16'hA019,4);
TASK_PP(16'hA01A,4);
TASK_PP(16'hA01B,4);
TASK_PP(16'hA01C,4);
TASK_PP(16'hA01D,4);
TASK_PP(16'hA01E,4);
TASK_PP(16'hA01F,4);
TASK_PP(16'hA020,4);
TASK_PP(16'hA021,4);
TASK_PP(16'hA022,4);
TASK_PP(16'hA023,4);
TASK_PP(16'hA024,4);
TASK_PP(16'hA025,4);
TASK_PP(16'hA026,4);
TASK_PP(16'hA027,4);
TASK_PP(16'hA028,4);
TASK_PP(16'hA029,4);
TASK_PP(16'hA02A,4);
TASK_PP(16'hA02B,4);
TASK_PP(16'hA02C,4);
TASK_PP(16'hA02D,4);
TASK_PP(16'hA02E,4);
TASK_PP(16'hA02F,4);
TASK_PP(16'hA030,4);
TASK_PP(16'hA031,4);
TASK_PP(16'hA032,4);
TASK_PP(16'hA033,4);
TASK_PP(16'hA034,4);
TASK_PP(16'hA035,4);
TASK_PP(16'hA036,4);
TASK_PP(16'hA037,4);
TASK_PP(16'hA038,4);
TASK_PP(16'hA039,4);
TASK_PP(16'hA03A,4);
TASK_PP(16'hA03B,4);
TASK_PP(16'hA03C,4);
TASK_PP(16'hA03D,4);
TASK_PP(16'hA03E,4);
TASK_PP(16'hA03F,4);
TASK_PP(16'hA040,4);
TASK_PP(16'hA041,4);
TASK_PP(16'hA042,4);
TASK_PP(16'hA043,4);
TASK_PP(16'hA044,4);
TASK_PP(16'hA045,4);
TASK_PP(16'hA046,4);
TASK_PP(16'hA047,4);
TASK_PP(16'hA048,4);
TASK_PP(16'hA049,4);
TASK_PP(16'hA04A,4);
TASK_PP(16'hA04B,4);
TASK_PP(16'hA04C,4);
TASK_PP(16'hA04D,4);
TASK_PP(16'hA04E,4);
TASK_PP(16'hA04F,4);
TASK_PP(16'hA050,4);
TASK_PP(16'hA051,4);
TASK_PP(16'hA052,4);
TASK_PP(16'hA053,4);
TASK_PP(16'hA054,4);
TASK_PP(16'hA055,4);
TASK_PP(16'hA056,4);
TASK_PP(16'hA057,4);
TASK_PP(16'hA058,4);
TASK_PP(16'hA059,4);
TASK_PP(16'hA05A,4);
TASK_PP(16'hA05B,4);
TASK_PP(16'hA05C,4);
TASK_PP(16'hA05D,4);
TASK_PP(16'hA05E,4);
TASK_PP(16'hA05F,4);
TASK_PP(16'hA060,4);
TASK_PP(16'hA061,4);
TASK_PP(16'hA062,4);
TASK_PP(16'hA063,4);
TASK_PP(16'hA064,4);
TASK_PP(16'hA065,4);
TASK_PP(16'hA066,4);
TASK_PP(16'hA067,4);
TASK_PP(16'hA068,4);
TASK_PP(16'hA069,4);
TASK_PP(16'hA06A,4);
TASK_PP(16'hA06B,4);
TASK_PP(16'hA06C,4);
TASK_PP(16'hA06D,4);
TASK_PP(16'hA06E,4);
TASK_PP(16'hA06F,4);
TASK_PP(16'hA070,4);
TASK_PP(16'hA071,4);
TASK_PP(16'hA072,4);
TASK_PP(16'hA073,4);
TASK_PP(16'hA074,4);
TASK_PP(16'hA075,4);
TASK_PP(16'hA076,4);
TASK_PP(16'hA077,4);
TASK_PP(16'hA078,4);
TASK_PP(16'hA079,4);
TASK_PP(16'hA07A,4);
TASK_PP(16'hA07B,4);
TASK_PP(16'hA07C,4);
TASK_PP(16'hA07D,4);
TASK_PP(16'hA07E,4);
TASK_PP(16'hA07F,4);
TASK_PP(16'hA080,4);
TASK_PP(16'hA081,4);
TASK_PP(16'hA082,4);
TASK_PP(16'hA083,4);
TASK_PP(16'hA084,4);
TASK_PP(16'hA085,4);
TASK_PP(16'hA086,4);
TASK_PP(16'hA087,4);
TASK_PP(16'hA088,4);
TASK_PP(16'hA089,4);
TASK_PP(16'hA08A,4);
TASK_PP(16'hA08B,4);
TASK_PP(16'hA08C,4);
TASK_PP(16'hA08D,4);
TASK_PP(16'hA08E,4);
TASK_PP(16'hA08F,4);
TASK_PP(16'hA090,4);
TASK_PP(16'hA091,4);
TASK_PP(16'hA092,4);
TASK_PP(16'hA093,4);
TASK_PP(16'hA094,4);
TASK_PP(16'hA095,4);
TASK_PP(16'hA096,4);
TASK_PP(16'hA097,4);
TASK_PP(16'hA098,4);
TASK_PP(16'hA099,4);
TASK_PP(16'hA09A,4);
TASK_PP(16'hA09B,4);
TASK_PP(16'hA09C,4);
TASK_PP(16'hA09D,4);
TASK_PP(16'hA09E,4);
TASK_PP(16'hA09F,4);
TASK_PP(16'hA0A0,4);
TASK_PP(16'hA0A1,4);
TASK_PP(16'hA0A2,4);
TASK_PP(16'hA0A3,4);
TASK_PP(16'hA0A4,4);
TASK_PP(16'hA0A5,4);
TASK_PP(16'hA0A6,4);
TASK_PP(16'hA0A7,4);
TASK_PP(16'hA0A8,4);
TASK_PP(16'hA0A9,4);
TASK_PP(16'hA0AA,4);
TASK_PP(16'hA0AB,4);
TASK_PP(16'hA0AC,4);
TASK_PP(16'hA0AD,4);
TASK_PP(16'hA0AE,4);
TASK_PP(16'hA0AF,4);
TASK_PP(16'hA0B0,4);
TASK_PP(16'hA0B1,4);
TASK_PP(16'hA0B2,4);
TASK_PP(16'hA0B3,4);
TASK_PP(16'hA0B4,4);
TASK_PP(16'hA0B5,4);
TASK_PP(16'hA0B6,4);
TASK_PP(16'hA0B7,4);
TASK_PP(16'hA0B8,4);
TASK_PP(16'hA0B9,4);
TASK_PP(16'hA0BA,4);
TASK_PP(16'hA0BB,4);
TASK_PP(16'hA0BC,4);
TASK_PP(16'hA0BD,4);
TASK_PP(16'hA0BE,4);
TASK_PP(16'hA0BF,4);
TASK_PP(16'hA0C0,4);
TASK_PP(16'hA0C1,4);
TASK_PP(16'hA0C2,4);
TASK_PP(16'hA0C3,4);
TASK_PP(16'hA0C4,4);
TASK_PP(16'hA0C5,4);
TASK_PP(16'hA0C6,4);
TASK_PP(16'hA0C7,4);
TASK_PP(16'hA0C8,4);
TASK_PP(16'hA0C9,4);
TASK_PP(16'hA0CA,4);
TASK_PP(16'hA0CB,4);
TASK_PP(16'hA0CC,4);
TASK_PP(16'hA0CD,4);
TASK_PP(16'hA0CE,4);
TASK_PP(16'hA0CF,4);
TASK_PP(16'hA0D0,4);
TASK_PP(16'hA0D1,4);
TASK_PP(16'hA0D2,4);
TASK_PP(16'hA0D3,4);
TASK_PP(16'hA0D4,4);
TASK_PP(16'hA0D5,4);
TASK_PP(16'hA0D6,4);
TASK_PP(16'hA0D7,4);
TASK_PP(16'hA0D8,4);
TASK_PP(16'hA0D9,4);
TASK_PP(16'hA0DA,4);
TASK_PP(16'hA0DB,4);
TASK_PP(16'hA0DC,4);
TASK_PP(16'hA0DD,4);
TASK_PP(16'hA0DE,4);
TASK_PP(16'hA0DF,4);
TASK_PP(16'hA0E0,4);
TASK_PP(16'hA0E1,4);
TASK_PP(16'hA0E2,4);
TASK_PP(16'hA0E3,4);
TASK_PP(16'hA0E4,4);
TASK_PP(16'hA0E5,4);
TASK_PP(16'hA0E6,4);
TASK_PP(16'hA0E7,4);
TASK_PP(16'hA0E8,4);
TASK_PP(16'hA0E9,4);
TASK_PP(16'hA0EA,4);
TASK_PP(16'hA0EB,4);
TASK_PP(16'hA0EC,4);
TASK_PP(16'hA0ED,4);
TASK_PP(16'hA0EE,4);
TASK_PP(16'hA0EF,4);
TASK_PP(16'hA0F0,4);
TASK_PP(16'hA0F1,4);
TASK_PP(16'hA0F2,4);
TASK_PP(16'hA0F3,4);
TASK_PP(16'hA0F4,4);
TASK_PP(16'hA0F5,4);
TASK_PP(16'hA0F6,4);
TASK_PP(16'hA0F7,4);
TASK_PP(16'hA0F8,4);
TASK_PP(16'hA0F9,4);
TASK_PP(16'hA0FA,4);
TASK_PP(16'hA0FB,4);
TASK_PP(16'hA0FC,4);
TASK_PP(16'hA0FD,4);
TASK_PP(16'hA0FE,4);
TASK_PP(16'hA0FF,4);
TASK_PP(16'hA100,4);
TASK_PP(16'hA101,4);
TASK_PP(16'hA102,4);
TASK_PP(16'hA103,4);
TASK_PP(16'hA104,4);
TASK_PP(16'hA105,4);
TASK_PP(16'hA106,4);
TASK_PP(16'hA107,4);
TASK_PP(16'hA108,4);
TASK_PP(16'hA109,4);
TASK_PP(16'hA10A,4);
TASK_PP(16'hA10B,4);
TASK_PP(16'hA10C,4);
TASK_PP(16'hA10D,4);
TASK_PP(16'hA10E,4);
TASK_PP(16'hA10F,4);
TASK_PP(16'hA110,4);
TASK_PP(16'hA111,4);
TASK_PP(16'hA112,4);
TASK_PP(16'hA113,4);
TASK_PP(16'hA114,4);
TASK_PP(16'hA115,4);
TASK_PP(16'hA116,4);
TASK_PP(16'hA117,4);
TASK_PP(16'hA118,4);
TASK_PP(16'hA119,4);
TASK_PP(16'hA11A,4);
TASK_PP(16'hA11B,4);
TASK_PP(16'hA11C,4);
TASK_PP(16'hA11D,4);
TASK_PP(16'hA11E,4);
TASK_PP(16'hA11F,4);
TASK_PP(16'hA120,4);
TASK_PP(16'hA121,4);
TASK_PP(16'hA122,4);
TASK_PP(16'hA123,4);
TASK_PP(16'hA124,4);
TASK_PP(16'hA125,4);
TASK_PP(16'hA126,4);
TASK_PP(16'hA127,4);
TASK_PP(16'hA128,4);
TASK_PP(16'hA129,4);
TASK_PP(16'hA12A,4);
TASK_PP(16'hA12B,4);
TASK_PP(16'hA12C,4);
TASK_PP(16'hA12D,4);
TASK_PP(16'hA12E,4);
TASK_PP(16'hA12F,4);
TASK_PP(16'hA130,4);
TASK_PP(16'hA131,4);
TASK_PP(16'hA132,4);
TASK_PP(16'hA133,4);
TASK_PP(16'hA134,4);
TASK_PP(16'hA135,4);
TASK_PP(16'hA136,4);
TASK_PP(16'hA137,4);
TASK_PP(16'hA138,4);
TASK_PP(16'hA139,4);
TASK_PP(16'hA13A,4);
TASK_PP(16'hA13B,4);
TASK_PP(16'hA13C,4);
TASK_PP(16'hA13D,4);
TASK_PP(16'hA13E,4);
TASK_PP(16'hA13F,4);
TASK_PP(16'hA140,4);
TASK_PP(16'hA141,4);
TASK_PP(16'hA142,4);
TASK_PP(16'hA143,4);
TASK_PP(16'hA144,4);
TASK_PP(16'hA145,4);
TASK_PP(16'hA146,4);
TASK_PP(16'hA147,4);
TASK_PP(16'hA148,4);
TASK_PP(16'hA149,4);
TASK_PP(16'hA14A,4);
TASK_PP(16'hA14B,4);
TASK_PP(16'hA14C,4);
TASK_PP(16'hA14D,4);
TASK_PP(16'hA14E,4);
TASK_PP(16'hA14F,4);
TASK_PP(16'hA150,4);
TASK_PP(16'hA151,4);
TASK_PP(16'hA152,4);
TASK_PP(16'hA153,4);
TASK_PP(16'hA154,4);
TASK_PP(16'hA155,4);
TASK_PP(16'hA156,4);
TASK_PP(16'hA157,4);
TASK_PP(16'hA158,4);
TASK_PP(16'hA159,4);
TASK_PP(16'hA15A,4);
TASK_PP(16'hA15B,4);
TASK_PP(16'hA15C,4);
TASK_PP(16'hA15D,4);
TASK_PP(16'hA15E,4);
TASK_PP(16'hA15F,4);
TASK_PP(16'hA160,4);
TASK_PP(16'hA161,4);
TASK_PP(16'hA162,4);
TASK_PP(16'hA163,4);
TASK_PP(16'hA164,4);
TASK_PP(16'hA165,4);
TASK_PP(16'hA166,4);
TASK_PP(16'hA167,4);
TASK_PP(16'hA168,4);
TASK_PP(16'hA169,4);
TASK_PP(16'hA16A,4);
TASK_PP(16'hA16B,4);
TASK_PP(16'hA16C,4);
TASK_PP(16'hA16D,4);
TASK_PP(16'hA16E,4);
TASK_PP(16'hA16F,4);
TASK_PP(16'hA170,4);
TASK_PP(16'hA171,4);
TASK_PP(16'hA172,4);
TASK_PP(16'hA173,4);
TASK_PP(16'hA174,4);
TASK_PP(16'hA175,4);
TASK_PP(16'hA176,4);
TASK_PP(16'hA177,4);
TASK_PP(16'hA178,4);
TASK_PP(16'hA179,4);
TASK_PP(16'hA17A,4);
TASK_PP(16'hA17B,4);
TASK_PP(16'hA17C,4);
TASK_PP(16'hA17D,4);
TASK_PP(16'hA17E,4);
TASK_PP(16'hA17F,4);
TASK_PP(16'hA180,4);
TASK_PP(16'hA181,4);
TASK_PP(16'hA182,4);
TASK_PP(16'hA183,4);
TASK_PP(16'hA184,4);
TASK_PP(16'hA185,4);
TASK_PP(16'hA186,4);
TASK_PP(16'hA187,4);
TASK_PP(16'hA188,4);
TASK_PP(16'hA189,4);
TASK_PP(16'hA18A,4);
TASK_PP(16'hA18B,4);
TASK_PP(16'hA18C,4);
TASK_PP(16'hA18D,4);
TASK_PP(16'hA18E,4);
TASK_PP(16'hA18F,4);
TASK_PP(16'hA190,4);
TASK_PP(16'hA191,4);
TASK_PP(16'hA192,4);
TASK_PP(16'hA193,4);
TASK_PP(16'hA194,4);
TASK_PP(16'hA195,4);
TASK_PP(16'hA196,4);
TASK_PP(16'hA197,4);
TASK_PP(16'hA198,4);
TASK_PP(16'hA199,4);
TASK_PP(16'hA19A,4);
TASK_PP(16'hA19B,4);
TASK_PP(16'hA19C,4);
TASK_PP(16'hA19D,4);
TASK_PP(16'hA19E,4);
TASK_PP(16'hA19F,4);
TASK_PP(16'hA1A0,4);
TASK_PP(16'hA1A1,4);
TASK_PP(16'hA1A2,4);
TASK_PP(16'hA1A3,4);
TASK_PP(16'hA1A4,4);
TASK_PP(16'hA1A5,4);
TASK_PP(16'hA1A6,4);
TASK_PP(16'hA1A7,4);
TASK_PP(16'hA1A8,4);
TASK_PP(16'hA1A9,4);
TASK_PP(16'hA1AA,4);
TASK_PP(16'hA1AB,4);
TASK_PP(16'hA1AC,4);
TASK_PP(16'hA1AD,4);
TASK_PP(16'hA1AE,4);
TASK_PP(16'hA1AF,4);
TASK_PP(16'hA1B0,4);
TASK_PP(16'hA1B1,4);
TASK_PP(16'hA1B2,4);
TASK_PP(16'hA1B3,4);
TASK_PP(16'hA1B4,4);
TASK_PP(16'hA1B5,4);
TASK_PP(16'hA1B6,4);
TASK_PP(16'hA1B7,4);
TASK_PP(16'hA1B8,4);
TASK_PP(16'hA1B9,4);
TASK_PP(16'hA1BA,4);
TASK_PP(16'hA1BB,4);
TASK_PP(16'hA1BC,4);
TASK_PP(16'hA1BD,4);
TASK_PP(16'hA1BE,4);
TASK_PP(16'hA1BF,4);
TASK_PP(16'hA1C0,4);
TASK_PP(16'hA1C1,4);
TASK_PP(16'hA1C2,4);
TASK_PP(16'hA1C3,4);
TASK_PP(16'hA1C4,4);
TASK_PP(16'hA1C5,4);
TASK_PP(16'hA1C6,4);
TASK_PP(16'hA1C7,4);
TASK_PP(16'hA1C8,4);
TASK_PP(16'hA1C9,4);
TASK_PP(16'hA1CA,4);
TASK_PP(16'hA1CB,4);
TASK_PP(16'hA1CC,4);
TASK_PP(16'hA1CD,4);
TASK_PP(16'hA1CE,4);
TASK_PP(16'hA1CF,4);
TASK_PP(16'hA1D0,4);
TASK_PP(16'hA1D1,4);
TASK_PP(16'hA1D2,4);
TASK_PP(16'hA1D3,4);
TASK_PP(16'hA1D4,4);
TASK_PP(16'hA1D5,4);
TASK_PP(16'hA1D6,4);
TASK_PP(16'hA1D7,4);
TASK_PP(16'hA1D8,4);
TASK_PP(16'hA1D9,4);
TASK_PP(16'hA1DA,4);
TASK_PP(16'hA1DB,4);
TASK_PP(16'hA1DC,4);
TASK_PP(16'hA1DD,4);
TASK_PP(16'hA1DE,4);
TASK_PP(16'hA1DF,4);
TASK_PP(16'hA1E0,4);
TASK_PP(16'hA1E1,4);
TASK_PP(16'hA1E2,4);
TASK_PP(16'hA1E3,4);
TASK_PP(16'hA1E4,4);
TASK_PP(16'hA1E5,4);
TASK_PP(16'hA1E6,4);
TASK_PP(16'hA1E7,4);
TASK_PP(16'hA1E8,4);
TASK_PP(16'hA1E9,4);
TASK_PP(16'hA1EA,4);
TASK_PP(16'hA1EB,4);
TASK_PP(16'hA1EC,4);
TASK_PP(16'hA1ED,4);
TASK_PP(16'hA1EE,4);
TASK_PP(16'hA1EF,4);
TASK_PP(16'hA1F0,4);
TASK_PP(16'hA1F1,4);
TASK_PP(16'hA1F2,4);
TASK_PP(16'hA1F3,4);
TASK_PP(16'hA1F4,4);
TASK_PP(16'hA1F5,4);
TASK_PP(16'hA1F6,4);
TASK_PP(16'hA1F7,4);
TASK_PP(16'hA1F8,4);
TASK_PP(16'hA1F9,4);
TASK_PP(16'hA1FA,4);
TASK_PP(16'hA1FB,4);
TASK_PP(16'hA1FC,4);
TASK_PP(16'hA1FD,4);
TASK_PP(16'hA1FE,4);
TASK_PP(16'hA1FF,4);
TASK_PP(16'hA200,4);
TASK_PP(16'hA201,4);
TASK_PP(16'hA202,4);
TASK_PP(16'hA203,4);
TASK_PP(16'hA204,4);
TASK_PP(16'hA205,4);
TASK_PP(16'hA206,4);
TASK_PP(16'hA207,4);
TASK_PP(16'hA208,4);
TASK_PP(16'hA209,4);
TASK_PP(16'hA20A,4);
TASK_PP(16'hA20B,4);
TASK_PP(16'hA20C,4);
TASK_PP(16'hA20D,4);
TASK_PP(16'hA20E,4);
TASK_PP(16'hA20F,4);
TASK_PP(16'hA210,4);
TASK_PP(16'hA211,4);
TASK_PP(16'hA212,4);
TASK_PP(16'hA213,4);
TASK_PP(16'hA214,4);
TASK_PP(16'hA215,4);
TASK_PP(16'hA216,4);
TASK_PP(16'hA217,4);
TASK_PP(16'hA218,4);
TASK_PP(16'hA219,4);
TASK_PP(16'hA21A,4);
TASK_PP(16'hA21B,4);
TASK_PP(16'hA21C,4);
TASK_PP(16'hA21D,4);
TASK_PP(16'hA21E,4);
TASK_PP(16'hA21F,4);
TASK_PP(16'hA220,4);
TASK_PP(16'hA221,4);
TASK_PP(16'hA222,4);
TASK_PP(16'hA223,4);
TASK_PP(16'hA224,4);
TASK_PP(16'hA225,4);
TASK_PP(16'hA226,4);
TASK_PP(16'hA227,4);
TASK_PP(16'hA228,4);
TASK_PP(16'hA229,4);
TASK_PP(16'hA22A,4);
TASK_PP(16'hA22B,4);
TASK_PP(16'hA22C,4);
TASK_PP(16'hA22D,4);
TASK_PP(16'hA22E,4);
TASK_PP(16'hA22F,4);
TASK_PP(16'hA230,4);
TASK_PP(16'hA231,4);
TASK_PP(16'hA232,4);
TASK_PP(16'hA233,4);
TASK_PP(16'hA234,4);
TASK_PP(16'hA235,4);
TASK_PP(16'hA236,4);
TASK_PP(16'hA237,4);
TASK_PP(16'hA238,4);
TASK_PP(16'hA239,4);
TASK_PP(16'hA23A,4);
TASK_PP(16'hA23B,4);
TASK_PP(16'hA23C,4);
TASK_PP(16'hA23D,4);
TASK_PP(16'hA23E,4);
TASK_PP(16'hA23F,4);
TASK_PP(16'hA240,4);
TASK_PP(16'hA241,4);
TASK_PP(16'hA242,4);
TASK_PP(16'hA243,4);
TASK_PP(16'hA244,4);
TASK_PP(16'hA245,4);
TASK_PP(16'hA246,4);
TASK_PP(16'hA247,4);
TASK_PP(16'hA248,4);
TASK_PP(16'hA249,4);
TASK_PP(16'hA24A,4);
TASK_PP(16'hA24B,4);
TASK_PP(16'hA24C,4);
TASK_PP(16'hA24D,4);
TASK_PP(16'hA24E,4);
TASK_PP(16'hA24F,4);
TASK_PP(16'hA250,4);
TASK_PP(16'hA251,4);
TASK_PP(16'hA252,4);
TASK_PP(16'hA253,4);
TASK_PP(16'hA254,4);
TASK_PP(16'hA255,4);
TASK_PP(16'hA256,4);
TASK_PP(16'hA257,4);
TASK_PP(16'hA258,4);
TASK_PP(16'hA259,4);
TASK_PP(16'hA25A,4);
TASK_PP(16'hA25B,4);
TASK_PP(16'hA25C,4);
TASK_PP(16'hA25D,4);
TASK_PP(16'hA25E,4);
TASK_PP(16'hA25F,4);
TASK_PP(16'hA260,4);
TASK_PP(16'hA261,4);
TASK_PP(16'hA262,4);
TASK_PP(16'hA263,4);
TASK_PP(16'hA264,4);
TASK_PP(16'hA265,4);
TASK_PP(16'hA266,4);
TASK_PP(16'hA267,4);
TASK_PP(16'hA268,4);
TASK_PP(16'hA269,4);
TASK_PP(16'hA26A,4);
TASK_PP(16'hA26B,4);
TASK_PP(16'hA26C,4);
TASK_PP(16'hA26D,4);
TASK_PP(16'hA26E,4);
TASK_PP(16'hA26F,4);
TASK_PP(16'hA270,4);
TASK_PP(16'hA271,4);
TASK_PP(16'hA272,4);
TASK_PP(16'hA273,4);
TASK_PP(16'hA274,4);
TASK_PP(16'hA275,4);
TASK_PP(16'hA276,4);
TASK_PP(16'hA277,4);
TASK_PP(16'hA278,4);
TASK_PP(16'hA279,4);
TASK_PP(16'hA27A,4);
TASK_PP(16'hA27B,4);
TASK_PP(16'hA27C,4);
TASK_PP(16'hA27D,4);
TASK_PP(16'hA27E,4);
TASK_PP(16'hA27F,4);
TASK_PP(16'hA280,4);
TASK_PP(16'hA281,4);
TASK_PP(16'hA282,4);
TASK_PP(16'hA283,4);
TASK_PP(16'hA284,4);
TASK_PP(16'hA285,4);
TASK_PP(16'hA286,4);
TASK_PP(16'hA287,4);
TASK_PP(16'hA288,4);
TASK_PP(16'hA289,4);
TASK_PP(16'hA28A,4);
TASK_PP(16'hA28B,4);
TASK_PP(16'hA28C,4);
TASK_PP(16'hA28D,4);
TASK_PP(16'hA28E,4);
TASK_PP(16'hA28F,4);
TASK_PP(16'hA290,4);
TASK_PP(16'hA291,4);
TASK_PP(16'hA292,4);
TASK_PP(16'hA293,4);
TASK_PP(16'hA294,4);
TASK_PP(16'hA295,4);
TASK_PP(16'hA296,4);
TASK_PP(16'hA297,4);
TASK_PP(16'hA298,4);
TASK_PP(16'hA299,4);
TASK_PP(16'hA29A,4);
TASK_PP(16'hA29B,4);
TASK_PP(16'hA29C,4);
TASK_PP(16'hA29D,4);
TASK_PP(16'hA29E,4);
TASK_PP(16'hA29F,4);
TASK_PP(16'hA2A0,4);
TASK_PP(16'hA2A1,4);
TASK_PP(16'hA2A2,4);
TASK_PP(16'hA2A3,4);
TASK_PP(16'hA2A4,4);
TASK_PP(16'hA2A5,4);
TASK_PP(16'hA2A6,4);
TASK_PP(16'hA2A7,4);
TASK_PP(16'hA2A8,4);
TASK_PP(16'hA2A9,4);
TASK_PP(16'hA2AA,4);
TASK_PP(16'hA2AB,4);
TASK_PP(16'hA2AC,4);
TASK_PP(16'hA2AD,4);
TASK_PP(16'hA2AE,4);
TASK_PP(16'hA2AF,4);
TASK_PP(16'hA2B0,4);
TASK_PP(16'hA2B1,4);
TASK_PP(16'hA2B2,4);
TASK_PP(16'hA2B3,4);
TASK_PP(16'hA2B4,4);
TASK_PP(16'hA2B5,4);
TASK_PP(16'hA2B6,4);
TASK_PP(16'hA2B7,4);
TASK_PP(16'hA2B8,4);
TASK_PP(16'hA2B9,4);
TASK_PP(16'hA2BA,4);
TASK_PP(16'hA2BB,4);
TASK_PP(16'hA2BC,4);
TASK_PP(16'hA2BD,4);
TASK_PP(16'hA2BE,4);
TASK_PP(16'hA2BF,4);
TASK_PP(16'hA2C0,4);
TASK_PP(16'hA2C1,4);
TASK_PP(16'hA2C2,4);
TASK_PP(16'hA2C3,4);
TASK_PP(16'hA2C4,4);
TASK_PP(16'hA2C5,4);
TASK_PP(16'hA2C6,4);
TASK_PP(16'hA2C7,4);
TASK_PP(16'hA2C8,4);
TASK_PP(16'hA2C9,4);
TASK_PP(16'hA2CA,4);
TASK_PP(16'hA2CB,4);
TASK_PP(16'hA2CC,4);
TASK_PP(16'hA2CD,4);
TASK_PP(16'hA2CE,4);
TASK_PP(16'hA2CF,4);
TASK_PP(16'hA2D0,4);
TASK_PP(16'hA2D1,4);
TASK_PP(16'hA2D2,4);
TASK_PP(16'hA2D3,4);
TASK_PP(16'hA2D4,4);
TASK_PP(16'hA2D5,4);
TASK_PP(16'hA2D6,4);
TASK_PP(16'hA2D7,4);
TASK_PP(16'hA2D8,4);
TASK_PP(16'hA2D9,4);
TASK_PP(16'hA2DA,4);
TASK_PP(16'hA2DB,4);
TASK_PP(16'hA2DC,4);
TASK_PP(16'hA2DD,4);
TASK_PP(16'hA2DE,4);
TASK_PP(16'hA2DF,4);
TASK_PP(16'hA2E0,4);
TASK_PP(16'hA2E1,4);
TASK_PP(16'hA2E2,4);
TASK_PP(16'hA2E3,4);
TASK_PP(16'hA2E4,4);
TASK_PP(16'hA2E5,4);
TASK_PP(16'hA2E6,4);
TASK_PP(16'hA2E7,4);
TASK_PP(16'hA2E8,4);
TASK_PP(16'hA2E9,4);
TASK_PP(16'hA2EA,4);
TASK_PP(16'hA2EB,4);
TASK_PP(16'hA2EC,4);
TASK_PP(16'hA2ED,4);
TASK_PP(16'hA2EE,4);
TASK_PP(16'hA2EF,4);
TASK_PP(16'hA2F0,4);
TASK_PP(16'hA2F1,4);
TASK_PP(16'hA2F2,4);
TASK_PP(16'hA2F3,4);
TASK_PP(16'hA2F4,4);
TASK_PP(16'hA2F5,4);
TASK_PP(16'hA2F6,4);
TASK_PP(16'hA2F7,4);
TASK_PP(16'hA2F8,4);
TASK_PP(16'hA2F9,4);
TASK_PP(16'hA2FA,4);
TASK_PP(16'hA2FB,4);
TASK_PP(16'hA2FC,4);
TASK_PP(16'hA2FD,4);
TASK_PP(16'hA2FE,4);
TASK_PP(16'hA2FF,4);
TASK_PP(16'hA300,4);
TASK_PP(16'hA301,4);
TASK_PP(16'hA302,4);
TASK_PP(16'hA303,4);
TASK_PP(16'hA304,4);
TASK_PP(16'hA305,4);
TASK_PP(16'hA306,4);
TASK_PP(16'hA307,4);
TASK_PP(16'hA308,4);
TASK_PP(16'hA309,4);
TASK_PP(16'hA30A,4);
TASK_PP(16'hA30B,4);
TASK_PP(16'hA30C,4);
TASK_PP(16'hA30D,4);
TASK_PP(16'hA30E,4);
TASK_PP(16'hA30F,4);
TASK_PP(16'hA310,4);
TASK_PP(16'hA311,4);
TASK_PP(16'hA312,4);
TASK_PP(16'hA313,4);
TASK_PP(16'hA314,4);
TASK_PP(16'hA315,4);
TASK_PP(16'hA316,4);
TASK_PP(16'hA317,4);
TASK_PP(16'hA318,4);
TASK_PP(16'hA319,4);
TASK_PP(16'hA31A,4);
TASK_PP(16'hA31B,4);
TASK_PP(16'hA31C,4);
TASK_PP(16'hA31D,4);
TASK_PP(16'hA31E,4);
TASK_PP(16'hA31F,4);
TASK_PP(16'hA320,4);
TASK_PP(16'hA321,4);
TASK_PP(16'hA322,4);
TASK_PP(16'hA323,4);
TASK_PP(16'hA324,4);
TASK_PP(16'hA325,4);
TASK_PP(16'hA326,4);
TASK_PP(16'hA327,4);
TASK_PP(16'hA328,4);
TASK_PP(16'hA329,4);
TASK_PP(16'hA32A,4);
TASK_PP(16'hA32B,4);
TASK_PP(16'hA32C,4);
TASK_PP(16'hA32D,4);
TASK_PP(16'hA32E,4);
TASK_PP(16'hA32F,4);
TASK_PP(16'hA330,4);
TASK_PP(16'hA331,4);
TASK_PP(16'hA332,4);
TASK_PP(16'hA333,4);
TASK_PP(16'hA334,4);
TASK_PP(16'hA335,4);
TASK_PP(16'hA336,4);
TASK_PP(16'hA337,4);
TASK_PP(16'hA338,4);
TASK_PP(16'hA339,4);
TASK_PP(16'hA33A,4);
TASK_PP(16'hA33B,4);
TASK_PP(16'hA33C,4);
TASK_PP(16'hA33D,4);
TASK_PP(16'hA33E,4);
TASK_PP(16'hA33F,4);
TASK_PP(16'hA340,4);
TASK_PP(16'hA341,4);
TASK_PP(16'hA342,4);
TASK_PP(16'hA343,4);
TASK_PP(16'hA344,4);
TASK_PP(16'hA345,4);
TASK_PP(16'hA346,4);
TASK_PP(16'hA347,4);
TASK_PP(16'hA348,4);
TASK_PP(16'hA349,4);
TASK_PP(16'hA34A,4);
TASK_PP(16'hA34B,4);
TASK_PP(16'hA34C,4);
TASK_PP(16'hA34D,4);
TASK_PP(16'hA34E,4);
TASK_PP(16'hA34F,4);
TASK_PP(16'hA350,4);
TASK_PP(16'hA351,4);
TASK_PP(16'hA352,4);
TASK_PP(16'hA353,4);
TASK_PP(16'hA354,4);
TASK_PP(16'hA355,4);
TASK_PP(16'hA356,4);
TASK_PP(16'hA357,4);
TASK_PP(16'hA358,4);
TASK_PP(16'hA359,4);
TASK_PP(16'hA35A,4);
TASK_PP(16'hA35B,4);
TASK_PP(16'hA35C,4);
TASK_PP(16'hA35D,4);
TASK_PP(16'hA35E,4);
TASK_PP(16'hA35F,4);
TASK_PP(16'hA360,4);
TASK_PP(16'hA361,4);
TASK_PP(16'hA362,4);
TASK_PP(16'hA363,4);
TASK_PP(16'hA364,4);
TASK_PP(16'hA365,4);
TASK_PP(16'hA366,4);
TASK_PP(16'hA367,4);
TASK_PP(16'hA368,4);
TASK_PP(16'hA369,4);
TASK_PP(16'hA36A,4);
TASK_PP(16'hA36B,4);
TASK_PP(16'hA36C,4);
TASK_PP(16'hA36D,4);
TASK_PP(16'hA36E,4);
TASK_PP(16'hA36F,4);
TASK_PP(16'hA370,4);
TASK_PP(16'hA371,4);
TASK_PP(16'hA372,4);
TASK_PP(16'hA373,4);
TASK_PP(16'hA374,4);
TASK_PP(16'hA375,4);
TASK_PP(16'hA376,4);
TASK_PP(16'hA377,4);
TASK_PP(16'hA378,4);
TASK_PP(16'hA379,4);
TASK_PP(16'hA37A,4);
TASK_PP(16'hA37B,4);
TASK_PP(16'hA37C,4);
TASK_PP(16'hA37D,4);
TASK_PP(16'hA37E,4);
TASK_PP(16'hA37F,4);
TASK_PP(16'hA380,4);
TASK_PP(16'hA381,4);
TASK_PP(16'hA382,4);
TASK_PP(16'hA383,4);
TASK_PP(16'hA384,4);
TASK_PP(16'hA385,4);
TASK_PP(16'hA386,4);
TASK_PP(16'hA387,4);
TASK_PP(16'hA388,4);
TASK_PP(16'hA389,4);
TASK_PP(16'hA38A,4);
TASK_PP(16'hA38B,4);
TASK_PP(16'hA38C,4);
TASK_PP(16'hA38D,4);
TASK_PP(16'hA38E,4);
TASK_PP(16'hA38F,4);
TASK_PP(16'hA390,4);
TASK_PP(16'hA391,4);
TASK_PP(16'hA392,4);
TASK_PP(16'hA393,4);
TASK_PP(16'hA394,4);
TASK_PP(16'hA395,4);
TASK_PP(16'hA396,4);
TASK_PP(16'hA397,4);
TASK_PP(16'hA398,4);
TASK_PP(16'hA399,4);
TASK_PP(16'hA39A,4);
TASK_PP(16'hA39B,4);
TASK_PP(16'hA39C,4);
TASK_PP(16'hA39D,4);
TASK_PP(16'hA39E,4);
TASK_PP(16'hA39F,4);
TASK_PP(16'hA3A0,4);
TASK_PP(16'hA3A1,4);
TASK_PP(16'hA3A2,4);
TASK_PP(16'hA3A3,4);
TASK_PP(16'hA3A4,4);
TASK_PP(16'hA3A5,4);
TASK_PP(16'hA3A6,4);
TASK_PP(16'hA3A7,4);
TASK_PP(16'hA3A8,4);
TASK_PP(16'hA3A9,4);
TASK_PP(16'hA3AA,4);
TASK_PP(16'hA3AB,4);
TASK_PP(16'hA3AC,4);
TASK_PP(16'hA3AD,4);
TASK_PP(16'hA3AE,4);
TASK_PP(16'hA3AF,4);
TASK_PP(16'hA3B0,4);
TASK_PP(16'hA3B1,4);
TASK_PP(16'hA3B2,4);
TASK_PP(16'hA3B3,4);
TASK_PP(16'hA3B4,4);
TASK_PP(16'hA3B5,4);
TASK_PP(16'hA3B6,4);
TASK_PP(16'hA3B7,4);
TASK_PP(16'hA3B8,4);
TASK_PP(16'hA3B9,4);
TASK_PP(16'hA3BA,4);
TASK_PP(16'hA3BB,4);
TASK_PP(16'hA3BC,4);
TASK_PP(16'hA3BD,4);
TASK_PP(16'hA3BE,4);
TASK_PP(16'hA3BF,4);
TASK_PP(16'hA3C0,4);
TASK_PP(16'hA3C1,4);
TASK_PP(16'hA3C2,4);
TASK_PP(16'hA3C3,4);
TASK_PP(16'hA3C4,4);
TASK_PP(16'hA3C5,4);
TASK_PP(16'hA3C6,4);
TASK_PP(16'hA3C7,4);
TASK_PP(16'hA3C8,4);
TASK_PP(16'hA3C9,4);
TASK_PP(16'hA3CA,4);
TASK_PP(16'hA3CB,4);
TASK_PP(16'hA3CC,4);
TASK_PP(16'hA3CD,4);
TASK_PP(16'hA3CE,4);
TASK_PP(16'hA3CF,4);
TASK_PP(16'hA3D0,4);
TASK_PP(16'hA3D1,4);
TASK_PP(16'hA3D2,4);
TASK_PP(16'hA3D3,4);
TASK_PP(16'hA3D4,4);
TASK_PP(16'hA3D5,4);
TASK_PP(16'hA3D6,4);
TASK_PP(16'hA3D7,4);
TASK_PP(16'hA3D8,4);
TASK_PP(16'hA3D9,4);
TASK_PP(16'hA3DA,4);
TASK_PP(16'hA3DB,4);
TASK_PP(16'hA3DC,4);
TASK_PP(16'hA3DD,4);
TASK_PP(16'hA3DE,4);
TASK_PP(16'hA3DF,4);
TASK_PP(16'hA3E0,4);
TASK_PP(16'hA3E1,4);
TASK_PP(16'hA3E2,4);
TASK_PP(16'hA3E3,4);
TASK_PP(16'hA3E4,4);
TASK_PP(16'hA3E5,4);
TASK_PP(16'hA3E6,4);
TASK_PP(16'hA3E7,4);
TASK_PP(16'hA3E8,4);
TASK_PP(16'hA3E9,4);
TASK_PP(16'hA3EA,4);
TASK_PP(16'hA3EB,4);
TASK_PP(16'hA3EC,4);
TASK_PP(16'hA3ED,4);
TASK_PP(16'hA3EE,4);
TASK_PP(16'hA3EF,4);
TASK_PP(16'hA3F0,4);
TASK_PP(16'hA3F1,4);
TASK_PP(16'hA3F2,4);
TASK_PP(16'hA3F3,4);
TASK_PP(16'hA3F4,4);
TASK_PP(16'hA3F5,4);
TASK_PP(16'hA3F6,4);
TASK_PP(16'hA3F7,4);
TASK_PP(16'hA3F8,4);
TASK_PP(16'hA3F9,4);
TASK_PP(16'hA3FA,4);
TASK_PP(16'hA3FB,4);
TASK_PP(16'hA3FC,4);
TASK_PP(16'hA3FD,4);
TASK_PP(16'hA3FE,4);
TASK_PP(16'hA3FF,4);
TASK_PP(16'hA400,4);
TASK_PP(16'hA401,4);
TASK_PP(16'hA402,4);
TASK_PP(16'hA403,4);
TASK_PP(16'hA404,4);
TASK_PP(16'hA405,4);
TASK_PP(16'hA406,4);
TASK_PP(16'hA407,4);
TASK_PP(16'hA408,4);
TASK_PP(16'hA409,4);
TASK_PP(16'hA40A,4);
TASK_PP(16'hA40B,4);
TASK_PP(16'hA40C,4);
TASK_PP(16'hA40D,4);
TASK_PP(16'hA40E,4);
TASK_PP(16'hA40F,4);
TASK_PP(16'hA410,4);
TASK_PP(16'hA411,4);
TASK_PP(16'hA412,4);
TASK_PP(16'hA413,4);
TASK_PP(16'hA414,4);
TASK_PP(16'hA415,4);
TASK_PP(16'hA416,4);
TASK_PP(16'hA417,4);
TASK_PP(16'hA418,4);
TASK_PP(16'hA419,4);
TASK_PP(16'hA41A,4);
TASK_PP(16'hA41B,4);
TASK_PP(16'hA41C,4);
TASK_PP(16'hA41D,4);
TASK_PP(16'hA41E,4);
TASK_PP(16'hA41F,4);
TASK_PP(16'hA420,4);
TASK_PP(16'hA421,4);
TASK_PP(16'hA422,4);
TASK_PP(16'hA423,4);
TASK_PP(16'hA424,4);
TASK_PP(16'hA425,4);
TASK_PP(16'hA426,4);
TASK_PP(16'hA427,4);
TASK_PP(16'hA428,4);
TASK_PP(16'hA429,4);
TASK_PP(16'hA42A,4);
TASK_PP(16'hA42B,4);
TASK_PP(16'hA42C,4);
TASK_PP(16'hA42D,4);
TASK_PP(16'hA42E,4);
TASK_PP(16'hA42F,4);
TASK_PP(16'hA430,4);
TASK_PP(16'hA431,4);
TASK_PP(16'hA432,4);
TASK_PP(16'hA433,4);
TASK_PP(16'hA434,4);
TASK_PP(16'hA435,4);
TASK_PP(16'hA436,4);
TASK_PP(16'hA437,4);
TASK_PP(16'hA438,4);
TASK_PP(16'hA439,4);
TASK_PP(16'hA43A,4);
TASK_PP(16'hA43B,4);
TASK_PP(16'hA43C,4);
TASK_PP(16'hA43D,4);
TASK_PP(16'hA43E,4);
TASK_PP(16'hA43F,4);
TASK_PP(16'hA440,4);
TASK_PP(16'hA441,4);
TASK_PP(16'hA442,4);
TASK_PP(16'hA443,4);
TASK_PP(16'hA444,4);
TASK_PP(16'hA445,4);
TASK_PP(16'hA446,4);
TASK_PP(16'hA447,4);
TASK_PP(16'hA448,4);
TASK_PP(16'hA449,4);
TASK_PP(16'hA44A,4);
TASK_PP(16'hA44B,4);
TASK_PP(16'hA44C,4);
TASK_PP(16'hA44D,4);
TASK_PP(16'hA44E,4);
TASK_PP(16'hA44F,4);
TASK_PP(16'hA450,4);
TASK_PP(16'hA451,4);
TASK_PP(16'hA452,4);
TASK_PP(16'hA453,4);
TASK_PP(16'hA454,4);
TASK_PP(16'hA455,4);
TASK_PP(16'hA456,4);
TASK_PP(16'hA457,4);
TASK_PP(16'hA458,4);
TASK_PP(16'hA459,4);
TASK_PP(16'hA45A,4);
TASK_PP(16'hA45B,4);
TASK_PP(16'hA45C,4);
TASK_PP(16'hA45D,4);
TASK_PP(16'hA45E,4);
TASK_PP(16'hA45F,4);
TASK_PP(16'hA460,4);
TASK_PP(16'hA461,4);
TASK_PP(16'hA462,4);
TASK_PP(16'hA463,4);
TASK_PP(16'hA464,4);
TASK_PP(16'hA465,4);
TASK_PP(16'hA466,4);
TASK_PP(16'hA467,4);
TASK_PP(16'hA468,4);
TASK_PP(16'hA469,4);
TASK_PP(16'hA46A,4);
TASK_PP(16'hA46B,4);
TASK_PP(16'hA46C,4);
TASK_PP(16'hA46D,4);
TASK_PP(16'hA46E,4);
TASK_PP(16'hA46F,4);
TASK_PP(16'hA470,4);
TASK_PP(16'hA471,4);
TASK_PP(16'hA472,4);
TASK_PP(16'hA473,4);
TASK_PP(16'hA474,4);
TASK_PP(16'hA475,4);
TASK_PP(16'hA476,4);
TASK_PP(16'hA477,4);
TASK_PP(16'hA478,4);
TASK_PP(16'hA479,4);
TASK_PP(16'hA47A,4);
TASK_PP(16'hA47B,4);
TASK_PP(16'hA47C,4);
TASK_PP(16'hA47D,4);
TASK_PP(16'hA47E,4);
TASK_PP(16'hA47F,4);
TASK_PP(16'hA480,4);
TASK_PP(16'hA481,4);
TASK_PP(16'hA482,4);
TASK_PP(16'hA483,4);
TASK_PP(16'hA484,4);
TASK_PP(16'hA485,4);
TASK_PP(16'hA486,4);
TASK_PP(16'hA487,4);
TASK_PP(16'hA488,4);
TASK_PP(16'hA489,4);
TASK_PP(16'hA48A,4);
TASK_PP(16'hA48B,4);
TASK_PP(16'hA48C,4);
TASK_PP(16'hA48D,4);
TASK_PP(16'hA48E,4);
TASK_PP(16'hA48F,4);
TASK_PP(16'hA490,4);
TASK_PP(16'hA491,4);
TASK_PP(16'hA492,4);
TASK_PP(16'hA493,4);
TASK_PP(16'hA494,4);
TASK_PP(16'hA495,4);
TASK_PP(16'hA496,4);
TASK_PP(16'hA497,4);
TASK_PP(16'hA498,4);
TASK_PP(16'hA499,4);
TASK_PP(16'hA49A,4);
TASK_PP(16'hA49B,4);
TASK_PP(16'hA49C,4);
TASK_PP(16'hA49D,4);
TASK_PP(16'hA49E,4);
TASK_PP(16'hA49F,4);
TASK_PP(16'hA4A0,4);
TASK_PP(16'hA4A1,4);
TASK_PP(16'hA4A2,4);
TASK_PP(16'hA4A3,4);
TASK_PP(16'hA4A4,4);
TASK_PP(16'hA4A5,4);
TASK_PP(16'hA4A6,4);
TASK_PP(16'hA4A7,4);
TASK_PP(16'hA4A8,4);
TASK_PP(16'hA4A9,4);
TASK_PP(16'hA4AA,4);
TASK_PP(16'hA4AB,4);
TASK_PP(16'hA4AC,4);
TASK_PP(16'hA4AD,4);
TASK_PP(16'hA4AE,4);
TASK_PP(16'hA4AF,4);
TASK_PP(16'hA4B0,4);
TASK_PP(16'hA4B1,4);
TASK_PP(16'hA4B2,4);
TASK_PP(16'hA4B3,4);
TASK_PP(16'hA4B4,4);
TASK_PP(16'hA4B5,4);
TASK_PP(16'hA4B6,4);
TASK_PP(16'hA4B7,4);
TASK_PP(16'hA4B8,4);
TASK_PP(16'hA4B9,4);
TASK_PP(16'hA4BA,4);
TASK_PP(16'hA4BB,4);
TASK_PP(16'hA4BC,4);
TASK_PP(16'hA4BD,4);
TASK_PP(16'hA4BE,4);
TASK_PP(16'hA4BF,4);
TASK_PP(16'hA4C0,4);
TASK_PP(16'hA4C1,4);
TASK_PP(16'hA4C2,4);
TASK_PP(16'hA4C3,4);
TASK_PP(16'hA4C4,4);
TASK_PP(16'hA4C5,4);
TASK_PP(16'hA4C6,4);
TASK_PP(16'hA4C7,4);
TASK_PP(16'hA4C8,4);
TASK_PP(16'hA4C9,4);
TASK_PP(16'hA4CA,4);
TASK_PP(16'hA4CB,4);
TASK_PP(16'hA4CC,4);
TASK_PP(16'hA4CD,4);
TASK_PP(16'hA4CE,4);
TASK_PP(16'hA4CF,4);
TASK_PP(16'hA4D0,4);
TASK_PP(16'hA4D1,4);
TASK_PP(16'hA4D2,4);
TASK_PP(16'hA4D3,4);
TASK_PP(16'hA4D4,4);
TASK_PP(16'hA4D5,4);
TASK_PP(16'hA4D6,4);
TASK_PP(16'hA4D7,4);
TASK_PP(16'hA4D8,4);
TASK_PP(16'hA4D9,4);
TASK_PP(16'hA4DA,4);
TASK_PP(16'hA4DB,4);
TASK_PP(16'hA4DC,4);
TASK_PP(16'hA4DD,4);
TASK_PP(16'hA4DE,4);
TASK_PP(16'hA4DF,4);
TASK_PP(16'hA4E0,4);
TASK_PP(16'hA4E1,4);
TASK_PP(16'hA4E2,4);
TASK_PP(16'hA4E3,4);
TASK_PP(16'hA4E4,4);
TASK_PP(16'hA4E5,4);
TASK_PP(16'hA4E6,4);
TASK_PP(16'hA4E7,4);
TASK_PP(16'hA4E8,4);
TASK_PP(16'hA4E9,4);
TASK_PP(16'hA4EA,4);
TASK_PP(16'hA4EB,4);
TASK_PP(16'hA4EC,4);
TASK_PP(16'hA4ED,4);
TASK_PP(16'hA4EE,4);
TASK_PP(16'hA4EF,4);
TASK_PP(16'hA4F0,4);
TASK_PP(16'hA4F1,4);
TASK_PP(16'hA4F2,4);
TASK_PP(16'hA4F3,4);
TASK_PP(16'hA4F4,4);
TASK_PP(16'hA4F5,4);
TASK_PP(16'hA4F6,4);
TASK_PP(16'hA4F7,4);
TASK_PP(16'hA4F8,4);
TASK_PP(16'hA4F9,4);
TASK_PP(16'hA4FA,4);
TASK_PP(16'hA4FB,4);
TASK_PP(16'hA4FC,4);
TASK_PP(16'hA4FD,4);
TASK_PP(16'hA4FE,4);
TASK_PP(16'hA4FF,4);
TASK_PP(16'hA500,4);
TASK_PP(16'hA501,4);
TASK_PP(16'hA502,4);
TASK_PP(16'hA503,4);
TASK_PP(16'hA504,4);
TASK_PP(16'hA505,4);
TASK_PP(16'hA506,4);
TASK_PP(16'hA507,4);
TASK_PP(16'hA508,4);
TASK_PP(16'hA509,4);
TASK_PP(16'hA50A,4);
TASK_PP(16'hA50B,4);
TASK_PP(16'hA50C,4);
TASK_PP(16'hA50D,4);
TASK_PP(16'hA50E,4);
TASK_PP(16'hA50F,4);
TASK_PP(16'hA510,4);
TASK_PP(16'hA511,4);
TASK_PP(16'hA512,4);
TASK_PP(16'hA513,4);
TASK_PP(16'hA514,4);
TASK_PP(16'hA515,4);
TASK_PP(16'hA516,4);
TASK_PP(16'hA517,4);
TASK_PP(16'hA518,4);
TASK_PP(16'hA519,4);
TASK_PP(16'hA51A,4);
TASK_PP(16'hA51B,4);
TASK_PP(16'hA51C,4);
TASK_PP(16'hA51D,4);
TASK_PP(16'hA51E,4);
TASK_PP(16'hA51F,4);
TASK_PP(16'hA520,4);
TASK_PP(16'hA521,4);
TASK_PP(16'hA522,4);
TASK_PP(16'hA523,4);
TASK_PP(16'hA524,4);
TASK_PP(16'hA525,4);
TASK_PP(16'hA526,4);
TASK_PP(16'hA527,4);
TASK_PP(16'hA528,4);
TASK_PP(16'hA529,4);
TASK_PP(16'hA52A,4);
TASK_PP(16'hA52B,4);
TASK_PP(16'hA52C,4);
TASK_PP(16'hA52D,4);
TASK_PP(16'hA52E,4);
TASK_PP(16'hA52F,4);
TASK_PP(16'hA530,4);
TASK_PP(16'hA531,4);
TASK_PP(16'hA532,4);
TASK_PP(16'hA533,4);
TASK_PP(16'hA534,4);
TASK_PP(16'hA535,4);
TASK_PP(16'hA536,4);
TASK_PP(16'hA537,4);
TASK_PP(16'hA538,4);
TASK_PP(16'hA539,4);
TASK_PP(16'hA53A,4);
TASK_PP(16'hA53B,4);
TASK_PP(16'hA53C,4);
TASK_PP(16'hA53D,4);
TASK_PP(16'hA53E,4);
TASK_PP(16'hA53F,4);
TASK_PP(16'hA540,4);
TASK_PP(16'hA541,4);
TASK_PP(16'hA542,4);
TASK_PP(16'hA543,4);
TASK_PP(16'hA544,4);
TASK_PP(16'hA545,4);
TASK_PP(16'hA546,4);
TASK_PP(16'hA547,4);
TASK_PP(16'hA548,4);
TASK_PP(16'hA549,4);
TASK_PP(16'hA54A,4);
TASK_PP(16'hA54B,4);
TASK_PP(16'hA54C,4);
TASK_PP(16'hA54D,4);
TASK_PP(16'hA54E,4);
TASK_PP(16'hA54F,4);
TASK_PP(16'hA550,4);
TASK_PP(16'hA551,4);
TASK_PP(16'hA552,4);
TASK_PP(16'hA553,4);
TASK_PP(16'hA554,4);
TASK_PP(16'hA555,4);
TASK_PP(16'hA556,4);
TASK_PP(16'hA557,4);
TASK_PP(16'hA558,4);
TASK_PP(16'hA559,4);
TASK_PP(16'hA55A,4);
TASK_PP(16'hA55B,4);
TASK_PP(16'hA55C,4);
TASK_PP(16'hA55D,4);
TASK_PP(16'hA55E,4);
TASK_PP(16'hA55F,4);
TASK_PP(16'hA560,4);
TASK_PP(16'hA561,4);
TASK_PP(16'hA562,4);
TASK_PP(16'hA563,4);
TASK_PP(16'hA564,4);
TASK_PP(16'hA565,4);
TASK_PP(16'hA566,4);
TASK_PP(16'hA567,4);
TASK_PP(16'hA568,4);
TASK_PP(16'hA569,4);
TASK_PP(16'hA56A,4);
TASK_PP(16'hA56B,4);
TASK_PP(16'hA56C,4);
TASK_PP(16'hA56D,4);
TASK_PP(16'hA56E,4);
TASK_PP(16'hA56F,4);
TASK_PP(16'hA570,4);
TASK_PP(16'hA571,4);
TASK_PP(16'hA572,4);
TASK_PP(16'hA573,4);
TASK_PP(16'hA574,4);
TASK_PP(16'hA575,4);
TASK_PP(16'hA576,4);
TASK_PP(16'hA577,4);
TASK_PP(16'hA578,4);
TASK_PP(16'hA579,4);
TASK_PP(16'hA57A,4);
TASK_PP(16'hA57B,4);
TASK_PP(16'hA57C,4);
TASK_PP(16'hA57D,4);
TASK_PP(16'hA57E,4);
TASK_PP(16'hA57F,4);
TASK_PP(16'hA580,4);
TASK_PP(16'hA581,4);
TASK_PP(16'hA582,4);
TASK_PP(16'hA583,4);
TASK_PP(16'hA584,4);
TASK_PP(16'hA585,4);
TASK_PP(16'hA586,4);
TASK_PP(16'hA587,4);
TASK_PP(16'hA588,4);
TASK_PP(16'hA589,4);
TASK_PP(16'hA58A,4);
TASK_PP(16'hA58B,4);
TASK_PP(16'hA58C,4);
TASK_PP(16'hA58D,4);
TASK_PP(16'hA58E,4);
TASK_PP(16'hA58F,4);
TASK_PP(16'hA590,4);
TASK_PP(16'hA591,4);
TASK_PP(16'hA592,4);
TASK_PP(16'hA593,4);
TASK_PP(16'hA594,4);
TASK_PP(16'hA595,4);
TASK_PP(16'hA596,4);
TASK_PP(16'hA597,4);
TASK_PP(16'hA598,4);
TASK_PP(16'hA599,4);
TASK_PP(16'hA59A,4);
TASK_PP(16'hA59B,4);
TASK_PP(16'hA59C,4);
TASK_PP(16'hA59D,4);
TASK_PP(16'hA59E,4);
TASK_PP(16'hA59F,4);
TASK_PP(16'hA5A0,4);
TASK_PP(16'hA5A1,4);
TASK_PP(16'hA5A2,4);
TASK_PP(16'hA5A3,4);
TASK_PP(16'hA5A4,4);
TASK_PP(16'hA5A5,4);
TASK_PP(16'hA5A6,4);
TASK_PP(16'hA5A7,4);
TASK_PP(16'hA5A8,4);
TASK_PP(16'hA5A9,4);
TASK_PP(16'hA5AA,4);
TASK_PP(16'hA5AB,4);
TASK_PP(16'hA5AC,4);
TASK_PP(16'hA5AD,4);
TASK_PP(16'hA5AE,4);
TASK_PP(16'hA5AF,4);
TASK_PP(16'hA5B0,4);
TASK_PP(16'hA5B1,4);
TASK_PP(16'hA5B2,4);
TASK_PP(16'hA5B3,4);
TASK_PP(16'hA5B4,4);
TASK_PP(16'hA5B5,4);
TASK_PP(16'hA5B6,4);
TASK_PP(16'hA5B7,4);
TASK_PP(16'hA5B8,4);
TASK_PP(16'hA5B9,4);
TASK_PP(16'hA5BA,4);
TASK_PP(16'hA5BB,4);
TASK_PP(16'hA5BC,4);
TASK_PP(16'hA5BD,4);
TASK_PP(16'hA5BE,4);
TASK_PP(16'hA5BF,4);
TASK_PP(16'hA5C0,4);
TASK_PP(16'hA5C1,4);
TASK_PP(16'hA5C2,4);
TASK_PP(16'hA5C3,4);
TASK_PP(16'hA5C4,4);
TASK_PP(16'hA5C5,4);
TASK_PP(16'hA5C6,4);
TASK_PP(16'hA5C7,4);
TASK_PP(16'hA5C8,4);
TASK_PP(16'hA5C9,4);
TASK_PP(16'hA5CA,4);
TASK_PP(16'hA5CB,4);
TASK_PP(16'hA5CC,4);
TASK_PP(16'hA5CD,4);
TASK_PP(16'hA5CE,4);
TASK_PP(16'hA5CF,4);
TASK_PP(16'hA5D0,4);
TASK_PP(16'hA5D1,4);
TASK_PP(16'hA5D2,4);
TASK_PP(16'hA5D3,4);
TASK_PP(16'hA5D4,4);
TASK_PP(16'hA5D5,4);
TASK_PP(16'hA5D6,4);
TASK_PP(16'hA5D7,4);
TASK_PP(16'hA5D8,4);
TASK_PP(16'hA5D9,4);
TASK_PP(16'hA5DA,4);
TASK_PP(16'hA5DB,4);
TASK_PP(16'hA5DC,4);
TASK_PP(16'hA5DD,4);
TASK_PP(16'hA5DE,4);
TASK_PP(16'hA5DF,4);
TASK_PP(16'hA5E0,4);
TASK_PP(16'hA5E1,4);
TASK_PP(16'hA5E2,4);
TASK_PP(16'hA5E3,4);
TASK_PP(16'hA5E4,4);
TASK_PP(16'hA5E5,4);
TASK_PP(16'hA5E6,4);
TASK_PP(16'hA5E7,4);
TASK_PP(16'hA5E8,4);
TASK_PP(16'hA5E9,4);
TASK_PP(16'hA5EA,4);
TASK_PP(16'hA5EB,4);
TASK_PP(16'hA5EC,4);
TASK_PP(16'hA5ED,4);
TASK_PP(16'hA5EE,4);
TASK_PP(16'hA5EF,4);
TASK_PP(16'hA5F0,4);
TASK_PP(16'hA5F1,4);
TASK_PP(16'hA5F2,4);
TASK_PP(16'hA5F3,4);
TASK_PP(16'hA5F4,4);
TASK_PP(16'hA5F5,4);
TASK_PP(16'hA5F6,4);
TASK_PP(16'hA5F7,4);
TASK_PP(16'hA5F8,4);
TASK_PP(16'hA5F9,4);
TASK_PP(16'hA5FA,4);
TASK_PP(16'hA5FB,4);
TASK_PP(16'hA5FC,4);
TASK_PP(16'hA5FD,4);
TASK_PP(16'hA5FE,4);
TASK_PP(16'hA5FF,4);
TASK_PP(16'hA600,4);
TASK_PP(16'hA601,4);
TASK_PP(16'hA602,4);
TASK_PP(16'hA603,4);
TASK_PP(16'hA604,4);
TASK_PP(16'hA605,4);
TASK_PP(16'hA606,4);
TASK_PP(16'hA607,4);
TASK_PP(16'hA608,4);
TASK_PP(16'hA609,4);
TASK_PP(16'hA60A,4);
TASK_PP(16'hA60B,4);
TASK_PP(16'hA60C,4);
TASK_PP(16'hA60D,4);
TASK_PP(16'hA60E,4);
TASK_PP(16'hA60F,4);
TASK_PP(16'hA610,4);
TASK_PP(16'hA611,4);
TASK_PP(16'hA612,4);
TASK_PP(16'hA613,4);
TASK_PP(16'hA614,4);
TASK_PP(16'hA615,4);
TASK_PP(16'hA616,4);
TASK_PP(16'hA617,4);
TASK_PP(16'hA618,4);
TASK_PP(16'hA619,4);
TASK_PP(16'hA61A,4);
TASK_PP(16'hA61B,4);
TASK_PP(16'hA61C,4);
TASK_PP(16'hA61D,4);
TASK_PP(16'hA61E,4);
TASK_PP(16'hA61F,4);
TASK_PP(16'hA620,4);
TASK_PP(16'hA621,4);
TASK_PP(16'hA622,4);
TASK_PP(16'hA623,4);
TASK_PP(16'hA624,4);
TASK_PP(16'hA625,4);
TASK_PP(16'hA626,4);
TASK_PP(16'hA627,4);
TASK_PP(16'hA628,4);
TASK_PP(16'hA629,4);
TASK_PP(16'hA62A,4);
TASK_PP(16'hA62B,4);
TASK_PP(16'hA62C,4);
TASK_PP(16'hA62D,4);
TASK_PP(16'hA62E,4);
TASK_PP(16'hA62F,4);
TASK_PP(16'hA630,4);
TASK_PP(16'hA631,4);
TASK_PP(16'hA632,4);
TASK_PP(16'hA633,4);
TASK_PP(16'hA634,4);
TASK_PP(16'hA635,4);
TASK_PP(16'hA636,4);
TASK_PP(16'hA637,4);
TASK_PP(16'hA638,4);
TASK_PP(16'hA639,4);
TASK_PP(16'hA63A,4);
TASK_PP(16'hA63B,4);
TASK_PP(16'hA63C,4);
TASK_PP(16'hA63D,4);
TASK_PP(16'hA63E,4);
TASK_PP(16'hA63F,4);
TASK_PP(16'hA640,4);
TASK_PP(16'hA641,4);
TASK_PP(16'hA642,4);
TASK_PP(16'hA643,4);
TASK_PP(16'hA644,4);
TASK_PP(16'hA645,4);
TASK_PP(16'hA646,4);
TASK_PP(16'hA647,4);
TASK_PP(16'hA648,4);
TASK_PP(16'hA649,4);
TASK_PP(16'hA64A,4);
TASK_PP(16'hA64B,4);
TASK_PP(16'hA64C,4);
TASK_PP(16'hA64D,4);
TASK_PP(16'hA64E,4);
TASK_PP(16'hA64F,4);
TASK_PP(16'hA650,4);
TASK_PP(16'hA651,4);
TASK_PP(16'hA652,4);
TASK_PP(16'hA653,4);
TASK_PP(16'hA654,4);
TASK_PP(16'hA655,4);
TASK_PP(16'hA656,4);
TASK_PP(16'hA657,4);
TASK_PP(16'hA658,4);
TASK_PP(16'hA659,4);
TASK_PP(16'hA65A,4);
TASK_PP(16'hA65B,4);
TASK_PP(16'hA65C,4);
TASK_PP(16'hA65D,4);
TASK_PP(16'hA65E,4);
TASK_PP(16'hA65F,4);
TASK_PP(16'hA660,4);
TASK_PP(16'hA661,4);
TASK_PP(16'hA662,4);
TASK_PP(16'hA663,4);
TASK_PP(16'hA664,4);
TASK_PP(16'hA665,4);
TASK_PP(16'hA666,4);
TASK_PP(16'hA667,4);
TASK_PP(16'hA668,4);
TASK_PP(16'hA669,4);
TASK_PP(16'hA66A,4);
TASK_PP(16'hA66B,4);
TASK_PP(16'hA66C,4);
TASK_PP(16'hA66D,4);
TASK_PP(16'hA66E,4);
TASK_PP(16'hA66F,4);
TASK_PP(16'hA670,4);
TASK_PP(16'hA671,4);
TASK_PP(16'hA672,4);
TASK_PP(16'hA673,4);
TASK_PP(16'hA674,4);
TASK_PP(16'hA675,4);
TASK_PP(16'hA676,4);
TASK_PP(16'hA677,4);
TASK_PP(16'hA678,4);
TASK_PP(16'hA679,4);
TASK_PP(16'hA67A,4);
TASK_PP(16'hA67B,4);
TASK_PP(16'hA67C,4);
TASK_PP(16'hA67D,4);
TASK_PP(16'hA67E,4);
TASK_PP(16'hA67F,4);
TASK_PP(16'hA680,4);
TASK_PP(16'hA681,4);
TASK_PP(16'hA682,4);
TASK_PP(16'hA683,4);
TASK_PP(16'hA684,4);
TASK_PP(16'hA685,4);
TASK_PP(16'hA686,4);
TASK_PP(16'hA687,4);
TASK_PP(16'hA688,4);
TASK_PP(16'hA689,4);
TASK_PP(16'hA68A,4);
TASK_PP(16'hA68B,4);
TASK_PP(16'hA68C,4);
TASK_PP(16'hA68D,4);
TASK_PP(16'hA68E,4);
TASK_PP(16'hA68F,4);
TASK_PP(16'hA690,4);
TASK_PP(16'hA691,4);
TASK_PP(16'hA692,4);
TASK_PP(16'hA693,4);
TASK_PP(16'hA694,4);
TASK_PP(16'hA695,4);
TASK_PP(16'hA696,4);
TASK_PP(16'hA697,4);
TASK_PP(16'hA698,4);
TASK_PP(16'hA699,4);
TASK_PP(16'hA69A,4);
TASK_PP(16'hA69B,4);
TASK_PP(16'hA69C,4);
TASK_PP(16'hA69D,4);
TASK_PP(16'hA69E,4);
TASK_PP(16'hA69F,4);
TASK_PP(16'hA6A0,4);
TASK_PP(16'hA6A1,4);
TASK_PP(16'hA6A2,4);
TASK_PP(16'hA6A3,4);
TASK_PP(16'hA6A4,4);
TASK_PP(16'hA6A5,4);
TASK_PP(16'hA6A6,4);
TASK_PP(16'hA6A7,4);
TASK_PP(16'hA6A8,4);
TASK_PP(16'hA6A9,4);
TASK_PP(16'hA6AA,4);
TASK_PP(16'hA6AB,4);
TASK_PP(16'hA6AC,4);
TASK_PP(16'hA6AD,4);
TASK_PP(16'hA6AE,4);
TASK_PP(16'hA6AF,4);
TASK_PP(16'hA6B0,4);
TASK_PP(16'hA6B1,4);
TASK_PP(16'hA6B2,4);
TASK_PP(16'hA6B3,4);
TASK_PP(16'hA6B4,4);
TASK_PP(16'hA6B5,4);
TASK_PP(16'hA6B6,4);
TASK_PP(16'hA6B7,4);
TASK_PP(16'hA6B8,4);
TASK_PP(16'hA6B9,4);
TASK_PP(16'hA6BA,4);
TASK_PP(16'hA6BB,4);
TASK_PP(16'hA6BC,4);
TASK_PP(16'hA6BD,4);
TASK_PP(16'hA6BE,4);
TASK_PP(16'hA6BF,4);
TASK_PP(16'hA6C0,4);
TASK_PP(16'hA6C1,4);
TASK_PP(16'hA6C2,4);
TASK_PP(16'hA6C3,4);
TASK_PP(16'hA6C4,4);
TASK_PP(16'hA6C5,4);
TASK_PP(16'hA6C6,4);
TASK_PP(16'hA6C7,4);
TASK_PP(16'hA6C8,4);
TASK_PP(16'hA6C9,4);
TASK_PP(16'hA6CA,4);
TASK_PP(16'hA6CB,4);
TASK_PP(16'hA6CC,4);
TASK_PP(16'hA6CD,4);
TASK_PP(16'hA6CE,4);
TASK_PP(16'hA6CF,4);
TASK_PP(16'hA6D0,4);
TASK_PP(16'hA6D1,4);
TASK_PP(16'hA6D2,4);
TASK_PP(16'hA6D3,4);
TASK_PP(16'hA6D4,4);
TASK_PP(16'hA6D5,4);
TASK_PP(16'hA6D6,4);
TASK_PP(16'hA6D7,4);
TASK_PP(16'hA6D8,4);
TASK_PP(16'hA6D9,4);
TASK_PP(16'hA6DA,4);
TASK_PP(16'hA6DB,4);
TASK_PP(16'hA6DC,4);
TASK_PP(16'hA6DD,4);
TASK_PP(16'hA6DE,4);
TASK_PP(16'hA6DF,4);
TASK_PP(16'hA6E0,4);
TASK_PP(16'hA6E1,4);
TASK_PP(16'hA6E2,4);
TASK_PP(16'hA6E3,4);
TASK_PP(16'hA6E4,4);
TASK_PP(16'hA6E5,4);
TASK_PP(16'hA6E6,4);
TASK_PP(16'hA6E7,4);
TASK_PP(16'hA6E8,4);
TASK_PP(16'hA6E9,4);
TASK_PP(16'hA6EA,4);
TASK_PP(16'hA6EB,4);
TASK_PP(16'hA6EC,4);
TASK_PP(16'hA6ED,4);
TASK_PP(16'hA6EE,4);
TASK_PP(16'hA6EF,4);
TASK_PP(16'hA6F0,4);
TASK_PP(16'hA6F1,4);
TASK_PP(16'hA6F2,4);
TASK_PP(16'hA6F3,4);
TASK_PP(16'hA6F4,4);
TASK_PP(16'hA6F5,4);
TASK_PP(16'hA6F6,4);
TASK_PP(16'hA6F7,4);
TASK_PP(16'hA6F8,4);
TASK_PP(16'hA6F9,4);
TASK_PP(16'hA6FA,4);
TASK_PP(16'hA6FB,4);
TASK_PP(16'hA6FC,4);
TASK_PP(16'hA6FD,4);
TASK_PP(16'hA6FE,4);
TASK_PP(16'hA6FF,4);
TASK_PP(16'hA700,4);
TASK_PP(16'hA701,4);
TASK_PP(16'hA702,4);
TASK_PP(16'hA703,4);
TASK_PP(16'hA704,4);
TASK_PP(16'hA705,4);
TASK_PP(16'hA706,4);
TASK_PP(16'hA707,4);
TASK_PP(16'hA708,4);
TASK_PP(16'hA709,4);
TASK_PP(16'hA70A,4);
TASK_PP(16'hA70B,4);
TASK_PP(16'hA70C,4);
TASK_PP(16'hA70D,4);
TASK_PP(16'hA70E,4);
TASK_PP(16'hA70F,4);
TASK_PP(16'hA710,4);
TASK_PP(16'hA711,4);
TASK_PP(16'hA712,4);
TASK_PP(16'hA713,4);
TASK_PP(16'hA714,4);
TASK_PP(16'hA715,4);
TASK_PP(16'hA716,4);
TASK_PP(16'hA717,4);
TASK_PP(16'hA718,4);
TASK_PP(16'hA719,4);
TASK_PP(16'hA71A,4);
TASK_PP(16'hA71B,4);
TASK_PP(16'hA71C,4);
TASK_PP(16'hA71D,4);
TASK_PP(16'hA71E,4);
TASK_PP(16'hA71F,4);
TASK_PP(16'hA720,4);
TASK_PP(16'hA721,4);
TASK_PP(16'hA722,4);
TASK_PP(16'hA723,4);
TASK_PP(16'hA724,4);
TASK_PP(16'hA725,4);
TASK_PP(16'hA726,4);
TASK_PP(16'hA727,4);
TASK_PP(16'hA728,4);
TASK_PP(16'hA729,4);
TASK_PP(16'hA72A,4);
TASK_PP(16'hA72B,4);
TASK_PP(16'hA72C,4);
TASK_PP(16'hA72D,4);
TASK_PP(16'hA72E,4);
TASK_PP(16'hA72F,4);
TASK_PP(16'hA730,4);
TASK_PP(16'hA731,4);
TASK_PP(16'hA732,4);
TASK_PP(16'hA733,4);
TASK_PP(16'hA734,4);
TASK_PP(16'hA735,4);
TASK_PP(16'hA736,4);
TASK_PP(16'hA737,4);
TASK_PP(16'hA738,4);
TASK_PP(16'hA739,4);
TASK_PP(16'hA73A,4);
TASK_PP(16'hA73B,4);
TASK_PP(16'hA73C,4);
TASK_PP(16'hA73D,4);
TASK_PP(16'hA73E,4);
TASK_PP(16'hA73F,4);
TASK_PP(16'hA740,4);
TASK_PP(16'hA741,4);
TASK_PP(16'hA742,4);
TASK_PP(16'hA743,4);
TASK_PP(16'hA744,4);
TASK_PP(16'hA745,4);
TASK_PP(16'hA746,4);
TASK_PP(16'hA747,4);
TASK_PP(16'hA748,4);
TASK_PP(16'hA749,4);
TASK_PP(16'hA74A,4);
TASK_PP(16'hA74B,4);
TASK_PP(16'hA74C,4);
TASK_PP(16'hA74D,4);
TASK_PP(16'hA74E,4);
TASK_PP(16'hA74F,4);
TASK_PP(16'hA750,4);
TASK_PP(16'hA751,4);
TASK_PP(16'hA752,4);
TASK_PP(16'hA753,4);
TASK_PP(16'hA754,4);
TASK_PP(16'hA755,4);
TASK_PP(16'hA756,4);
TASK_PP(16'hA757,4);
TASK_PP(16'hA758,4);
TASK_PP(16'hA759,4);
TASK_PP(16'hA75A,4);
TASK_PP(16'hA75B,4);
TASK_PP(16'hA75C,4);
TASK_PP(16'hA75D,4);
TASK_PP(16'hA75E,4);
TASK_PP(16'hA75F,4);
TASK_PP(16'hA760,4);
TASK_PP(16'hA761,4);
TASK_PP(16'hA762,4);
TASK_PP(16'hA763,4);
TASK_PP(16'hA764,4);
TASK_PP(16'hA765,4);
TASK_PP(16'hA766,4);
TASK_PP(16'hA767,4);
TASK_PP(16'hA768,4);
TASK_PP(16'hA769,4);
TASK_PP(16'hA76A,4);
TASK_PP(16'hA76B,4);
TASK_PP(16'hA76C,4);
TASK_PP(16'hA76D,4);
TASK_PP(16'hA76E,4);
TASK_PP(16'hA76F,4);
TASK_PP(16'hA770,4);
TASK_PP(16'hA771,4);
TASK_PP(16'hA772,4);
TASK_PP(16'hA773,4);
TASK_PP(16'hA774,4);
TASK_PP(16'hA775,4);
TASK_PP(16'hA776,4);
TASK_PP(16'hA777,4);
TASK_PP(16'hA778,4);
TASK_PP(16'hA779,4);
TASK_PP(16'hA77A,4);
TASK_PP(16'hA77B,4);
TASK_PP(16'hA77C,4);
TASK_PP(16'hA77D,4);
TASK_PP(16'hA77E,4);
TASK_PP(16'hA77F,4);
TASK_PP(16'hA780,4);
TASK_PP(16'hA781,4);
TASK_PP(16'hA782,4);
TASK_PP(16'hA783,4);
TASK_PP(16'hA784,4);
TASK_PP(16'hA785,4);
TASK_PP(16'hA786,4);
TASK_PP(16'hA787,4);
TASK_PP(16'hA788,4);
TASK_PP(16'hA789,4);
TASK_PP(16'hA78A,4);
TASK_PP(16'hA78B,4);
TASK_PP(16'hA78C,4);
TASK_PP(16'hA78D,4);
TASK_PP(16'hA78E,4);
TASK_PP(16'hA78F,4);
TASK_PP(16'hA790,4);
TASK_PP(16'hA791,4);
TASK_PP(16'hA792,4);
TASK_PP(16'hA793,4);
TASK_PP(16'hA794,4);
TASK_PP(16'hA795,4);
TASK_PP(16'hA796,4);
TASK_PP(16'hA797,4);
TASK_PP(16'hA798,4);
TASK_PP(16'hA799,4);
TASK_PP(16'hA79A,4);
TASK_PP(16'hA79B,4);
TASK_PP(16'hA79C,4);
TASK_PP(16'hA79D,4);
TASK_PP(16'hA79E,4);
TASK_PP(16'hA79F,4);
TASK_PP(16'hA7A0,4);
TASK_PP(16'hA7A1,4);
TASK_PP(16'hA7A2,4);
TASK_PP(16'hA7A3,4);
TASK_PP(16'hA7A4,4);
TASK_PP(16'hA7A5,4);
TASK_PP(16'hA7A6,4);
TASK_PP(16'hA7A7,4);
TASK_PP(16'hA7A8,4);
TASK_PP(16'hA7A9,4);
TASK_PP(16'hA7AA,4);
TASK_PP(16'hA7AB,4);
TASK_PP(16'hA7AC,4);
TASK_PP(16'hA7AD,4);
TASK_PP(16'hA7AE,4);
TASK_PP(16'hA7AF,4);
TASK_PP(16'hA7B0,4);
TASK_PP(16'hA7B1,4);
TASK_PP(16'hA7B2,4);
TASK_PP(16'hA7B3,4);
TASK_PP(16'hA7B4,4);
TASK_PP(16'hA7B5,4);
TASK_PP(16'hA7B6,4);
TASK_PP(16'hA7B7,4);
TASK_PP(16'hA7B8,4);
TASK_PP(16'hA7B9,4);
TASK_PP(16'hA7BA,4);
TASK_PP(16'hA7BB,4);
TASK_PP(16'hA7BC,4);
TASK_PP(16'hA7BD,4);
TASK_PP(16'hA7BE,4);
TASK_PP(16'hA7BF,4);
TASK_PP(16'hA7C0,4);
TASK_PP(16'hA7C1,4);
TASK_PP(16'hA7C2,4);
TASK_PP(16'hA7C3,4);
TASK_PP(16'hA7C4,4);
TASK_PP(16'hA7C5,4);
TASK_PP(16'hA7C6,4);
TASK_PP(16'hA7C7,4);
TASK_PP(16'hA7C8,4);
TASK_PP(16'hA7C9,4);
TASK_PP(16'hA7CA,4);
TASK_PP(16'hA7CB,4);
TASK_PP(16'hA7CC,4);
TASK_PP(16'hA7CD,4);
TASK_PP(16'hA7CE,4);
TASK_PP(16'hA7CF,4);
TASK_PP(16'hA7D0,4);
TASK_PP(16'hA7D1,4);
TASK_PP(16'hA7D2,4);
TASK_PP(16'hA7D3,4);
TASK_PP(16'hA7D4,4);
TASK_PP(16'hA7D5,4);
TASK_PP(16'hA7D6,4);
TASK_PP(16'hA7D7,4);
TASK_PP(16'hA7D8,4);
TASK_PP(16'hA7D9,4);
TASK_PP(16'hA7DA,4);
TASK_PP(16'hA7DB,4);
TASK_PP(16'hA7DC,4);
TASK_PP(16'hA7DD,4);
TASK_PP(16'hA7DE,4);
TASK_PP(16'hA7DF,4);
TASK_PP(16'hA7E0,4);
TASK_PP(16'hA7E1,4);
TASK_PP(16'hA7E2,4);
TASK_PP(16'hA7E3,4);
TASK_PP(16'hA7E4,4);
TASK_PP(16'hA7E5,4);
TASK_PP(16'hA7E6,4);
TASK_PP(16'hA7E7,4);
TASK_PP(16'hA7E8,4);
TASK_PP(16'hA7E9,4);
TASK_PP(16'hA7EA,4);
TASK_PP(16'hA7EB,4);
TASK_PP(16'hA7EC,4);
TASK_PP(16'hA7ED,4);
TASK_PP(16'hA7EE,4);
TASK_PP(16'hA7EF,4);
TASK_PP(16'hA7F0,4);
TASK_PP(16'hA7F1,4);
TASK_PP(16'hA7F2,4);
TASK_PP(16'hA7F3,4);
TASK_PP(16'hA7F4,4);
TASK_PP(16'hA7F5,4);
TASK_PP(16'hA7F6,4);
TASK_PP(16'hA7F7,4);
TASK_PP(16'hA7F8,4);
TASK_PP(16'hA7F9,4);
TASK_PP(16'hA7FA,4);
TASK_PP(16'hA7FB,4);
TASK_PP(16'hA7FC,4);
TASK_PP(16'hA7FD,4);
TASK_PP(16'hA7FE,4);
TASK_PP(16'hA7FF,4);
TASK_PP(16'hA800,4);
TASK_PP(16'hA801,4);
TASK_PP(16'hA802,4);
TASK_PP(16'hA803,4);
TASK_PP(16'hA804,4);
TASK_PP(16'hA805,4);
TASK_PP(16'hA806,4);
TASK_PP(16'hA807,4);
TASK_PP(16'hA808,4);
TASK_PP(16'hA809,4);
TASK_PP(16'hA80A,4);
TASK_PP(16'hA80B,4);
TASK_PP(16'hA80C,4);
TASK_PP(16'hA80D,4);
TASK_PP(16'hA80E,4);
TASK_PP(16'hA80F,4);
TASK_PP(16'hA810,4);
TASK_PP(16'hA811,4);
TASK_PP(16'hA812,4);
TASK_PP(16'hA813,4);
TASK_PP(16'hA814,4);
TASK_PP(16'hA815,4);
TASK_PP(16'hA816,4);
TASK_PP(16'hA817,4);
TASK_PP(16'hA818,4);
TASK_PP(16'hA819,4);
TASK_PP(16'hA81A,4);
TASK_PP(16'hA81B,4);
TASK_PP(16'hA81C,4);
TASK_PP(16'hA81D,4);
TASK_PP(16'hA81E,4);
TASK_PP(16'hA81F,4);
TASK_PP(16'hA820,4);
TASK_PP(16'hA821,4);
TASK_PP(16'hA822,4);
TASK_PP(16'hA823,4);
TASK_PP(16'hA824,4);
TASK_PP(16'hA825,4);
TASK_PP(16'hA826,4);
TASK_PP(16'hA827,4);
TASK_PP(16'hA828,4);
TASK_PP(16'hA829,4);
TASK_PP(16'hA82A,4);
TASK_PP(16'hA82B,4);
TASK_PP(16'hA82C,4);
TASK_PP(16'hA82D,4);
TASK_PP(16'hA82E,4);
TASK_PP(16'hA82F,4);
TASK_PP(16'hA830,4);
TASK_PP(16'hA831,4);
TASK_PP(16'hA832,4);
TASK_PP(16'hA833,4);
TASK_PP(16'hA834,4);
TASK_PP(16'hA835,4);
TASK_PP(16'hA836,4);
TASK_PP(16'hA837,4);
TASK_PP(16'hA838,4);
TASK_PP(16'hA839,4);
TASK_PP(16'hA83A,4);
TASK_PP(16'hA83B,4);
TASK_PP(16'hA83C,4);
TASK_PP(16'hA83D,4);
TASK_PP(16'hA83E,4);
TASK_PP(16'hA83F,4);
TASK_PP(16'hA840,4);
TASK_PP(16'hA841,4);
TASK_PP(16'hA842,4);
TASK_PP(16'hA843,4);
TASK_PP(16'hA844,4);
TASK_PP(16'hA845,4);
TASK_PP(16'hA846,4);
TASK_PP(16'hA847,4);
TASK_PP(16'hA848,4);
TASK_PP(16'hA849,4);
TASK_PP(16'hA84A,4);
TASK_PP(16'hA84B,4);
TASK_PP(16'hA84C,4);
TASK_PP(16'hA84D,4);
TASK_PP(16'hA84E,4);
TASK_PP(16'hA84F,4);
TASK_PP(16'hA850,4);
TASK_PP(16'hA851,4);
TASK_PP(16'hA852,4);
TASK_PP(16'hA853,4);
TASK_PP(16'hA854,4);
TASK_PP(16'hA855,4);
TASK_PP(16'hA856,4);
TASK_PP(16'hA857,4);
TASK_PP(16'hA858,4);
TASK_PP(16'hA859,4);
TASK_PP(16'hA85A,4);
TASK_PP(16'hA85B,4);
TASK_PP(16'hA85C,4);
TASK_PP(16'hA85D,4);
TASK_PP(16'hA85E,4);
TASK_PP(16'hA85F,4);
TASK_PP(16'hA860,4);
TASK_PP(16'hA861,4);
TASK_PP(16'hA862,4);
TASK_PP(16'hA863,4);
TASK_PP(16'hA864,4);
TASK_PP(16'hA865,4);
TASK_PP(16'hA866,4);
TASK_PP(16'hA867,4);
TASK_PP(16'hA868,4);
TASK_PP(16'hA869,4);
TASK_PP(16'hA86A,4);
TASK_PP(16'hA86B,4);
TASK_PP(16'hA86C,4);
TASK_PP(16'hA86D,4);
TASK_PP(16'hA86E,4);
TASK_PP(16'hA86F,4);
TASK_PP(16'hA870,4);
TASK_PP(16'hA871,4);
TASK_PP(16'hA872,4);
TASK_PP(16'hA873,4);
TASK_PP(16'hA874,4);
TASK_PP(16'hA875,4);
TASK_PP(16'hA876,4);
TASK_PP(16'hA877,4);
TASK_PP(16'hA878,4);
TASK_PP(16'hA879,4);
TASK_PP(16'hA87A,4);
TASK_PP(16'hA87B,4);
TASK_PP(16'hA87C,4);
TASK_PP(16'hA87D,4);
TASK_PP(16'hA87E,4);
TASK_PP(16'hA87F,4);
TASK_PP(16'hA880,4);
TASK_PP(16'hA881,4);
TASK_PP(16'hA882,4);
TASK_PP(16'hA883,4);
TASK_PP(16'hA884,4);
TASK_PP(16'hA885,4);
TASK_PP(16'hA886,4);
TASK_PP(16'hA887,4);
TASK_PP(16'hA888,4);
TASK_PP(16'hA889,4);
TASK_PP(16'hA88A,4);
TASK_PP(16'hA88B,4);
TASK_PP(16'hA88C,4);
TASK_PP(16'hA88D,4);
TASK_PP(16'hA88E,4);
TASK_PP(16'hA88F,4);
TASK_PP(16'hA890,4);
TASK_PP(16'hA891,4);
TASK_PP(16'hA892,4);
TASK_PP(16'hA893,4);
TASK_PP(16'hA894,4);
TASK_PP(16'hA895,4);
TASK_PP(16'hA896,4);
TASK_PP(16'hA897,4);
TASK_PP(16'hA898,4);
TASK_PP(16'hA899,4);
TASK_PP(16'hA89A,4);
TASK_PP(16'hA89B,4);
TASK_PP(16'hA89C,4);
TASK_PP(16'hA89D,4);
TASK_PP(16'hA89E,4);
TASK_PP(16'hA89F,4);
TASK_PP(16'hA8A0,4);
TASK_PP(16'hA8A1,4);
TASK_PP(16'hA8A2,4);
TASK_PP(16'hA8A3,4);
TASK_PP(16'hA8A4,4);
TASK_PP(16'hA8A5,4);
TASK_PP(16'hA8A6,4);
TASK_PP(16'hA8A7,4);
TASK_PP(16'hA8A8,4);
TASK_PP(16'hA8A9,4);
TASK_PP(16'hA8AA,4);
TASK_PP(16'hA8AB,4);
TASK_PP(16'hA8AC,4);
TASK_PP(16'hA8AD,4);
TASK_PP(16'hA8AE,4);
TASK_PP(16'hA8AF,4);
TASK_PP(16'hA8B0,4);
TASK_PP(16'hA8B1,4);
TASK_PP(16'hA8B2,4);
TASK_PP(16'hA8B3,4);
TASK_PP(16'hA8B4,4);
TASK_PP(16'hA8B5,4);
TASK_PP(16'hA8B6,4);
TASK_PP(16'hA8B7,4);
TASK_PP(16'hA8B8,4);
TASK_PP(16'hA8B9,4);
TASK_PP(16'hA8BA,4);
TASK_PP(16'hA8BB,4);
TASK_PP(16'hA8BC,4);
TASK_PP(16'hA8BD,4);
TASK_PP(16'hA8BE,4);
TASK_PP(16'hA8BF,4);
TASK_PP(16'hA8C0,4);
TASK_PP(16'hA8C1,4);
TASK_PP(16'hA8C2,4);
TASK_PP(16'hA8C3,4);
TASK_PP(16'hA8C4,4);
TASK_PP(16'hA8C5,4);
TASK_PP(16'hA8C6,4);
TASK_PP(16'hA8C7,4);
TASK_PP(16'hA8C8,4);
TASK_PP(16'hA8C9,4);
TASK_PP(16'hA8CA,4);
TASK_PP(16'hA8CB,4);
TASK_PP(16'hA8CC,4);
TASK_PP(16'hA8CD,4);
TASK_PP(16'hA8CE,4);
TASK_PP(16'hA8CF,4);
TASK_PP(16'hA8D0,4);
TASK_PP(16'hA8D1,4);
TASK_PP(16'hA8D2,4);
TASK_PP(16'hA8D3,4);
TASK_PP(16'hA8D4,4);
TASK_PP(16'hA8D5,4);
TASK_PP(16'hA8D6,4);
TASK_PP(16'hA8D7,4);
TASK_PP(16'hA8D8,4);
TASK_PP(16'hA8D9,4);
TASK_PP(16'hA8DA,4);
TASK_PP(16'hA8DB,4);
TASK_PP(16'hA8DC,4);
TASK_PP(16'hA8DD,4);
TASK_PP(16'hA8DE,4);
TASK_PP(16'hA8DF,4);
TASK_PP(16'hA8E0,4);
TASK_PP(16'hA8E1,4);
TASK_PP(16'hA8E2,4);
TASK_PP(16'hA8E3,4);
TASK_PP(16'hA8E4,4);
TASK_PP(16'hA8E5,4);
TASK_PP(16'hA8E6,4);
TASK_PP(16'hA8E7,4);
TASK_PP(16'hA8E8,4);
TASK_PP(16'hA8E9,4);
TASK_PP(16'hA8EA,4);
TASK_PP(16'hA8EB,4);
TASK_PP(16'hA8EC,4);
TASK_PP(16'hA8ED,4);
TASK_PP(16'hA8EE,4);
TASK_PP(16'hA8EF,4);
TASK_PP(16'hA8F0,4);
TASK_PP(16'hA8F1,4);
TASK_PP(16'hA8F2,4);
TASK_PP(16'hA8F3,4);
TASK_PP(16'hA8F4,4);
TASK_PP(16'hA8F5,4);
TASK_PP(16'hA8F6,4);
TASK_PP(16'hA8F7,4);
TASK_PP(16'hA8F8,4);
TASK_PP(16'hA8F9,4);
TASK_PP(16'hA8FA,4);
TASK_PP(16'hA8FB,4);
TASK_PP(16'hA8FC,4);
TASK_PP(16'hA8FD,4);
TASK_PP(16'hA8FE,4);
TASK_PP(16'hA8FF,4);
TASK_PP(16'hA900,4);
TASK_PP(16'hA901,4);
TASK_PP(16'hA902,4);
TASK_PP(16'hA903,4);
TASK_PP(16'hA904,4);
TASK_PP(16'hA905,4);
TASK_PP(16'hA906,4);
TASK_PP(16'hA907,4);
TASK_PP(16'hA908,4);
TASK_PP(16'hA909,4);
TASK_PP(16'hA90A,4);
TASK_PP(16'hA90B,4);
TASK_PP(16'hA90C,4);
TASK_PP(16'hA90D,4);
TASK_PP(16'hA90E,4);
TASK_PP(16'hA90F,4);
TASK_PP(16'hA910,4);
TASK_PP(16'hA911,4);
TASK_PP(16'hA912,4);
TASK_PP(16'hA913,4);
TASK_PP(16'hA914,4);
TASK_PP(16'hA915,4);
TASK_PP(16'hA916,4);
TASK_PP(16'hA917,4);
TASK_PP(16'hA918,4);
TASK_PP(16'hA919,4);
TASK_PP(16'hA91A,4);
TASK_PP(16'hA91B,4);
TASK_PP(16'hA91C,4);
TASK_PP(16'hA91D,4);
TASK_PP(16'hA91E,4);
TASK_PP(16'hA91F,4);
TASK_PP(16'hA920,4);
TASK_PP(16'hA921,4);
TASK_PP(16'hA922,4);
TASK_PP(16'hA923,4);
TASK_PP(16'hA924,4);
TASK_PP(16'hA925,4);
TASK_PP(16'hA926,4);
TASK_PP(16'hA927,4);
TASK_PP(16'hA928,4);
TASK_PP(16'hA929,4);
TASK_PP(16'hA92A,4);
TASK_PP(16'hA92B,4);
TASK_PP(16'hA92C,4);
TASK_PP(16'hA92D,4);
TASK_PP(16'hA92E,4);
TASK_PP(16'hA92F,4);
TASK_PP(16'hA930,4);
TASK_PP(16'hA931,4);
TASK_PP(16'hA932,4);
TASK_PP(16'hA933,4);
TASK_PP(16'hA934,4);
TASK_PP(16'hA935,4);
TASK_PP(16'hA936,4);
TASK_PP(16'hA937,4);
TASK_PP(16'hA938,4);
TASK_PP(16'hA939,4);
TASK_PP(16'hA93A,4);
TASK_PP(16'hA93B,4);
TASK_PP(16'hA93C,4);
TASK_PP(16'hA93D,4);
TASK_PP(16'hA93E,4);
TASK_PP(16'hA93F,4);
TASK_PP(16'hA940,4);
TASK_PP(16'hA941,4);
TASK_PP(16'hA942,4);
TASK_PP(16'hA943,4);
TASK_PP(16'hA944,4);
TASK_PP(16'hA945,4);
TASK_PP(16'hA946,4);
TASK_PP(16'hA947,4);
TASK_PP(16'hA948,4);
TASK_PP(16'hA949,4);
TASK_PP(16'hA94A,4);
TASK_PP(16'hA94B,4);
TASK_PP(16'hA94C,4);
TASK_PP(16'hA94D,4);
TASK_PP(16'hA94E,4);
TASK_PP(16'hA94F,4);
TASK_PP(16'hA950,4);
TASK_PP(16'hA951,4);
TASK_PP(16'hA952,4);
TASK_PP(16'hA953,4);
TASK_PP(16'hA954,4);
TASK_PP(16'hA955,4);
TASK_PP(16'hA956,4);
TASK_PP(16'hA957,4);
TASK_PP(16'hA958,4);
TASK_PP(16'hA959,4);
TASK_PP(16'hA95A,4);
TASK_PP(16'hA95B,4);
TASK_PP(16'hA95C,4);
TASK_PP(16'hA95D,4);
TASK_PP(16'hA95E,4);
TASK_PP(16'hA95F,4);
TASK_PP(16'hA960,4);
TASK_PP(16'hA961,4);
TASK_PP(16'hA962,4);
TASK_PP(16'hA963,4);
TASK_PP(16'hA964,4);
TASK_PP(16'hA965,4);
TASK_PP(16'hA966,4);
TASK_PP(16'hA967,4);
TASK_PP(16'hA968,4);
TASK_PP(16'hA969,4);
TASK_PP(16'hA96A,4);
TASK_PP(16'hA96B,4);
TASK_PP(16'hA96C,4);
TASK_PP(16'hA96D,4);
TASK_PP(16'hA96E,4);
TASK_PP(16'hA96F,4);
TASK_PP(16'hA970,4);
TASK_PP(16'hA971,4);
TASK_PP(16'hA972,4);
TASK_PP(16'hA973,4);
TASK_PP(16'hA974,4);
TASK_PP(16'hA975,4);
TASK_PP(16'hA976,4);
TASK_PP(16'hA977,4);
TASK_PP(16'hA978,4);
TASK_PP(16'hA979,4);
TASK_PP(16'hA97A,4);
TASK_PP(16'hA97B,4);
TASK_PP(16'hA97C,4);
TASK_PP(16'hA97D,4);
TASK_PP(16'hA97E,4);
TASK_PP(16'hA97F,4);
TASK_PP(16'hA980,4);
TASK_PP(16'hA981,4);
TASK_PP(16'hA982,4);
TASK_PP(16'hA983,4);
TASK_PP(16'hA984,4);
TASK_PP(16'hA985,4);
TASK_PP(16'hA986,4);
TASK_PP(16'hA987,4);
TASK_PP(16'hA988,4);
TASK_PP(16'hA989,4);
TASK_PP(16'hA98A,4);
TASK_PP(16'hA98B,4);
TASK_PP(16'hA98C,4);
TASK_PP(16'hA98D,4);
TASK_PP(16'hA98E,4);
TASK_PP(16'hA98F,4);
TASK_PP(16'hA990,4);
TASK_PP(16'hA991,4);
TASK_PP(16'hA992,4);
TASK_PP(16'hA993,4);
TASK_PP(16'hA994,4);
TASK_PP(16'hA995,4);
TASK_PP(16'hA996,4);
TASK_PP(16'hA997,4);
TASK_PP(16'hA998,4);
TASK_PP(16'hA999,4);
TASK_PP(16'hA99A,4);
TASK_PP(16'hA99B,4);
TASK_PP(16'hA99C,4);
TASK_PP(16'hA99D,4);
TASK_PP(16'hA99E,4);
TASK_PP(16'hA99F,4);
TASK_PP(16'hA9A0,4);
TASK_PP(16'hA9A1,4);
TASK_PP(16'hA9A2,4);
TASK_PP(16'hA9A3,4);
TASK_PP(16'hA9A4,4);
TASK_PP(16'hA9A5,4);
TASK_PP(16'hA9A6,4);
TASK_PP(16'hA9A7,4);
TASK_PP(16'hA9A8,4);
TASK_PP(16'hA9A9,4);
TASK_PP(16'hA9AA,4);
TASK_PP(16'hA9AB,4);
TASK_PP(16'hA9AC,4);
TASK_PP(16'hA9AD,4);
TASK_PP(16'hA9AE,4);
TASK_PP(16'hA9AF,4);
TASK_PP(16'hA9B0,4);
TASK_PP(16'hA9B1,4);
TASK_PP(16'hA9B2,4);
TASK_PP(16'hA9B3,4);
TASK_PP(16'hA9B4,4);
TASK_PP(16'hA9B5,4);
TASK_PP(16'hA9B6,4);
TASK_PP(16'hA9B7,4);
TASK_PP(16'hA9B8,4);
TASK_PP(16'hA9B9,4);
TASK_PP(16'hA9BA,4);
TASK_PP(16'hA9BB,4);
TASK_PP(16'hA9BC,4);
TASK_PP(16'hA9BD,4);
TASK_PP(16'hA9BE,4);
TASK_PP(16'hA9BF,4);
TASK_PP(16'hA9C0,4);
TASK_PP(16'hA9C1,4);
TASK_PP(16'hA9C2,4);
TASK_PP(16'hA9C3,4);
TASK_PP(16'hA9C4,4);
TASK_PP(16'hA9C5,4);
TASK_PP(16'hA9C6,4);
TASK_PP(16'hA9C7,4);
TASK_PP(16'hA9C8,4);
TASK_PP(16'hA9C9,4);
TASK_PP(16'hA9CA,4);
TASK_PP(16'hA9CB,4);
TASK_PP(16'hA9CC,4);
TASK_PP(16'hA9CD,4);
TASK_PP(16'hA9CE,4);
TASK_PP(16'hA9CF,4);
TASK_PP(16'hA9D0,4);
TASK_PP(16'hA9D1,4);
TASK_PP(16'hA9D2,4);
TASK_PP(16'hA9D3,4);
TASK_PP(16'hA9D4,4);
TASK_PP(16'hA9D5,4);
TASK_PP(16'hA9D6,4);
TASK_PP(16'hA9D7,4);
TASK_PP(16'hA9D8,4);
TASK_PP(16'hA9D9,4);
TASK_PP(16'hA9DA,4);
TASK_PP(16'hA9DB,4);
TASK_PP(16'hA9DC,4);
TASK_PP(16'hA9DD,4);
TASK_PP(16'hA9DE,4);
TASK_PP(16'hA9DF,4);
TASK_PP(16'hA9E0,4);
TASK_PP(16'hA9E1,4);
TASK_PP(16'hA9E2,4);
TASK_PP(16'hA9E3,4);
TASK_PP(16'hA9E4,4);
TASK_PP(16'hA9E5,4);
TASK_PP(16'hA9E6,4);
TASK_PP(16'hA9E7,4);
TASK_PP(16'hA9E8,4);
TASK_PP(16'hA9E9,4);
TASK_PP(16'hA9EA,4);
TASK_PP(16'hA9EB,4);
TASK_PP(16'hA9EC,4);
TASK_PP(16'hA9ED,4);
TASK_PP(16'hA9EE,4);
TASK_PP(16'hA9EF,4);
TASK_PP(16'hA9F0,4);
TASK_PP(16'hA9F1,4);
TASK_PP(16'hA9F2,4);
TASK_PP(16'hA9F3,4);
TASK_PP(16'hA9F4,4);
TASK_PP(16'hA9F5,4);
TASK_PP(16'hA9F6,4);
TASK_PP(16'hA9F7,4);
TASK_PP(16'hA9F8,4);
TASK_PP(16'hA9F9,4);
TASK_PP(16'hA9FA,4);
TASK_PP(16'hA9FB,4);
TASK_PP(16'hA9FC,4);
TASK_PP(16'hA9FD,4);
TASK_PP(16'hA9FE,4);
TASK_PP(16'hA9FF,4);
TASK_PP(16'hAA00,4);
TASK_PP(16'hAA01,4);
TASK_PP(16'hAA02,4);
TASK_PP(16'hAA03,4);
TASK_PP(16'hAA04,4);
TASK_PP(16'hAA05,4);
TASK_PP(16'hAA06,4);
TASK_PP(16'hAA07,4);
TASK_PP(16'hAA08,4);
TASK_PP(16'hAA09,4);
TASK_PP(16'hAA0A,4);
TASK_PP(16'hAA0B,4);
TASK_PP(16'hAA0C,4);
TASK_PP(16'hAA0D,4);
TASK_PP(16'hAA0E,4);
TASK_PP(16'hAA0F,4);
TASK_PP(16'hAA10,4);
TASK_PP(16'hAA11,4);
TASK_PP(16'hAA12,4);
TASK_PP(16'hAA13,4);
TASK_PP(16'hAA14,4);
TASK_PP(16'hAA15,4);
TASK_PP(16'hAA16,4);
TASK_PP(16'hAA17,4);
TASK_PP(16'hAA18,4);
TASK_PP(16'hAA19,4);
TASK_PP(16'hAA1A,4);
TASK_PP(16'hAA1B,4);
TASK_PP(16'hAA1C,4);
TASK_PP(16'hAA1D,4);
TASK_PP(16'hAA1E,4);
TASK_PP(16'hAA1F,4);
TASK_PP(16'hAA20,4);
TASK_PP(16'hAA21,4);
TASK_PP(16'hAA22,4);
TASK_PP(16'hAA23,4);
TASK_PP(16'hAA24,4);
TASK_PP(16'hAA25,4);
TASK_PP(16'hAA26,4);
TASK_PP(16'hAA27,4);
TASK_PP(16'hAA28,4);
TASK_PP(16'hAA29,4);
TASK_PP(16'hAA2A,4);
TASK_PP(16'hAA2B,4);
TASK_PP(16'hAA2C,4);
TASK_PP(16'hAA2D,4);
TASK_PP(16'hAA2E,4);
TASK_PP(16'hAA2F,4);
TASK_PP(16'hAA30,4);
TASK_PP(16'hAA31,4);
TASK_PP(16'hAA32,4);
TASK_PP(16'hAA33,4);
TASK_PP(16'hAA34,4);
TASK_PP(16'hAA35,4);
TASK_PP(16'hAA36,4);
TASK_PP(16'hAA37,4);
TASK_PP(16'hAA38,4);
TASK_PP(16'hAA39,4);
TASK_PP(16'hAA3A,4);
TASK_PP(16'hAA3B,4);
TASK_PP(16'hAA3C,4);
TASK_PP(16'hAA3D,4);
TASK_PP(16'hAA3E,4);
TASK_PP(16'hAA3F,4);
TASK_PP(16'hAA40,4);
TASK_PP(16'hAA41,4);
TASK_PP(16'hAA42,4);
TASK_PP(16'hAA43,4);
TASK_PP(16'hAA44,4);
TASK_PP(16'hAA45,4);
TASK_PP(16'hAA46,4);
TASK_PP(16'hAA47,4);
TASK_PP(16'hAA48,4);
TASK_PP(16'hAA49,4);
TASK_PP(16'hAA4A,4);
TASK_PP(16'hAA4B,4);
TASK_PP(16'hAA4C,4);
TASK_PP(16'hAA4D,4);
TASK_PP(16'hAA4E,4);
TASK_PP(16'hAA4F,4);
TASK_PP(16'hAA50,4);
TASK_PP(16'hAA51,4);
TASK_PP(16'hAA52,4);
TASK_PP(16'hAA53,4);
TASK_PP(16'hAA54,4);
TASK_PP(16'hAA55,4);
TASK_PP(16'hAA56,4);
TASK_PP(16'hAA57,4);
TASK_PP(16'hAA58,4);
TASK_PP(16'hAA59,4);
TASK_PP(16'hAA5A,4);
TASK_PP(16'hAA5B,4);
TASK_PP(16'hAA5C,4);
TASK_PP(16'hAA5D,4);
TASK_PP(16'hAA5E,4);
TASK_PP(16'hAA5F,4);
TASK_PP(16'hAA60,4);
TASK_PP(16'hAA61,4);
TASK_PP(16'hAA62,4);
TASK_PP(16'hAA63,4);
TASK_PP(16'hAA64,4);
TASK_PP(16'hAA65,4);
TASK_PP(16'hAA66,4);
TASK_PP(16'hAA67,4);
TASK_PP(16'hAA68,4);
TASK_PP(16'hAA69,4);
TASK_PP(16'hAA6A,4);
TASK_PP(16'hAA6B,4);
TASK_PP(16'hAA6C,4);
TASK_PP(16'hAA6D,4);
TASK_PP(16'hAA6E,4);
TASK_PP(16'hAA6F,4);
TASK_PP(16'hAA70,4);
TASK_PP(16'hAA71,4);
TASK_PP(16'hAA72,4);
TASK_PP(16'hAA73,4);
TASK_PP(16'hAA74,4);
TASK_PP(16'hAA75,4);
TASK_PP(16'hAA76,4);
TASK_PP(16'hAA77,4);
TASK_PP(16'hAA78,4);
TASK_PP(16'hAA79,4);
TASK_PP(16'hAA7A,4);
TASK_PP(16'hAA7B,4);
TASK_PP(16'hAA7C,4);
TASK_PP(16'hAA7D,4);
TASK_PP(16'hAA7E,4);
TASK_PP(16'hAA7F,4);
TASK_PP(16'hAA80,4);
TASK_PP(16'hAA81,4);
TASK_PP(16'hAA82,4);
TASK_PP(16'hAA83,4);
TASK_PP(16'hAA84,4);
TASK_PP(16'hAA85,4);
TASK_PP(16'hAA86,4);
TASK_PP(16'hAA87,4);
TASK_PP(16'hAA88,4);
TASK_PP(16'hAA89,4);
TASK_PP(16'hAA8A,4);
TASK_PP(16'hAA8B,4);
TASK_PP(16'hAA8C,4);
TASK_PP(16'hAA8D,4);
TASK_PP(16'hAA8E,4);
TASK_PP(16'hAA8F,4);
TASK_PP(16'hAA90,4);
TASK_PP(16'hAA91,4);
TASK_PP(16'hAA92,4);
TASK_PP(16'hAA93,4);
TASK_PP(16'hAA94,4);
TASK_PP(16'hAA95,4);
TASK_PP(16'hAA96,4);
TASK_PP(16'hAA97,4);
TASK_PP(16'hAA98,4);
TASK_PP(16'hAA99,4);
TASK_PP(16'hAA9A,4);
TASK_PP(16'hAA9B,4);
TASK_PP(16'hAA9C,4);
TASK_PP(16'hAA9D,4);
TASK_PP(16'hAA9E,4);
TASK_PP(16'hAA9F,4);
TASK_PP(16'hAAA0,4);
TASK_PP(16'hAAA1,4);
TASK_PP(16'hAAA2,4);
TASK_PP(16'hAAA3,4);
TASK_PP(16'hAAA4,4);
TASK_PP(16'hAAA5,4);
TASK_PP(16'hAAA6,4);
TASK_PP(16'hAAA7,4);
TASK_PP(16'hAAA8,4);
TASK_PP(16'hAAA9,4);
TASK_PP(16'hAAAA,4);
TASK_PP(16'hAAAB,4);
TASK_PP(16'hAAAC,4);
TASK_PP(16'hAAAD,4);
TASK_PP(16'hAAAE,4);
TASK_PP(16'hAAAF,4);
TASK_PP(16'hAAB0,4);
TASK_PP(16'hAAB1,4);
TASK_PP(16'hAAB2,4);
TASK_PP(16'hAAB3,4);
TASK_PP(16'hAAB4,4);
TASK_PP(16'hAAB5,4);
TASK_PP(16'hAAB6,4);
TASK_PP(16'hAAB7,4);
TASK_PP(16'hAAB8,4);
TASK_PP(16'hAAB9,4);
TASK_PP(16'hAABA,4);
TASK_PP(16'hAABB,4);
TASK_PP(16'hAABC,4);
TASK_PP(16'hAABD,4);
TASK_PP(16'hAABE,4);
TASK_PP(16'hAABF,4);
TASK_PP(16'hAAC0,4);
TASK_PP(16'hAAC1,4);
TASK_PP(16'hAAC2,4);
TASK_PP(16'hAAC3,4);
TASK_PP(16'hAAC4,4);
TASK_PP(16'hAAC5,4);
TASK_PP(16'hAAC6,4);
TASK_PP(16'hAAC7,4);
TASK_PP(16'hAAC8,4);
TASK_PP(16'hAAC9,4);
TASK_PP(16'hAACA,4);
TASK_PP(16'hAACB,4);
TASK_PP(16'hAACC,4);
TASK_PP(16'hAACD,4);
TASK_PP(16'hAACE,4);
TASK_PP(16'hAACF,4);
TASK_PP(16'hAAD0,4);
TASK_PP(16'hAAD1,4);
TASK_PP(16'hAAD2,4);
TASK_PP(16'hAAD3,4);
TASK_PP(16'hAAD4,4);
TASK_PP(16'hAAD5,4);
TASK_PP(16'hAAD6,4);
TASK_PP(16'hAAD7,4);
TASK_PP(16'hAAD8,4);
TASK_PP(16'hAAD9,4);
TASK_PP(16'hAADA,4);
TASK_PP(16'hAADB,4);
TASK_PP(16'hAADC,4);
TASK_PP(16'hAADD,4);
TASK_PP(16'hAADE,4);
TASK_PP(16'hAADF,4);
TASK_PP(16'hAAE0,4);
TASK_PP(16'hAAE1,4);
TASK_PP(16'hAAE2,4);
TASK_PP(16'hAAE3,4);
TASK_PP(16'hAAE4,4);
TASK_PP(16'hAAE5,4);
TASK_PP(16'hAAE6,4);
TASK_PP(16'hAAE7,4);
TASK_PP(16'hAAE8,4);
TASK_PP(16'hAAE9,4);
TASK_PP(16'hAAEA,4);
TASK_PP(16'hAAEB,4);
TASK_PP(16'hAAEC,4);
TASK_PP(16'hAAED,4);
TASK_PP(16'hAAEE,4);
TASK_PP(16'hAAEF,4);
TASK_PP(16'hAAF0,4);
TASK_PP(16'hAAF1,4);
TASK_PP(16'hAAF2,4);
TASK_PP(16'hAAF3,4);
TASK_PP(16'hAAF4,4);
TASK_PP(16'hAAF5,4);
TASK_PP(16'hAAF6,4);
TASK_PP(16'hAAF7,4);
TASK_PP(16'hAAF8,4);
TASK_PP(16'hAAF9,4);
TASK_PP(16'hAAFA,4);
TASK_PP(16'hAAFB,4);
TASK_PP(16'hAAFC,4);
TASK_PP(16'hAAFD,4);
TASK_PP(16'hAAFE,4);
TASK_PP(16'hAAFF,4);
TASK_PP(16'hAB00,4);
TASK_PP(16'hAB01,4);
TASK_PP(16'hAB02,4);
TASK_PP(16'hAB03,4);
TASK_PP(16'hAB04,4);
TASK_PP(16'hAB05,4);
TASK_PP(16'hAB06,4);
TASK_PP(16'hAB07,4);
TASK_PP(16'hAB08,4);
TASK_PP(16'hAB09,4);
TASK_PP(16'hAB0A,4);
TASK_PP(16'hAB0B,4);
TASK_PP(16'hAB0C,4);
TASK_PP(16'hAB0D,4);
TASK_PP(16'hAB0E,4);
TASK_PP(16'hAB0F,4);
TASK_PP(16'hAB10,4);
TASK_PP(16'hAB11,4);
TASK_PP(16'hAB12,4);
TASK_PP(16'hAB13,4);
TASK_PP(16'hAB14,4);
TASK_PP(16'hAB15,4);
TASK_PP(16'hAB16,4);
TASK_PP(16'hAB17,4);
TASK_PP(16'hAB18,4);
TASK_PP(16'hAB19,4);
TASK_PP(16'hAB1A,4);
TASK_PP(16'hAB1B,4);
TASK_PP(16'hAB1C,4);
TASK_PP(16'hAB1D,4);
TASK_PP(16'hAB1E,4);
TASK_PP(16'hAB1F,4);
TASK_PP(16'hAB20,4);
TASK_PP(16'hAB21,4);
TASK_PP(16'hAB22,4);
TASK_PP(16'hAB23,4);
TASK_PP(16'hAB24,4);
TASK_PP(16'hAB25,4);
TASK_PP(16'hAB26,4);
TASK_PP(16'hAB27,4);
TASK_PP(16'hAB28,4);
TASK_PP(16'hAB29,4);
TASK_PP(16'hAB2A,4);
TASK_PP(16'hAB2B,4);
TASK_PP(16'hAB2C,4);
TASK_PP(16'hAB2D,4);
TASK_PP(16'hAB2E,4);
TASK_PP(16'hAB2F,4);
TASK_PP(16'hAB30,4);
TASK_PP(16'hAB31,4);
TASK_PP(16'hAB32,4);
TASK_PP(16'hAB33,4);
TASK_PP(16'hAB34,4);
TASK_PP(16'hAB35,4);
TASK_PP(16'hAB36,4);
TASK_PP(16'hAB37,4);
TASK_PP(16'hAB38,4);
TASK_PP(16'hAB39,4);
TASK_PP(16'hAB3A,4);
TASK_PP(16'hAB3B,4);
TASK_PP(16'hAB3C,4);
TASK_PP(16'hAB3D,4);
TASK_PP(16'hAB3E,4);
TASK_PP(16'hAB3F,4);
TASK_PP(16'hAB40,4);
TASK_PP(16'hAB41,4);
TASK_PP(16'hAB42,4);
TASK_PP(16'hAB43,4);
TASK_PP(16'hAB44,4);
TASK_PP(16'hAB45,4);
TASK_PP(16'hAB46,4);
TASK_PP(16'hAB47,4);
TASK_PP(16'hAB48,4);
TASK_PP(16'hAB49,4);
TASK_PP(16'hAB4A,4);
TASK_PP(16'hAB4B,4);
TASK_PP(16'hAB4C,4);
TASK_PP(16'hAB4D,4);
TASK_PP(16'hAB4E,4);
TASK_PP(16'hAB4F,4);
TASK_PP(16'hAB50,4);
TASK_PP(16'hAB51,4);
TASK_PP(16'hAB52,4);
TASK_PP(16'hAB53,4);
TASK_PP(16'hAB54,4);
TASK_PP(16'hAB55,4);
TASK_PP(16'hAB56,4);
TASK_PP(16'hAB57,4);
TASK_PP(16'hAB58,4);
TASK_PP(16'hAB59,4);
TASK_PP(16'hAB5A,4);
TASK_PP(16'hAB5B,4);
TASK_PP(16'hAB5C,4);
TASK_PP(16'hAB5D,4);
TASK_PP(16'hAB5E,4);
TASK_PP(16'hAB5F,4);
TASK_PP(16'hAB60,4);
TASK_PP(16'hAB61,4);
TASK_PP(16'hAB62,4);
TASK_PP(16'hAB63,4);
TASK_PP(16'hAB64,4);
TASK_PP(16'hAB65,4);
TASK_PP(16'hAB66,4);
TASK_PP(16'hAB67,4);
TASK_PP(16'hAB68,4);
TASK_PP(16'hAB69,4);
TASK_PP(16'hAB6A,4);
TASK_PP(16'hAB6B,4);
TASK_PP(16'hAB6C,4);
TASK_PP(16'hAB6D,4);
TASK_PP(16'hAB6E,4);
TASK_PP(16'hAB6F,4);
TASK_PP(16'hAB70,4);
TASK_PP(16'hAB71,4);
TASK_PP(16'hAB72,4);
TASK_PP(16'hAB73,4);
TASK_PP(16'hAB74,4);
TASK_PP(16'hAB75,4);
TASK_PP(16'hAB76,4);
TASK_PP(16'hAB77,4);
TASK_PP(16'hAB78,4);
TASK_PP(16'hAB79,4);
TASK_PP(16'hAB7A,4);
TASK_PP(16'hAB7B,4);
TASK_PP(16'hAB7C,4);
TASK_PP(16'hAB7D,4);
TASK_PP(16'hAB7E,4);
TASK_PP(16'hAB7F,4);
TASK_PP(16'hAB80,4);
TASK_PP(16'hAB81,4);
TASK_PP(16'hAB82,4);
TASK_PP(16'hAB83,4);
TASK_PP(16'hAB84,4);
TASK_PP(16'hAB85,4);
TASK_PP(16'hAB86,4);
TASK_PP(16'hAB87,4);
TASK_PP(16'hAB88,4);
TASK_PP(16'hAB89,4);
TASK_PP(16'hAB8A,4);
TASK_PP(16'hAB8B,4);
TASK_PP(16'hAB8C,4);
TASK_PP(16'hAB8D,4);
TASK_PP(16'hAB8E,4);
TASK_PP(16'hAB8F,4);
TASK_PP(16'hAB90,4);
TASK_PP(16'hAB91,4);
TASK_PP(16'hAB92,4);
TASK_PP(16'hAB93,4);
TASK_PP(16'hAB94,4);
TASK_PP(16'hAB95,4);
TASK_PP(16'hAB96,4);
TASK_PP(16'hAB97,4);
TASK_PP(16'hAB98,4);
TASK_PP(16'hAB99,4);
TASK_PP(16'hAB9A,4);
TASK_PP(16'hAB9B,4);
TASK_PP(16'hAB9C,4);
TASK_PP(16'hAB9D,4);
TASK_PP(16'hAB9E,4);
TASK_PP(16'hAB9F,4);
TASK_PP(16'hABA0,4);
TASK_PP(16'hABA1,4);
TASK_PP(16'hABA2,4);
TASK_PP(16'hABA3,4);
TASK_PP(16'hABA4,4);
TASK_PP(16'hABA5,4);
TASK_PP(16'hABA6,4);
TASK_PP(16'hABA7,4);
TASK_PP(16'hABA8,4);
TASK_PP(16'hABA9,4);
TASK_PP(16'hABAA,4);
TASK_PP(16'hABAB,4);
TASK_PP(16'hABAC,4);
TASK_PP(16'hABAD,4);
TASK_PP(16'hABAE,4);
TASK_PP(16'hABAF,4);
TASK_PP(16'hABB0,4);
TASK_PP(16'hABB1,4);
TASK_PP(16'hABB2,4);
TASK_PP(16'hABB3,4);
TASK_PP(16'hABB4,4);
TASK_PP(16'hABB5,4);
TASK_PP(16'hABB6,4);
TASK_PP(16'hABB7,4);
TASK_PP(16'hABB8,4);
TASK_PP(16'hABB9,4);
TASK_PP(16'hABBA,4);
TASK_PP(16'hABBB,4);
TASK_PP(16'hABBC,4);
TASK_PP(16'hABBD,4);
TASK_PP(16'hABBE,4);
TASK_PP(16'hABBF,4);
TASK_PP(16'hABC0,4);
TASK_PP(16'hABC1,4);
TASK_PP(16'hABC2,4);
TASK_PP(16'hABC3,4);
TASK_PP(16'hABC4,4);
TASK_PP(16'hABC5,4);
TASK_PP(16'hABC6,4);
TASK_PP(16'hABC7,4);
TASK_PP(16'hABC8,4);
TASK_PP(16'hABC9,4);
TASK_PP(16'hABCA,4);
TASK_PP(16'hABCB,4);
TASK_PP(16'hABCC,4);
TASK_PP(16'hABCD,4);
TASK_PP(16'hABCE,4);
TASK_PP(16'hABCF,4);
TASK_PP(16'hABD0,4);
TASK_PP(16'hABD1,4);
TASK_PP(16'hABD2,4);
TASK_PP(16'hABD3,4);
TASK_PP(16'hABD4,4);
TASK_PP(16'hABD5,4);
TASK_PP(16'hABD6,4);
TASK_PP(16'hABD7,4);
TASK_PP(16'hABD8,4);
TASK_PP(16'hABD9,4);
TASK_PP(16'hABDA,4);
TASK_PP(16'hABDB,4);
TASK_PP(16'hABDC,4);
TASK_PP(16'hABDD,4);
TASK_PP(16'hABDE,4);
TASK_PP(16'hABDF,4);
TASK_PP(16'hABE0,4);
TASK_PP(16'hABE1,4);
TASK_PP(16'hABE2,4);
TASK_PP(16'hABE3,4);
TASK_PP(16'hABE4,4);
TASK_PP(16'hABE5,4);
TASK_PP(16'hABE6,4);
TASK_PP(16'hABE7,4);
TASK_PP(16'hABE8,4);
TASK_PP(16'hABE9,4);
TASK_PP(16'hABEA,4);
TASK_PP(16'hABEB,4);
TASK_PP(16'hABEC,4);
TASK_PP(16'hABED,4);
TASK_PP(16'hABEE,4);
TASK_PP(16'hABEF,4);
TASK_PP(16'hABF0,4);
TASK_PP(16'hABF1,4);
TASK_PP(16'hABF2,4);
TASK_PP(16'hABF3,4);
TASK_PP(16'hABF4,4);
TASK_PP(16'hABF5,4);
TASK_PP(16'hABF6,4);
TASK_PP(16'hABF7,4);
TASK_PP(16'hABF8,4);
TASK_PP(16'hABF9,4);
TASK_PP(16'hABFA,4);
TASK_PP(16'hABFB,4);
TASK_PP(16'hABFC,4);
TASK_PP(16'hABFD,4);
TASK_PP(16'hABFE,4);
TASK_PP(16'hABFF,4);
TASK_PP(16'hAC00,4);
TASK_PP(16'hAC01,4);
TASK_PP(16'hAC02,4);
TASK_PP(16'hAC03,4);
TASK_PP(16'hAC04,4);
TASK_PP(16'hAC05,4);
TASK_PP(16'hAC06,4);
TASK_PP(16'hAC07,4);
TASK_PP(16'hAC08,4);
TASK_PP(16'hAC09,4);
TASK_PP(16'hAC0A,4);
TASK_PP(16'hAC0B,4);
TASK_PP(16'hAC0C,4);
TASK_PP(16'hAC0D,4);
TASK_PP(16'hAC0E,4);
TASK_PP(16'hAC0F,4);
TASK_PP(16'hAC10,4);
TASK_PP(16'hAC11,4);
TASK_PP(16'hAC12,4);
TASK_PP(16'hAC13,4);
TASK_PP(16'hAC14,4);
TASK_PP(16'hAC15,4);
TASK_PP(16'hAC16,4);
TASK_PP(16'hAC17,4);
TASK_PP(16'hAC18,4);
TASK_PP(16'hAC19,4);
TASK_PP(16'hAC1A,4);
TASK_PP(16'hAC1B,4);
TASK_PP(16'hAC1C,4);
TASK_PP(16'hAC1D,4);
TASK_PP(16'hAC1E,4);
TASK_PP(16'hAC1F,4);
TASK_PP(16'hAC20,4);
TASK_PP(16'hAC21,4);
TASK_PP(16'hAC22,4);
TASK_PP(16'hAC23,4);
TASK_PP(16'hAC24,4);
TASK_PP(16'hAC25,4);
TASK_PP(16'hAC26,4);
TASK_PP(16'hAC27,4);
TASK_PP(16'hAC28,4);
TASK_PP(16'hAC29,4);
TASK_PP(16'hAC2A,4);
TASK_PP(16'hAC2B,4);
TASK_PP(16'hAC2C,4);
TASK_PP(16'hAC2D,4);
TASK_PP(16'hAC2E,4);
TASK_PP(16'hAC2F,4);
TASK_PP(16'hAC30,4);
TASK_PP(16'hAC31,4);
TASK_PP(16'hAC32,4);
TASK_PP(16'hAC33,4);
TASK_PP(16'hAC34,4);
TASK_PP(16'hAC35,4);
TASK_PP(16'hAC36,4);
TASK_PP(16'hAC37,4);
TASK_PP(16'hAC38,4);
TASK_PP(16'hAC39,4);
TASK_PP(16'hAC3A,4);
TASK_PP(16'hAC3B,4);
TASK_PP(16'hAC3C,4);
TASK_PP(16'hAC3D,4);
TASK_PP(16'hAC3E,4);
TASK_PP(16'hAC3F,4);
TASK_PP(16'hAC40,4);
TASK_PP(16'hAC41,4);
TASK_PP(16'hAC42,4);
TASK_PP(16'hAC43,4);
TASK_PP(16'hAC44,4);
TASK_PP(16'hAC45,4);
TASK_PP(16'hAC46,4);
TASK_PP(16'hAC47,4);
TASK_PP(16'hAC48,4);
TASK_PP(16'hAC49,4);
TASK_PP(16'hAC4A,4);
TASK_PP(16'hAC4B,4);
TASK_PP(16'hAC4C,4);
TASK_PP(16'hAC4D,4);
TASK_PP(16'hAC4E,4);
TASK_PP(16'hAC4F,4);
TASK_PP(16'hAC50,4);
TASK_PP(16'hAC51,4);
TASK_PP(16'hAC52,4);
TASK_PP(16'hAC53,4);
TASK_PP(16'hAC54,4);
TASK_PP(16'hAC55,4);
TASK_PP(16'hAC56,4);
TASK_PP(16'hAC57,4);
TASK_PP(16'hAC58,4);
TASK_PP(16'hAC59,4);
TASK_PP(16'hAC5A,4);
TASK_PP(16'hAC5B,4);
TASK_PP(16'hAC5C,4);
TASK_PP(16'hAC5D,4);
TASK_PP(16'hAC5E,4);
TASK_PP(16'hAC5F,4);
TASK_PP(16'hAC60,4);
TASK_PP(16'hAC61,4);
TASK_PP(16'hAC62,4);
TASK_PP(16'hAC63,4);
TASK_PP(16'hAC64,4);
TASK_PP(16'hAC65,4);
TASK_PP(16'hAC66,4);
TASK_PP(16'hAC67,4);
TASK_PP(16'hAC68,4);
TASK_PP(16'hAC69,4);
TASK_PP(16'hAC6A,4);
TASK_PP(16'hAC6B,4);
TASK_PP(16'hAC6C,4);
TASK_PP(16'hAC6D,4);
TASK_PP(16'hAC6E,4);
TASK_PP(16'hAC6F,4);
TASK_PP(16'hAC70,4);
TASK_PP(16'hAC71,4);
TASK_PP(16'hAC72,4);
TASK_PP(16'hAC73,4);
TASK_PP(16'hAC74,4);
TASK_PP(16'hAC75,4);
TASK_PP(16'hAC76,4);
TASK_PP(16'hAC77,4);
TASK_PP(16'hAC78,4);
TASK_PP(16'hAC79,4);
TASK_PP(16'hAC7A,4);
TASK_PP(16'hAC7B,4);
TASK_PP(16'hAC7C,4);
TASK_PP(16'hAC7D,4);
TASK_PP(16'hAC7E,4);
TASK_PP(16'hAC7F,4);
TASK_PP(16'hAC80,4);
TASK_PP(16'hAC81,4);
TASK_PP(16'hAC82,4);
TASK_PP(16'hAC83,4);
TASK_PP(16'hAC84,4);
TASK_PP(16'hAC85,4);
TASK_PP(16'hAC86,4);
TASK_PP(16'hAC87,4);
TASK_PP(16'hAC88,4);
TASK_PP(16'hAC89,4);
TASK_PP(16'hAC8A,4);
TASK_PP(16'hAC8B,4);
TASK_PP(16'hAC8C,4);
TASK_PP(16'hAC8D,4);
TASK_PP(16'hAC8E,4);
TASK_PP(16'hAC8F,4);
TASK_PP(16'hAC90,4);
TASK_PP(16'hAC91,4);
TASK_PP(16'hAC92,4);
TASK_PP(16'hAC93,4);
TASK_PP(16'hAC94,4);
TASK_PP(16'hAC95,4);
TASK_PP(16'hAC96,4);
TASK_PP(16'hAC97,4);
TASK_PP(16'hAC98,4);
TASK_PP(16'hAC99,4);
TASK_PP(16'hAC9A,4);
TASK_PP(16'hAC9B,4);
TASK_PP(16'hAC9C,4);
TASK_PP(16'hAC9D,4);
TASK_PP(16'hAC9E,4);
TASK_PP(16'hAC9F,4);
TASK_PP(16'hACA0,4);
TASK_PP(16'hACA1,4);
TASK_PP(16'hACA2,4);
TASK_PP(16'hACA3,4);
TASK_PP(16'hACA4,4);
TASK_PP(16'hACA5,4);
TASK_PP(16'hACA6,4);
TASK_PP(16'hACA7,4);
TASK_PP(16'hACA8,4);
TASK_PP(16'hACA9,4);
TASK_PP(16'hACAA,4);
TASK_PP(16'hACAB,4);
TASK_PP(16'hACAC,4);
TASK_PP(16'hACAD,4);
TASK_PP(16'hACAE,4);
TASK_PP(16'hACAF,4);
TASK_PP(16'hACB0,4);
TASK_PP(16'hACB1,4);
TASK_PP(16'hACB2,4);
TASK_PP(16'hACB3,4);
TASK_PP(16'hACB4,4);
TASK_PP(16'hACB5,4);
TASK_PP(16'hACB6,4);
TASK_PP(16'hACB7,4);
TASK_PP(16'hACB8,4);
TASK_PP(16'hACB9,4);
TASK_PP(16'hACBA,4);
TASK_PP(16'hACBB,4);
TASK_PP(16'hACBC,4);
TASK_PP(16'hACBD,4);
TASK_PP(16'hACBE,4);
TASK_PP(16'hACBF,4);
TASK_PP(16'hACC0,4);
TASK_PP(16'hACC1,4);
TASK_PP(16'hACC2,4);
TASK_PP(16'hACC3,4);
TASK_PP(16'hACC4,4);
TASK_PP(16'hACC5,4);
TASK_PP(16'hACC6,4);
TASK_PP(16'hACC7,4);
TASK_PP(16'hACC8,4);
TASK_PP(16'hACC9,4);
TASK_PP(16'hACCA,4);
TASK_PP(16'hACCB,4);
TASK_PP(16'hACCC,4);
TASK_PP(16'hACCD,4);
TASK_PP(16'hACCE,4);
TASK_PP(16'hACCF,4);
TASK_PP(16'hACD0,4);
TASK_PP(16'hACD1,4);
TASK_PP(16'hACD2,4);
TASK_PP(16'hACD3,4);
TASK_PP(16'hACD4,4);
TASK_PP(16'hACD5,4);
TASK_PP(16'hACD6,4);
TASK_PP(16'hACD7,4);
TASK_PP(16'hACD8,4);
TASK_PP(16'hACD9,4);
TASK_PP(16'hACDA,4);
TASK_PP(16'hACDB,4);
TASK_PP(16'hACDC,4);
TASK_PP(16'hACDD,4);
TASK_PP(16'hACDE,4);
TASK_PP(16'hACDF,4);
TASK_PP(16'hACE0,4);
TASK_PP(16'hACE1,4);
TASK_PP(16'hACE2,4);
TASK_PP(16'hACE3,4);
TASK_PP(16'hACE4,4);
TASK_PP(16'hACE5,4);
TASK_PP(16'hACE6,4);
TASK_PP(16'hACE7,4);
TASK_PP(16'hACE8,4);
TASK_PP(16'hACE9,4);
TASK_PP(16'hACEA,4);
TASK_PP(16'hACEB,4);
TASK_PP(16'hACEC,4);
TASK_PP(16'hACED,4);
TASK_PP(16'hACEE,4);
TASK_PP(16'hACEF,4);
TASK_PP(16'hACF0,4);
TASK_PP(16'hACF1,4);
TASK_PP(16'hACF2,4);
TASK_PP(16'hACF3,4);
TASK_PP(16'hACF4,4);
TASK_PP(16'hACF5,4);
TASK_PP(16'hACF6,4);
TASK_PP(16'hACF7,4);
TASK_PP(16'hACF8,4);
TASK_PP(16'hACF9,4);
TASK_PP(16'hACFA,4);
TASK_PP(16'hACFB,4);
TASK_PP(16'hACFC,4);
TASK_PP(16'hACFD,4);
TASK_PP(16'hACFE,4);
TASK_PP(16'hACFF,4);
TASK_PP(16'hAD00,4);
TASK_PP(16'hAD01,4);
TASK_PP(16'hAD02,4);
TASK_PP(16'hAD03,4);
TASK_PP(16'hAD04,4);
TASK_PP(16'hAD05,4);
TASK_PP(16'hAD06,4);
TASK_PP(16'hAD07,4);
TASK_PP(16'hAD08,4);
TASK_PP(16'hAD09,4);
TASK_PP(16'hAD0A,4);
TASK_PP(16'hAD0B,4);
TASK_PP(16'hAD0C,4);
TASK_PP(16'hAD0D,4);
TASK_PP(16'hAD0E,4);
TASK_PP(16'hAD0F,4);
TASK_PP(16'hAD10,4);
TASK_PP(16'hAD11,4);
TASK_PP(16'hAD12,4);
TASK_PP(16'hAD13,4);
TASK_PP(16'hAD14,4);
TASK_PP(16'hAD15,4);
TASK_PP(16'hAD16,4);
TASK_PP(16'hAD17,4);
TASK_PP(16'hAD18,4);
TASK_PP(16'hAD19,4);
TASK_PP(16'hAD1A,4);
TASK_PP(16'hAD1B,4);
TASK_PP(16'hAD1C,4);
TASK_PP(16'hAD1D,4);
TASK_PP(16'hAD1E,4);
TASK_PP(16'hAD1F,4);
TASK_PP(16'hAD20,4);
TASK_PP(16'hAD21,4);
TASK_PP(16'hAD22,4);
TASK_PP(16'hAD23,4);
TASK_PP(16'hAD24,4);
TASK_PP(16'hAD25,4);
TASK_PP(16'hAD26,4);
TASK_PP(16'hAD27,4);
TASK_PP(16'hAD28,4);
TASK_PP(16'hAD29,4);
TASK_PP(16'hAD2A,4);
TASK_PP(16'hAD2B,4);
TASK_PP(16'hAD2C,4);
TASK_PP(16'hAD2D,4);
TASK_PP(16'hAD2E,4);
TASK_PP(16'hAD2F,4);
TASK_PP(16'hAD30,4);
TASK_PP(16'hAD31,4);
TASK_PP(16'hAD32,4);
TASK_PP(16'hAD33,4);
TASK_PP(16'hAD34,4);
TASK_PP(16'hAD35,4);
TASK_PP(16'hAD36,4);
TASK_PP(16'hAD37,4);
TASK_PP(16'hAD38,4);
TASK_PP(16'hAD39,4);
TASK_PP(16'hAD3A,4);
TASK_PP(16'hAD3B,4);
TASK_PP(16'hAD3C,4);
TASK_PP(16'hAD3D,4);
TASK_PP(16'hAD3E,4);
TASK_PP(16'hAD3F,4);
TASK_PP(16'hAD40,4);
TASK_PP(16'hAD41,4);
TASK_PP(16'hAD42,4);
TASK_PP(16'hAD43,4);
TASK_PP(16'hAD44,4);
TASK_PP(16'hAD45,4);
TASK_PP(16'hAD46,4);
TASK_PP(16'hAD47,4);
TASK_PP(16'hAD48,4);
TASK_PP(16'hAD49,4);
TASK_PP(16'hAD4A,4);
TASK_PP(16'hAD4B,4);
TASK_PP(16'hAD4C,4);
TASK_PP(16'hAD4D,4);
TASK_PP(16'hAD4E,4);
TASK_PP(16'hAD4F,4);
TASK_PP(16'hAD50,4);
TASK_PP(16'hAD51,4);
TASK_PP(16'hAD52,4);
TASK_PP(16'hAD53,4);
TASK_PP(16'hAD54,4);
TASK_PP(16'hAD55,4);
TASK_PP(16'hAD56,4);
TASK_PP(16'hAD57,4);
TASK_PP(16'hAD58,4);
TASK_PP(16'hAD59,4);
TASK_PP(16'hAD5A,4);
TASK_PP(16'hAD5B,4);
TASK_PP(16'hAD5C,4);
TASK_PP(16'hAD5D,4);
TASK_PP(16'hAD5E,4);
TASK_PP(16'hAD5F,4);
TASK_PP(16'hAD60,4);
TASK_PP(16'hAD61,4);
TASK_PP(16'hAD62,4);
TASK_PP(16'hAD63,4);
TASK_PP(16'hAD64,4);
TASK_PP(16'hAD65,4);
TASK_PP(16'hAD66,4);
TASK_PP(16'hAD67,4);
TASK_PP(16'hAD68,4);
TASK_PP(16'hAD69,4);
TASK_PP(16'hAD6A,4);
TASK_PP(16'hAD6B,4);
TASK_PP(16'hAD6C,4);
TASK_PP(16'hAD6D,4);
TASK_PP(16'hAD6E,4);
TASK_PP(16'hAD6F,4);
TASK_PP(16'hAD70,4);
TASK_PP(16'hAD71,4);
TASK_PP(16'hAD72,4);
TASK_PP(16'hAD73,4);
TASK_PP(16'hAD74,4);
TASK_PP(16'hAD75,4);
TASK_PP(16'hAD76,4);
TASK_PP(16'hAD77,4);
TASK_PP(16'hAD78,4);
TASK_PP(16'hAD79,4);
TASK_PP(16'hAD7A,4);
TASK_PP(16'hAD7B,4);
TASK_PP(16'hAD7C,4);
TASK_PP(16'hAD7D,4);
TASK_PP(16'hAD7E,4);
TASK_PP(16'hAD7F,4);
TASK_PP(16'hAD80,4);
TASK_PP(16'hAD81,4);
TASK_PP(16'hAD82,4);
TASK_PP(16'hAD83,4);
TASK_PP(16'hAD84,4);
TASK_PP(16'hAD85,4);
TASK_PP(16'hAD86,4);
TASK_PP(16'hAD87,4);
TASK_PP(16'hAD88,4);
TASK_PP(16'hAD89,4);
TASK_PP(16'hAD8A,4);
TASK_PP(16'hAD8B,4);
TASK_PP(16'hAD8C,4);
TASK_PP(16'hAD8D,4);
TASK_PP(16'hAD8E,4);
TASK_PP(16'hAD8F,4);
TASK_PP(16'hAD90,4);
TASK_PP(16'hAD91,4);
TASK_PP(16'hAD92,4);
TASK_PP(16'hAD93,4);
TASK_PP(16'hAD94,4);
TASK_PP(16'hAD95,4);
TASK_PP(16'hAD96,4);
TASK_PP(16'hAD97,4);
TASK_PP(16'hAD98,4);
TASK_PP(16'hAD99,4);
TASK_PP(16'hAD9A,4);
TASK_PP(16'hAD9B,4);
TASK_PP(16'hAD9C,4);
TASK_PP(16'hAD9D,4);
TASK_PP(16'hAD9E,4);
TASK_PP(16'hAD9F,4);
TASK_PP(16'hADA0,4);
TASK_PP(16'hADA1,4);
TASK_PP(16'hADA2,4);
TASK_PP(16'hADA3,4);
TASK_PP(16'hADA4,4);
TASK_PP(16'hADA5,4);
TASK_PP(16'hADA6,4);
TASK_PP(16'hADA7,4);
TASK_PP(16'hADA8,4);
TASK_PP(16'hADA9,4);
TASK_PP(16'hADAA,4);
TASK_PP(16'hADAB,4);
TASK_PP(16'hADAC,4);
TASK_PP(16'hADAD,4);
TASK_PP(16'hADAE,4);
TASK_PP(16'hADAF,4);
TASK_PP(16'hADB0,4);
TASK_PP(16'hADB1,4);
TASK_PP(16'hADB2,4);
TASK_PP(16'hADB3,4);
TASK_PP(16'hADB4,4);
TASK_PP(16'hADB5,4);
TASK_PP(16'hADB6,4);
TASK_PP(16'hADB7,4);
TASK_PP(16'hADB8,4);
TASK_PP(16'hADB9,4);
TASK_PP(16'hADBA,4);
TASK_PP(16'hADBB,4);
TASK_PP(16'hADBC,4);
TASK_PP(16'hADBD,4);
TASK_PP(16'hADBE,4);
TASK_PP(16'hADBF,4);
TASK_PP(16'hADC0,4);
TASK_PP(16'hADC1,4);
TASK_PP(16'hADC2,4);
TASK_PP(16'hADC3,4);
TASK_PP(16'hADC4,4);
TASK_PP(16'hADC5,4);
TASK_PP(16'hADC6,4);
TASK_PP(16'hADC7,4);
TASK_PP(16'hADC8,4);
TASK_PP(16'hADC9,4);
TASK_PP(16'hADCA,4);
TASK_PP(16'hADCB,4);
TASK_PP(16'hADCC,4);
TASK_PP(16'hADCD,4);
TASK_PP(16'hADCE,4);
TASK_PP(16'hADCF,4);
TASK_PP(16'hADD0,4);
TASK_PP(16'hADD1,4);
TASK_PP(16'hADD2,4);
TASK_PP(16'hADD3,4);
TASK_PP(16'hADD4,4);
TASK_PP(16'hADD5,4);
TASK_PP(16'hADD6,4);
TASK_PP(16'hADD7,4);
TASK_PP(16'hADD8,4);
TASK_PP(16'hADD9,4);
TASK_PP(16'hADDA,4);
TASK_PP(16'hADDB,4);
TASK_PP(16'hADDC,4);
TASK_PP(16'hADDD,4);
TASK_PP(16'hADDE,4);
TASK_PP(16'hADDF,4);
TASK_PP(16'hADE0,4);
TASK_PP(16'hADE1,4);
TASK_PP(16'hADE2,4);
TASK_PP(16'hADE3,4);
TASK_PP(16'hADE4,4);
TASK_PP(16'hADE5,4);
TASK_PP(16'hADE6,4);
TASK_PP(16'hADE7,4);
TASK_PP(16'hADE8,4);
TASK_PP(16'hADE9,4);
TASK_PP(16'hADEA,4);
TASK_PP(16'hADEB,4);
TASK_PP(16'hADEC,4);
TASK_PP(16'hADED,4);
TASK_PP(16'hADEE,4);
TASK_PP(16'hADEF,4);
TASK_PP(16'hADF0,4);
TASK_PP(16'hADF1,4);
TASK_PP(16'hADF2,4);
TASK_PP(16'hADF3,4);
TASK_PP(16'hADF4,4);
TASK_PP(16'hADF5,4);
TASK_PP(16'hADF6,4);
TASK_PP(16'hADF7,4);
TASK_PP(16'hADF8,4);
TASK_PP(16'hADF9,4);
TASK_PP(16'hADFA,4);
TASK_PP(16'hADFB,4);
TASK_PP(16'hADFC,4);
TASK_PP(16'hADFD,4);
TASK_PP(16'hADFE,4);
TASK_PP(16'hADFF,4);
TASK_PP(16'hAE00,4);
TASK_PP(16'hAE01,4);
TASK_PP(16'hAE02,4);
TASK_PP(16'hAE03,4);
TASK_PP(16'hAE04,4);
TASK_PP(16'hAE05,4);
TASK_PP(16'hAE06,4);
TASK_PP(16'hAE07,4);
TASK_PP(16'hAE08,4);
TASK_PP(16'hAE09,4);
TASK_PP(16'hAE0A,4);
TASK_PP(16'hAE0B,4);
TASK_PP(16'hAE0C,4);
TASK_PP(16'hAE0D,4);
TASK_PP(16'hAE0E,4);
TASK_PP(16'hAE0F,4);
TASK_PP(16'hAE10,4);
TASK_PP(16'hAE11,4);
TASK_PP(16'hAE12,4);
TASK_PP(16'hAE13,4);
TASK_PP(16'hAE14,4);
TASK_PP(16'hAE15,4);
TASK_PP(16'hAE16,4);
TASK_PP(16'hAE17,4);
TASK_PP(16'hAE18,4);
TASK_PP(16'hAE19,4);
TASK_PP(16'hAE1A,4);
TASK_PP(16'hAE1B,4);
TASK_PP(16'hAE1C,4);
TASK_PP(16'hAE1D,4);
TASK_PP(16'hAE1E,4);
TASK_PP(16'hAE1F,4);
TASK_PP(16'hAE20,4);
TASK_PP(16'hAE21,4);
TASK_PP(16'hAE22,4);
TASK_PP(16'hAE23,4);
TASK_PP(16'hAE24,4);
TASK_PP(16'hAE25,4);
TASK_PP(16'hAE26,4);
TASK_PP(16'hAE27,4);
TASK_PP(16'hAE28,4);
TASK_PP(16'hAE29,4);
TASK_PP(16'hAE2A,4);
TASK_PP(16'hAE2B,4);
TASK_PP(16'hAE2C,4);
TASK_PP(16'hAE2D,4);
TASK_PP(16'hAE2E,4);
TASK_PP(16'hAE2F,4);
TASK_PP(16'hAE30,4);
TASK_PP(16'hAE31,4);
TASK_PP(16'hAE32,4);
TASK_PP(16'hAE33,4);
TASK_PP(16'hAE34,4);
TASK_PP(16'hAE35,4);
TASK_PP(16'hAE36,4);
TASK_PP(16'hAE37,4);
TASK_PP(16'hAE38,4);
TASK_PP(16'hAE39,4);
TASK_PP(16'hAE3A,4);
TASK_PP(16'hAE3B,4);
TASK_PP(16'hAE3C,4);
TASK_PP(16'hAE3D,4);
TASK_PP(16'hAE3E,4);
TASK_PP(16'hAE3F,4);
TASK_PP(16'hAE40,4);
TASK_PP(16'hAE41,4);
TASK_PP(16'hAE42,4);
TASK_PP(16'hAE43,4);
TASK_PP(16'hAE44,4);
TASK_PP(16'hAE45,4);
TASK_PP(16'hAE46,4);
TASK_PP(16'hAE47,4);
TASK_PP(16'hAE48,4);
TASK_PP(16'hAE49,4);
TASK_PP(16'hAE4A,4);
TASK_PP(16'hAE4B,4);
TASK_PP(16'hAE4C,4);
TASK_PP(16'hAE4D,4);
TASK_PP(16'hAE4E,4);
TASK_PP(16'hAE4F,4);
TASK_PP(16'hAE50,4);
TASK_PP(16'hAE51,4);
TASK_PP(16'hAE52,4);
TASK_PP(16'hAE53,4);
TASK_PP(16'hAE54,4);
TASK_PP(16'hAE55,4);
TASK_PP(16'hAE56,4);
TASK_PP(16'hAE57,4);
TASK_PP(16'hAE58,4);
TASK_PP(16'hAE59,4);
TASK_PP(16'hAE5A,4);
TASK_PP(16'hAE5B,4);
TASK_PP(16'hAE5C,4);
TASK_PP(16'hAE5D,4);
TASK_PP(16'hAE5E,4);
TASK_PP(16'hAE5F,4);
TASK_PP(16'hAE60,4);
TASK_PP(16'hAE61,4);
TASK_PP(16'hAE62,4);
TASK_PP(16'hAE63,4);
TASK_PP(16'hAE64,4);
TASK_PP(16'hAE65,4);
TASK_PP(16'hAE66,4);
TASK_PP(16'hAE67,4);
TASK_PP(16'hAE68,4);
TASK_PP(16'hAE69,4);
TASK_PP(16'hAE6A,4);
TASK_PP(16'hAE6B,4);
TASK_PP(16'hAE6C,4);
TASK_PP(16'hAE6D,4);
TASK_PP(16'hAE6E,4);
TASK_PP(16'hAE6F,4);
TASK_PP(16'hAE70,4);
TASK_PP(16'hAE71,4);
TASK_PP(16'hAE72,4);
TASK_PP(16'hAE73,4);
TASK_PP(16'hAE74,4);
TASK_PP(16'hAE75,4);
TASK_PP(16'hAE76,4);
TASK_PP(16'hAE77,4);
TASK_PP(16'hAE78,4);
TASK_PP(16'hAE79,4);
TASK_PP(16'hAE7A,4);
TASK_PP(16'hAE7B,4);
TASK_PP(16'hAE7C,4);
TASK_PP(16'hAE7D,4);
TASK_PP(16'hAE7E,4);
TASK_PP(16'hAE7F,4);
TASK_PP(16'hAE80,4);
TASK_PP(16'hAE81,4);
TASK_PP(16'hAE82,4);
TASK_PP(16'hAE83,4);
TASK_PP(16'hAE84,4);
TASK_PP(16'hAE85,4);
TASK_PP(16'hAE86,4);
TASK_PP(16'hAE87,4);
TASK_PP(16'hAE88,4);
TASK_PP(16'hAE89,4);
TASK_PP(16'hAE8A,4);
TASK_PP(16'hAE8B,4);
TASK_PP(16'hAE8C,4);
TASK_PP(16'hAE8D,4);
TASK_PP(16'hAE8E,4);
TASK_PP(16'hAE8F,4);
TASK_PP(16'hAE90,4);
TASK_PP(16'hAE91,4);
TASK_PP(16'hAE92,4);
TASK_PP(16'hAE93,4);
TASK_PP(16'hAE94,4);
TASK_PP(16'hAE95,4);
TASK_PP(16'hAE96,4);
TASK_PP(16'hAE97,4);
TASK_PP(16'hAE98,4);
TASK_PP(16'hAE99,4);
TASK_PP(16'hAE9A,4);
TASK_PP(16'hAE9B,4);
TASK_PP(16'hAE9C,4);
TASK_PP(16'hAE9D,4);
TASK_PP(16'hAE9E,4);
TASK_PP(16'hAE9F,4);
TASK_PP(16'hAEA0,4);
TASK_PP(16'hAEA1,4);
TASK_PP(16'hAEA2,4);
TASK_PP(16'hAEA3,4);
TASK_PP(16'hAEA4,4);
TASK_PP(16'hAEA5,4);
TASK_PP(16'hAEA6,4);
TASK_PP(16'hAEA7,4);
TASK_PP(16'hAEA8,4);
TASK_PP(16'hAEA9,4);
TASK_PP(16'hAEAA,4);
TASK_PP(16'hAEAB,4);
TASK_PP(16'hAEAC,4);
TASK_PP(16'hAEAD,4);
TASK_PP(16'hAEAE,4);
TASK_PP(16'hAEAF,4);
TASK_PP(16'hAEB0,4);
TASK_PP(16'hAEB1,4);
TASK_PP(16'hAEB2,4);
TASK_PP(16'hAEB3,4);
TASK_PP(16'hAEB4,4);
TASK_PP(16'hAEB5,4);
TASK_PP(16'hAEB6,4);
TASK_PP(16'hAEB7,4);
TASK_PP(16'hAEB8,4);
TASK_PP(16'hAEB9,4);
TASK_PP(16'hAEBA,4);
TASK_PP(16'hAEBB,4);
TASK_PP(16'hAEBC,4);
TASK_PP(16'hAEBD,4);
TASK_PP(16'hAEBE,4);
TASK_PP(16'hAEBF,4);
TASK_PP(16'hAEC0,4);
TASK_PP(16'hAEC1,4);
TASK_PP(16'hAEC2,4);
TASK_PP(16'hAEC3,4);
TASK_PP(16'hAEC4,4);
TASK_PP(16'hAEC5,4);
TASK_PP(16'hAEC6,4);
TASK_PP(16'hAEC7,4);
TASK_PP(16'hAEC8,4);
TASK_PP(16'hAEC9,4);
TASK_PP(16'hAECA,4);
TASK_PP(16'hAECB,4);
TASK_PP(16'hAECC,4);
TASK_PP(16'hAECD,4);
TASK_PP(16'hAECE,4);
TASK_PP(16'hAECF,4);
TASK_PP(16'hAED0,4);
TASK_PP(16'hAED1,4);
TASK_PP(16'hAED2,4);
TASK_PP(16'hAED3,4);
TASK_PP(16'hAED4,4);
TASK_PP(16'hAED5,4);
TASK_PP(16'hAED6,4);
TASK_PP(16'hAED7,4);
TASK_PP(16'hAED8,4);
TASK_PP(16'hAED9,4);
TASK_PP(16'hAEDA,4);
TASK_PP(16'hAEDB,4);
TASK_PP(16'hAEDC,4);
TASK_PP(16'hAEDD,4);
TASK_PP(16'hAEDE,4);
TASK_PP(16'hAEDF,4);
TASK_PP(16'hAEE0,4);
TASK_PP(16'hAEE1,4);
TASK_PP(16'hAEE2,4);
TASK_PP(16'hAEE3,4);
TASK_PP(16'hAEE4,4);
TASK_PP(16'hAEE5,4);
TASK_PP(16'hAEE6,4);
TASK_PP(16'hAEE7,4);
TASK_PP(16'hAEE8,4);
TASK_PP(16'hAEE9,4);
TASK_PP(16'hAEEA,4);
TASK_PP(16'hAEEB,4);
TASK_PP(16'hAEEC,4);
TASK_PP(16'hAEED,4);
TASK_PP(16'hAEEE,4);
TASK_PP(16'hAEEF,4);
TASK_PP(16'hAEF0,4);
TASK_PP(16'hAEF1,4);
TASK_PP(16'hAEF2,4);
TASK_PP(16'hAEF3,4);
TASK_PP(16'hAEF4,4);
TASK_PP(16'hAEF5,4);
TASK_PP(16'hAEF6,4);
TASK_PP(16'hAEF7,4);
TASK_PP(16'hAEF8,4);
TASK_PP(16'hAEF9,4);
TASK_PP(16'hAEFA,4);
TASK_PP(16'hAEFB,4);
TASK_PP(16'hAEFC,4);
TASK_PP(16'hAEFD,4);
TASK_PP(16'hAEFE,4);
TASK_PP(16'hAEFF,4);
TASK_PP(16'hAF00,4);
TASK_PP(16'hAF01,4);
TASK_PP(16'hAF02,4);
TASK_PP(16'hAF03,4);
TASK_PP(16'hAF04,4);
TASK_PP(16'hAF05,4);
TASK_PP(16'hAF06,4);
TASK_PP(16'hAF07,4);
TASK_PP(16'hAF08,4);
TASK_PP(16'hAF09,4);
TASK_PP(16'hAF0A,4);
TASK_PP(16'hAF0B,4);
TASK_PP(16'hAF0C,4);
TASK_PP(16'hAF0D,4);
TASK_PP(16'hAF0E,4);
TASK_PP(16'hAF0F,4);
TASK_PP(16'hAF10,4);
TASK_PP(16'hAF11,4);
TASK_PP(16'hAF12,4);
TASK_PP(16'hAF13,4);
TASK_PP(16'hAF14,4);
TASK_PP(16'hAF15,4);
TASK_PP(16'hAF16,4);
TASK_PP(16'hAF17,4);
TASK_PP(16'hAF18,4);
TASK_PP(16'hAF19,4);
TASK_PP(16'hAF1A,4);
TASK_PP(16'hAF1B,4);
TASK_PP(16'hAF1C,4);
TASK_PP(16'hAF1D,4);
TASK_PP(16'hAF1E,4);
TASK_PP(16'hAF1F,4);
TASK_PP(16'hAF20,4);
TASK_PP(16'hAF21,4);
TASK_PP(16'hAF22,4);
TASK_PP(16'hAF23,4);
TASK_PP(16'hAF24,4);
TASK_PP(16'hAF25,4);
TASK_PP(16'hAF26,4);
TASK_PP(16'hAF27,4);
TASK_PP(16'hAF28,4);
TASK_PP(16'hAF29,4);
TASK_PP(16'hAF2A,4);
TASK_PP(16'hAF2B,4);
TASK_PP(16'hAF2C,4);
TASK_PP(16'hAF2D,4);
TASK_PP(16'hAF2E,4);
TASK_PP(16'hAF2F,4);
TASK_PP(16'hAF30,4);
TASK_PP(16'hAF31,4);
TASK_PP(16'hAF32,4);
TASK_PP(16'hAF33,4);
TASK_PP(16'hAF34,4);
TASK_PP(16'hAF35,4);
TASK_PP(16'hAF36,4);
TASK_PP(16'hAF37,4);
TASK_PP(16'hAF38,4);
TASK_PP(16'hAF39,4);
TASK_PP(16'hAF3A,4);
TASK_PP(16'hAF3B,4);
TASK_PP(16'hAF3C,4);
TASK_PP(16'hAF3D,4);
TASK_PP(16'hAF3E,4);
TASK_PP(16'hAF3F,4);
TASK_PP(16'hAF40,4);
TASK_PP(16'hAF41,4);
TASK_PP(16'hAF42,4);
TASK_PP(16'hAF43,4);
TASK_PP(16'hAF44,4);
TASK_PP(16'hAF45,4);
TASK_PP(16'hAF46,4);
TASK_PP(16'hAF47,4);
TASK_PP(16'hAF48,4);
TASK_PP(16'hAF49,4);
TASK_PP(16'hAF4A,4);
TASK_PP(16'hAF4B,4);
TASK_PP(16'hAF4C,4);
TASK_PP(16'hAF4D,4);
TASK_PP(16'hAF4E,4);
TASK_PP(16'hAF4F,4);
TASK_PP(16'hAF50,4);
TASK_PP(16'hAF51,4);
TASK_PP(16'hAF52,4);
TASK_PP(16'hAF53,4);
TASK_PP(16'hAF54,4);
TASK_PP(16'hAF55,4);
TASK_PP(16'hAF56,4);
TASK_PP(16'hAF57,4);
TASK_PP(16'hAF58,4);
TASK_PP(16'hAF59,4);
TASK_PP(16'hAF5A,4);
TASK_PP(16'hAF5B,4);
TASK_PP(16'hAF5C,4);
TASK_PP(16'hAF5D,4);
TASK_PP(16'hAF5E,4);
TASK_PP(16'hAF5F,4);
TASK_PP(16'hAF60,4);
TASK_PP(16'hAF61,4);
TASK_PP(16'hAF62,4);
TASK_PP(16'hAF63,4);
TASK_PP(16'hAF64,4);
TASK_PP(16'hAF65,4);
TASK_PP(16'hAF66,4);
TASK_PP(16'hAF67,4);
TASK_PP(16'hAF68,4);
TASK_PP(16'hAF69,4);
TASK_PP(16'hAF6A,4);
TASK_PP(16'hAF6B,4);
TASK_PP(16'hAF6C,4);
TASK_PP(16'hAF6D,4);
TASK_PP(16'hAF6E,4);
TASK_PP(16'hAF6F,4);
TASK_PP(16'hAF70,4);
TASK_PP(16'hAF71,4);
TASK_PP(16'hAF72,4);
TASK_PP(16'hAF73,4);
TASK_PP(16'hAF74,4);
TASK_PP(16'hAF75,4);
TASK_PP(16'hAF76,4);
TASK_PP(16'hAF77,4);
TASK_PP(16'hAF78,4);
TASK_PP(16'hAF79,4);
TASK_PP(16'hAF7A,4);
TASK_PP(16'hAF7B,4);
TASK_PP(16'hAF7C,4);
TASK_PP(16'hAF7D,4);
TASK_PP(16'hAF7E,4);
TASK_PP(16'hAF7F,4);
TASK_PP(16'hAF80,4);
TASK_PP(16'hAF81,4);
TASK_PP(16'hAF82,4);
TASK_PP(16'hAF83,4);
TASK_PP(16'hAF84,4);
TASK_PP(16'hAF85,4);
TASK_PP(16'hAF86,4);
TASK_PP(16'hAF87,4);
TASK_PP(16'hAF88,4);
TASK_PP(16'hAF89,4);
TASK_PP(16'hAF8A,4);
TASK_PP(16'hAF8B,4);
TASK_PP(16'hAF8C,4);
TASK_PP(16'hAF8D,4);
TASK_PP(16'hAF8E,4);
TASK_PP(16'hAF8F,4);
TASK_PP(16'hAF90,4);
TASK_PP(16'hAF91,4);
TASK_PP(16'hAF92,4);
TASK_PP(16'hAF93,4);
TASK_PP(16'hAF94,4);
TASK_PP(16'hAF95,4);
TASK_PP(16'hAF96,4);
TASK_PP(16'hAF97,4);
TASK_PP(16'hAF98,4);
TASK_PP(16'hAF99,4);
TASK_PP(16'hAF9A,4);
TASK_PP(16'hAF9B,4);
TASK_PP(16'hAF9C,4);
TASK_PP(16'hAF9D,4);
TASK_PP(16'hAF9E,4);
TASK_PP(16'hAF9F,4);
TASK_PP(16'hAFA0,4);
TASK_PP(16'hAFA1,4);
TASK_PP(16'hAFA2,4);
TASK_PP(16'hAFA3,4);
TASK_PP(16'hAFA4,4);
TASK_PP(16'hAFA5,4);
TASK_PP(16'hAFA6,4);
TASK_PP(16'hAFA7,4);
TASK_PP(16'hAFA8,4);
TASK_PP(16'hAFA9,4);
TASK_PP(16'hAFAA,4);
TASK_PP(16'hAFAB,4);
TASK_PP(16'hAFAC,4);
TASK_PP(16'hAFAD,4);
TASK_PP(16'hAFAE,4);
TASK_PP(16'hAFAF,4);
TASK_PP(16'hAFB0,4);
TASK_PP(16'hAFB1,4);
TASK_PP(16'hAFB2,4);
TASK_PP(16'hAFB3,4);
TASK_PP(16'hAFB4,4);
TASK_PP(16'hAFB5,4);
TASK_PP(16'hAFB6,4);
TASK_PP(16'hAFB7,4);
TASK_PP(16'hAFB8,4);
TASK_PP(16'hAFB9,4);
TASK_PP(16'hAFBA,4);
TASK_PP(16'hAFBB,4);
TASK_PP(16'hAFBC,4);
TASK_PP(16'hAFBD,4);
TASK_PP(16'hAFBE,4);
TASK_PP(16'hAFBF,4);
TASK_PP(16'hAFC0,4);
TASK_PP(16'hAFC1,4);
TASK_PP(16'hAFC2,4);
TASK_PP(16'hAFC3,4);
TASK_PP(16'hAFC4,4);
TASK_PP(16'hAFC5,4);
TASK_PP(16'hAFC6,4);
TASK_PP(16'hAFC7,4);
TASK_PP(16'hAFC8,4);
TASK_PP(16'hAFC9,4);
TASK_PP(16'hAFCA,4);
TASK_PP(16'hAFCB,4);
TASK_PP(16'hAFCC,4);
TASK_PP(16'hAFCD,4);
TASK_PP(16'hAFCE,4);
TASK_PP(16'hAFCF,4);
TASK_PP(16'hAFD0,4);
TASK_PP(16'hAFD1,4);
TASK_PP(16'hAFD2,4);
TASK_PP(16'hAFD3,4);
TASK_PP(16'hAFD4,4);
TASK_PP(16'hAFD5,4);
TASK_PP(16'hAFD6,4);
TASK_PP(16'hAFD7,4);
TASK_PP(16'hAFD8,4);
TASK_PP(16'hAFD9,4);
TASK_PP(16'hAFDA,4);
TASK_PP(16'hAFDB,4);
TASK_PP(16'hAFDC,4);
TASK_PP(16'hAFDD,4);
TASK_PP(16'hAFDE,4);
TASK_PP(16'hAFDF,4);
TASK_PP(16'hAFE0,4);
TASK_PP(16'hAFE1,4);
TASK_PP(16'hAFE2,4);
TASK_PP(16'hAFE3,4);
TASK_PP(16'hAFE4,4);
TASK_PP(16'hAFE5,4);
TASK_PP(16'hAFE6,4);
TASK_PP(16'hAFE7,4);
TASK_PP(16'hAFE8,4);
TASK_PP(16'hAFE9,4);
TASK_PP(16'hAFEA,4);
TASK_PP(16'hAFEB,4);
TASK_PP(16'hAFEC,4);
TASK_PP(16'hAFED,4);
TASK_PP(16'hAFEE,4);
TASK_PP(16'hAFEF,4);
TASK_PP(16'hAFF0,4);
TASK_PP(16'hAFF1,4);
TASK_PP(16'hAFF2,4);
TASK_PP(16'hAFF3,4);
TASK_PP(16'hAFF4,4);
TASK_PP(16'hAFF5,4);
TASK_PP(16'hAFF6,4);
TASK_PP(16'hAFF7,4);
TASK_PP(16'hAFF8,4);
TASK_PP(16'hAFF9,4);
TASK_PP(16'hAFFA,4);
TASK_PP(16'hAFFB,4);
TASK_PP(16'hAFFC,4);
TASK_PP(16'hAFFD,4);
TASK_PP(16'hAFFE,4);
TASK_PP(16'hAFFF,4);
TASK_PP(16'hB000,4);
TASK_PP(16'hB001,4);
TASK_PP(16'hB002,4);
TASK_PP(16'hB003,4);
TASK_PP(16'hB004,4);
TASK_PP(16'hB005,4);
TASK_PP(16'hB006,4);
TASK_PP(16'hB007,4);
TASK_PP(16'hB008,4);
TASK_PP(16'hB009,4);
TASK_PP(16'hB00A,4);
TASK_PP(16'hB00B,4);
TASK_PP(16'hB00C,4);
TASK_PP(16'hB00D,4);
TASK_PP(16'hB00E,4);
TASK_PP(16'hB00F,4);
TASK_PP(16'hB010,4);
TASK_PP(16'hB011,4);
TASK_PP(16'hB012,4);
TASK_PP(16'hB013,4);
TASK_PP(16'hB014,4);
TASK_PP(16'hB015,4);
TASK_PP(16'hB016,4);
TASK_PP(16'hB017,4);
TASK_PP(16'hB018,4);
TASK_PP(16'hB019,4);
TASK_PP(16'hB01A,4);
TASK_PP(16'hB01B,4);
TASK_PP(16'hB01C,4);
TASK_PP(16'hB01D,4);
TASK_PP(16'hB01E,4);
TASK_PP(16'hB01F,4);
TASK_PP(16'hB020,4);
TASK_PP(16'hB021,4);
TASK_PP(16'hB022,4);
TASK_PP(16'hB023,4);
TASK_PP(16'hB024,4);
TASK_PP(16'hB025,4);
TASK_PP(16'hB026,4);
TASK_PP(16'hB027,4);
TASK_PP(16'hB028,4);
TASK_PP(16'hB029,4);
TASK_PP(16'hB02A,4);
TASK_PP(16'hB02B,4);
TASK_PP(16'hB02C,4);
TASK_PP(16'hB02D,4);
TASK_PP(16'hB02E,4);
TASK_PP(16'hB02F,4);
TASK_PP(16'hB030,4);
TASK_PP(16'hB031,4);
TASK_PP(16'hB032,4);
TASK_PP(16'hB033,4);
TASK_PP(16'hB034,4);
TASK_PP(16'hB035,4);
TASK_PP(16'hB036,4);
TASK_PP(16'hB037,4);
TASK_PP(16'hB038,4);
TASK_PP(16'hB039,4);
TASK_PP(16'hB03A,4);
TASK_PP(16'hB03B,4);
TASK_PP(16'hB03C,4);
TASK_PP(16'hB03D,4);
TASK_PP(16'hB03E,4);
TASK_PP(16'hB03F,4);
TASK_PP(16'hB040,4);
TASK_PP(16'hB041,4);
TASK_PP(16'hB042,4);
TASK_PP(16'hB043,4);
TASK_PP(16'hB044,4);
TASK_PP(16'hB045,4);
TASK_PP(16'hB046,4);
TASK_PP(16'hB047,4);
TASK_PP(16'hB048,4);
TASK_PP(16'hB049,4);
TASK_PP(16'hB04A,4);
TASK_PP(16'hB04B,4);
TASK_PP(16'hB04C,4);
TASK_PP(16'hB04D,4);
TASK_PP(16'hB04E,4);
TASK_PP(16'hB04F,4);
TASK_PP(16'hB050,4);
TASK_PP(16'hB051,4);
TASK_PP(16'hB052,4);
TASK_PP(16'hB053,4);
TASK_PP(16'hB054,4);
TASK_PP(16'hB055,4);
TASK_PP(16'hB056,4);
TASK_PP(16'hB057,4);
TASK_PP(16'hB058,4);
TASK_PP(16'hB059,4);
TASK_PP(16'hB05A,4);
TASK_PP(16'hB05B,4);
TASK_PP(16'hB05C,4);
TASK_PP(16'hB05D,4);
TASK_PP(16'hB05E,4);
TASK_PP(16'hB05F,4);
TASK_PP(16'hB060,4);
TASK_PP(16'hB061,4);
TASK_PP(16'hB062,4);
TASK_PP(16'hB063,4);
TASK_PP(16'hB064,4);
TASK_PP(16'hB065,4);
TASK_PP(16'hB066,4);
TASK_PP(16'hB067,4);
TASK_PP(16'hB068,4);
TASK_PP(16'hB069,4);
TASK_PP(16'hB06A,4);
TASK_PP(16'hB06B,4);
TASK_PP(16'hB06C,4);
TASK_PP(16'hB06D,4);
TASK_PP(16'hB06E,4);
TASK_PP(16'hB06F,4);
TASK_PP(16'hB070,4);
TASK_PP(16'hB071,4);
TASK_PP(16'hB072,4);
TASK_PP(16'hB073,4);
TASK_PP(16'hB074,4);
TASK_PP(16'hB075,4);
TASK_PP(16'hB076,4);
TASK_PP(16'hB077,4);
TASK_PP(16'hB078,4);
TASK_PP(16'hB079,4);
TASK_PP(16'hB07A,4);
TASK_PP(16'hB07B,4);
TASK_PP(16'hB07C,4);
TASK_PP(16'hB07D,4);
TASK_PP(16'hB07E,4);
TASK_PP(16'hB07F,4);
TASK_PP(16'hB080,4);
TASK_PP(16'hB081,4);
TASK_PP(16'hB082,4);
TASK_PP(16'hB083,4);
TASK_PP(16'hB084,4);
TASK_PP(16'hB085,4);
TASK_PP(16'hB086,4);
TASK_PP(16'hB087,4);
TASK_PP(16'hB088,4);
TASK_PP(16'hB089,4);
TASK_PP(16'hB08A,4);
TASK_PP(16'hB08B,4);
TASK_PP(16'hB08C,4);
TASK_PP(16'hB08D,4);
TASK_PP(16'hB08E,4);
TASK_PP(16'hB08F,4);
TASK_PP(16'hB090,4);
TASK_PP(16'hB091,4);
TASK_PP(16'hB092,4);
TASK_PP(16'hB093,4);
TASK_PP(16'hB094,4);
TASK_PP(16'hB095,4);
TASK_PP(16'hB096,4);
TASK_PP(16'hB097,4);
TASK_PP(16'hB098,4);
TASK_PP(16'hB099,4);
TASK_PP(16'hB09A,4);
TASK_PP(16'hB09B,4);
TASK_PP(16'hB09C,4);
TASK_PP(16'hB09D,4);
TASK_PP(16'hB09E,4);
TASK_PP(16'hB09F,4);
TASK_PP(16'hB0A0,4);
TASK_PP(16'hB0A1,4);
TASK_PP(16'hB0A2,4);
TASK_PP(16'hB0A3,4);
TASK_PP(16'hB0A4,4);
TASK_PP(16'hB0A5,4);
TASK_PP(16'hB0A6,4);
TASK_PP(16'hB0A7,4);
TASK_PP(16'hB0A8,4);
TASK_PP(16'hB0A9,4);
TASK_PP(16'hB0AA,4);
TASK_PP(16'hB0AB,4);
TASK_PP(16'hB0AC,4);
TASK_PP(16'hB0AD,4);
TASK_PP(16'hB0AE,4);
TASK_PP(16'hB0AF,4);
TASK_PP(16'hB0B0,4);
TASK_PP(16'hB0B1,4);
TASK_PP(16'hB0B2,4);
TASK_PP(16'hB0B3,4);
TASK_PP(16'hB0B4,4);
TASK_PP(16'hB0B5,4);
TASK_PP(16'hB0B6,4);
TASK_PP(16'hB0B7,4);
TASK_PP(16'hB0B8,4);
TASK_PP(16'hB0B9,4);
TASK_PP(16'hB0BA,4);
TASK_PP(16'hB0BB,4);
TASK_PP(16'hB0BC,4);
TASK_PP(16'hB0BD,4);
TASK_PP(16'hB0BE,4);
TASK_PP(16'hB0BF,4);
TASK_PP(16'hB0C0,4);
TASK_PP(16'hB0C1,4);
TASK_PP(16'hB0C2,4);
TASK_PP(16'hB0C3,4);
TASK_PP(16'hB0C4,4);
TASK_PP(16'hB0C5,4);
TASK_PP(16'hB0C6,4);
TASK_PP(16'hB0C7,4);
TASK_PP(16'hB0C8,4);
TASK_PP(16'hB0C9,4);
TASK_PP(16'hB0CA,4);
TASK_PP(16'hB0CB,4);
TASK_PP(16'hB0CC,4);
TASK_PP(16'hB0CD,4);
TASK_PP(16'hB0CE,4);
TASK_PP(16'hB0CF,4);
TASK_PP(16'hB0D0,4);
TASK_PP(16'hB0D1,4);
TASK_PP(16'hB0D2,4);
TASK_PP(16'hB0D3,4);
TASK_PP(16'hB0D4,4);
TASK_PP(16'hB0D5,4);
TASK_PP(16'hB0D6,4);
TASK_PP(16'hB0D7,4);
TASK_PP(16'hB0D8,4);
TASK_PP(16'hB0D9,4);
TASK_PP(16'hB0DA,4);
TASK_PP(16'hB0DB,4);
TASK_PP(16'hB0DC,4);
TASK_PP(16'hB0DD,4);
TASK_PP(16'hB0DE,4);
TASK_PP(16'hB0DF,4);
TASK_PP(16'hB0E0,4);
TASK_PP(16'hB0E1,4);
TASK_PP(16'hB0E2,4);
TASK_PP(16'hB0E3,4);
TASK_PP(16'hB0E4,4);
TASK_PP(16'hB0E5,4);
TASK_PP(16'hB0E6,4);
TASK_PP(16'hB0E7,4);
TASK_PP(16'hB0E8,4);
TASK_PP(16'hB0E9,4);
TASK_PP(16'hB0EA,4);
TASK_PP(16'hB0EB,4);
TASK_PP(16'hB0EC,4);
TASK_PP(16'hB0ED,4);
TASK_PP(16'hB0EE,4);
TASK_PP(16'hB0EF,4);
TASK_PP(16'hB0F0,4);
TASK_PP(16'hB0F1,4);
TASK_PP(16'hB0F2,4);
TASK_PP(16'hB0F3,4);
TASK_PP(16'hB0F4,4);
TASK_PP(16'hB0F5,4);
TASK_PP(16'hB0F6,4);
TASK_PP(16'hB0F7,4);
TASK_PP(16'hB0F8,4);
TASK_PP(16'hB0F9,4);
TASK_PP(16'hB0FA,4);
TASK_PP(16'hB0FB,4);
TASK_PP(16'hB0FC,4);
TASK_PP(16'hB0FD,4);
TASK_PP(16'hB0FE,4);
TASK_PP(16'hB0FF,4);
TASK_PP(16'hB100,4);
TASK_PP(16'hB101,4);
TASK_PP(16'hB102,4);
TASK_PP(16'hB103,4);
TASK_PP(16'hB104,4);
TASK_PP(16'hB105,4);
TASK_PP(16'hB106,4);
TASK_PP(16'hB107,4);
TASK_PP(16'hB108,4);
TASK_PP(16'hB109,4);
TASK_PP(16'hB10A,4);
TASK_PP(16'hB10B,4);
TASK_PP(16'hB10C,4);
TASK_PP(16'hB10D,4);
TASK_PP(16'hB10E,4);
TASK_PP(16'hB10F,4);
TASK_PP(16'hB110,4);
TASK_PP(16'hB111,4);
TASK_PP(16'hB112,4);
TASK_PP(16'hB113,4);
TASK_PP(16'hB114,4);
TASK_PP(16'hB115,4);
TASK_PP(16'hB116,4);
TASK_PP(16'hB117,4);
TASK_PP(16'hB118,4);
TASK_PP(16'hB119,4);
TASK_PP(16'hB11A,4);
TASK_PP(16'hB11B,4);
TASK_PP(16'hB11C,4);
TASK_PP(16'hB11D,4);
TASK_PP(16'hB11E,4);
TASK_PP(16'hB11F,4);
TASK_PP(16'hB120,4);
TASK_PP(16'hB121,4);
TASK_PP(16'hB122,4);
TASK_PP(16'hB123,4);
TASK_PP(16'hB124,4);
TASK_PP(16'hB125,4);
TASK_PP(16'hB126,4);
TASK_PP(16'hB127,4);
TASK_PP(16'hB128,4);
TASK_PP(16'hB129,4);
TASK_PP(16'hB12A,4);
TASK_PP(16'hB12B,4);
TASK_PP(16'hB12C,4);
TASK_PP(16'hB12D,4);
TASK_PP(16'hB12E,4);
TASK_PP(16'hB12F,4);
TASK_PP(16'hB130,4);
TASK_PP(16'hB131,4);
TASK_PP(16'hB132,4);
TASK_PP(16'hB133,4);
TASK_PP(16'hB134,4);
TASK_PP(16'hB135,4);
TASK_PP(16'hB136,4);
TASK_PP(16'hB137,4);
TASK_PP(16'hB138,4);
TASK_PP(16'hB139,4);
TASK_PP(16'hB13A,4);
TASK_PP(16'hB13B,4);
TASK_PP(16'hB13C,4);
TASK_PP(16'hB13D,4);
TASK_PP(16'hB13E,4);
TASK_PP(16'hB13F,4);
TASK_PP(16'hB140,4);
TASK_PP(16'hB141,4);
TASK_PP(16'hB142,4);
TASK_PP(16'hB143,4);
TASK_PP(16'hB144,4);
TASK_PP(16'hB145,4);
TASK_PP(16'hB146,4);
TASK_PP(16'hB147,4);
TASK_PP(16'hB148,4);
TASK_PP(16'hB149,4);
TASK_PP(16'hB14A,4);
TASK_PP(16'hB14B,4);
TASK_PP(16'hB14C,4);
TASK_PP(16'hB14D,4);
TASK_PP(16'hB14E,4);
TASK_PP(16'hB14F,4);
TASK_PP(16'hB150,4);
TASK_PP(16'hB151,4);
TASK_PP(16'hB152,4);
TASK_PP(16'hB153,4);
TASK_PP(16'hB154,4);
TASK_PP(16'hB155,4);
TASK_PP(16'hB156,4);
TASK_PP(16'hB157,4);
TASK_PP(16'hB158,4);
TASK_PP(16'hB159,4);
TASK_PP(16'hB15A,4);
TASK_PP(16'hB15B,4);
TASK_PP(16'hB15C,4);
TASK_PP(16'hB15D,4);
TASK_PP(16'hB15E,4);
TASK_PP(16'hB15F,4);
TASK_PP(16'hB160,4);
TASK_PP(16'hB161,4);
TASK_PP(16'hB162,4);
TASK_PP(16'hB163,4);
TASK_PP(16'hB164,4);
TASK_PP(16'hB165,4);
TASK_PP(16'hB166,4);
TASK_PP(16'hB167,4);
TASK_PP(16'hB168,4);
TASK_PP(16'hB169,4);
TASK_PP(16'hB16A,4);
TASK_PP(16'hB16B,4);
TASK_PP(16'hB16C,4);
TASK_PP(16'hB16D,4);
TASK_PP(16'hB16E,4);
TASK_PP(16'hB16F,4);
TASK_PP(16'hB170,4);
TASK_PP(16'hB171,4);
TASK_PP(16'hB172,4);
TASK_PP(16'hB173,4);
TASK_PP(16'hB174,4);
TASK_PP(16'hB175,4);
TASK_PP(16'hB176,4);
TASK_PP(16'hB177,4);
TASK_PP(16'hB178,4);
TASK_PP(16'hB179,4);
TASK_PP(16'hB17A,4);
TASK_PP(16'hB17B,4);
TASK_PP(16'hB17C,4);
TASK_PP(16'hB17D,4);
TASK_PP(16'hB17E,4);
TASK_PP(16'hB17F,4);
TASK_PP(16'hB180,4);
TASK_PP(16'hB181,4);
TASK_PP(16'hB182,4);
TASK_PP(16'hB183,4);
TASK_PP(16'hB184,4);
TASK_PP(16'hB185,4);
TASK_PP(16'hB186,4);
TASK_PP(16'hB187,4);
TASK_PP(16'hB188,4);
TASK_PP(16'hB189,4);
TASK_PP(16'hB18A,4);
TASK_PP(16'hB18B,4);
TASK_PP(16'hB18C,4);
TASK_PP(16'hB18D,4);
TASK_PP(16'hB18E,4);
TASK_PP(16'hB18F,4);
TASK_PP(16'hB190,4);
TASK_PP(16'hB191,4);
TASK_PP(16'hB192,4);
TASK_PP(16'hB193,4);
TASK_PP(16'hB194,4);
TASK_PP(16'hB195,4);
TASK_PP(16'hB196,4);
TASK_PP(16'hB197,4);
TASK_PP(16'hB198,4);
TASK_PP(16'hB199,4);
TASK_PP(16'hB19A,4);
TASK_PP(16'hB19B,4);
TASK_PP(16'hB19C,4);
TASK_PP(16'hB19D,4);
TASK_PP(16'hB19E,4);
TASK_PP(16'hB19F,4);
TASK_PP(16'hB1A0,4);
TASK_PP(16'hB1A1,4);
TASK_PP(16'hB1A2,4);
TASK_PP(16'hB1A3,4);
TASK_PP(16'hB1A4,4);
TASK_PP(16'hB1A5,4);
TASK_PP(16'hB1A6,4);
TASK_PP(16'hB1A7,4);
TASK_PP(16'hB1A8,4);
TASK_PP(16'hB1A9,4);
TASK_PP(16'hB1AA,4);
TASK_PP(16'hB1AB,4);
TASK_PP(16'hB1AC,4);
TASK_PP(16'hB1AD,4);
TASK_PP(16'hB1AE,4);
TASK_PP(16'hB1AF,4);
TASK_PP(16'hB1B0,4);
TASK_PP(16'hB1B1,4);
TASK_PP(16'hB1B2,4);
TASK_PP(16'hB1B3,4);
TASK_PP(16'hB1B4,4);
TASK_PP(16'hB1B5,4);
TASK_PP(16'hB1B6,4);
TASK_PP(16'hB1B7,4);
TASK_PP(16'hB1B8,4);
TASK_PP(16'hB1B9,4);
TASK_PP(16'hB1BA,4);
TASK_PP(16'hB1BB,4);
TASK_PP(16'hB1BC,4);
TASK_PP(16'hB1BD,4);
TASK_PP(16'hB1BE,4);
TASK_PP(16'hB1BF,4);
TASK_PP(16'hB1C0,4);
TASK_PP(16'hB1C1,4);
TASK_PP(16'hB1C2,4);
TASK_PP(16'hB1C3,4);
TASK_PP(16'hB1C4,4);
TASK_PP(16'hB1C5,4);
TASK_PP(16'hB1C6,4);
TASK_PP(16'hB1C7,4);
TASK_PP(16'hB1C8,4);
TASK_PP(16'hB1C9,4);
TASK_PP(16'hB1CA,4);
TASK_PP(16'hB1CB,4);
TASK_PP(16'hB1CC,4);
TASK_PP(16'hB1CD,4);
TASK_PP(16'hB1CE,4);
TASK_PP(16'hB1CF,4);
TASK_PP(16'hB1D0,4);
TASK_PP(16'hB1D1,4);
TASK_PP(16'hB1D2,4);
TASK_PP(16'hB1D3,4);
TASK_PP(16'hB1D4,4);
TASK_PP(16'hB1D5,4);
TASK_PP(16'hB1D6,4);
TASK_PP(16'hB1D7,4);
TASK_PP(16'hB1D8,4);
TASK_PP(16'hB1D9,4);
TASK_PP(16'hB1DA,4);
TASK_PP(16'hB1DB,4);
TASK_PP(16'hB1DC,4);
TASK_PP(16'hB1DD,4);
TASK_PP(16'hB1DE,4);
TASK_PP(16'hB1DF,4);
TASK_PP(16'hB1E0,4);
TASK_PP(16'hB1E1,4);
TASK_PP(16'hB1E2,4);
TASK_PP(16'hB1E3,4);
TASK_PP(16'hB1E4,4);
TASK_PP(16'hB1E5,4);
TASK_PP(16'hB1E6,4);
TASK_PP(16'hB1E7,4);
TASK_PP(16'hB1E8,4);
TASK_PP(16'hB1E9,4);
TASK_PP(16'hB1EA,4);
TASK_PP(16'hB1EB,4);
TASK_PP(16'hB1EC,4);
TASK_PP(16'hB1ED,4);
TASK_PP(16'hB1EE,4);
TASK_PP(16'hB1EF,4);
TASK_PP(16'hB1F0,4);
TASK_PP(16'hB1F1,4);
TASK_PP(16'hB1F2,4);
TASK_PP(16'hB1F3,4);
TASK_PP(16'hB1F4,4);
TASK_PP(16'hB1F5,4);
TASK_PP(16'hB1F6,4);
TASK_PP(16'hB1F7,4);
TASK_PP(16'hB1F8,4);
TASK_PP(16'hB1F9,4);
TASK_PP(16'hB1FA,4);
TASK_PP(16'hB1FB,4);
TASK_PP(16'hB1FC,4);
TASK_PP(16'hB1FD,4);
TASK_PP(16'hB1FE,4);
TASK_PP(16'hB1FF,4);
TASK_PP(16'hB200,4);
TASK_PP(16'hB201,4);
TASK_PP(16'hB202,4);
TASK_PP(16'hB203,4);
TASK_PP(16'hB204,4);
TASK_PP(16'hB205,4);
TASK_PP(16'hB206,4);
TASK_PP(16'hB207,4);
TASK_PP(16'hB208,4);
TASK_PP(16'hB209,4);
TASK_PP(16'hB20A,4);
TASK_PP(16'hB20B,4);
TASK_PP(16'hB20C,4);
TASK_PP(16'hB20D,4);
TASK_PP(16'hB20E,4);
TASK_PP(16'hB20F,4);
TASK_PP(16'hB210,4);
TASK_PP(16'hB211,4);
TASK_PP(16'hB212,4);
TASK_PP(16'hB213,4);
TASK_PP(16'hB214,4);
TASK_PP(16'hB215,4);
TASK_PP(16'hB216,4);
TASK_PP(16'hB217,4);
TASK_PP(16'hB218,4);
TASK_PP(16'hB219,4);
TASK_PP(16'hB21A,4);
TASK_PP(16'hB21B,4);
TASK_PP(16'hB21C,4);
TASK_PP(16'hB21D,4);
TASK_PP(16'hB21E,4);
TASK_PP(16'hB21F,4);
TASK_PP(16'hB220,4);
TASK_PP(16'hB221,4);
TASK_PP(16'hB222,4);
TASK_PP(16'hB223,4);
TASK_PP(16'hB224,4);
TASK_PP(16'hB225,4);
TASK_PP(16'hB226,4);
TASK_PP(16'hB227,4);
TASK_PP(16'hB228,4);
TASK_PP(16'hB229,4);
TASK_PP(16'hB22A,4);
TASK_PP(16'hB22B,4);
TASK_PP(16'hB22C,4);
TASK_PP(16'hB22D,4);
TASK_PP(16'hB22E,4);
TASK_PP(16'hB22F,4);
TASK_PP(16'hB230,4);
TASK_PP(16'hB231,4);
TASK_PP(16'hB232,4);
TASK_PP(16'hB233,4);
TASK_PP(16'hB234,4);
TASK_PP(16'hB235,4);
TASK_PP(16'hB236,4);
TASK_PP(16'hB237,4);
TASK_PP(16'hB238,4);
TASK_PP(16'hB239,4);
TASK_PP(16'hB23A,4);
TASK_PP(16'hB23B,4);
TASK_PP(16'hB23C,4);
TASK_PP(16'hB23D,4);
TASK_PP(16'hB23E,4);
TASK_PP(16'hB23F,4);
TASK_PP(16'hB240,4);
TASK_PP(16'hB241,4);
TASK_PP(16'hB242,4);
TASK_PP(16'hB243,4);
TASK_PP(16'hB244,4);
TASK_PP(16'hB245,4);
TASK_PP(16'hB246,4);
TASK_PP(16'hB247,4);
TASK_PP(16'hB248,4);
TASK_PP(16'hB249,4);
TASK_PP(16'hB24A,4);
TASK_PP(16'hB24B,4);
TASK_PP(16'hB24C,4);
TASK_PP(16'hB24D,4);
TASK_PP(16'hB24E,4);
TASK_PP(16'hB24F,4);
TASK_PP(16'hB250,4);
TASK_PP(16'hB251,4);
TASK_PP(16'hB252,4);
TASK_PP(16'hB253,4);
TASK_PP(16'hB254,4);
TASK_PP(16'hB255,4);
TASK_PP(16'hB256,4);
TASK_PP(16'hB257,4);
TASK_PP(16'hB258,4);
TASK_PP(16'hB259,4);
TASK_PP(16'hB25A,4);
TASK_PP(16'hB25B,4);
TASK_PP(16'hB25C,4);
TASK_PP(16'hB25D,4);
TASK_PP(16'hB25E,4);
TASK_PP(16'hB25F,4);
TASK_PP(16'hB260,4);
TASK_PP(16'hB261,4);
TASK_PP(16'hB262,4);
TASK_PP(16'hB263,4);
TASK_PP(16'hB264,4);
TASK_PP(16'hB265,4);
TASK_PP(16'hB266,4);
TASK_PP(16'hB267,4);
TASK_PP(16'hB268,4);
TASK_PP(16'hB269,4);
TASK_PP(16'hB26A,4);
TASK_PP(16'hB26B,4);
TASK_PP(16'hB26C,4);
TASK_PP(16'hB26D,4);
TASK_PP(16'hB26E,4);
TASK_PP(16'hB26F,4);
TASK_PP(16'hB270,4);
TASK_PP(16'hB271,4);
TASK_PP(16'hB272,4);
TASK_PP(16'hB273,4);
TASK_PP(16'hB274,4);
TASK_PP(16'hB275,4);
TASK_PP(16'hB276,4);
TASK_PP(16'hB277,4);
TASK_PP(16'hB278,4);
TASK_PP(16'hB279,4);
TASK_PP(16'hB27A,4);
TASK_PP(16'hB27B,4);
TASK_PP(16'hB27C,4);
TASK_PP(16'hB27D,4);
TASK_PP(16'hB27E,4);
TASK_PP(16'hB27F,4);
TASK_PP(16'hB280,4);
TASK_PP(16'hB281,4);
TASK_PP(16'hB282,4);
TASK_PP(16'hB283,4);
TASK_PP(16'hB284,4);
TASK_PP(16'hB285,4);
TASK_PP(16'hB286,4);
TASK_PP(16'hB287,4);
TASK_PP(16'hB288,4);
TASK_PP(16'hB289,4);
TASK_PP(16'hB28A,4);
TASK_PP(16'hB28B,4);
TASK_PP(16'hB28C,4);
TASK_PP(16'hB28D,4);
TASK_PP(16'hB28E,4);
TASK_PP(16'hB28F,4);
TASK_PP(16'hB290,4);
TASK_PP(16'hB291,4);
TASK_PP(16'hB292,4);
TASK_PP(16'hB293,4);
TASK_PP(16'hB294,4);
TASK_PP(16'hB295,4);
TASK_PP(16'hB296,4);
TASK_PP(16'hB297,4);
TASK_PP(16'hB298,4);
TASK_PP(16'hB299,4);
TASK_PP(16'hB29A,4);
TASK_PP(16'hB29B,4);
TASK_PP(16'hB29C,4);
TASK_PP(16'hB29D,4);
TASK_PP(16'hB29E,4);
TASK_PP(16'hB29F,4);
TASK_PP(16'hB2A0,4);
TASK_PP(16'hB2A1,4);
TASK_PP(16'hB2A2,4);
TASK_PP(16'hB2A3,4);
TASK_PP(16'hB2A4,4);
TASK_PP(16'hB2A5,4);
TASK_PP(16'hB2A6,4);
TASK_PP(16'hB2A7,4);
TASK_PP(16'hB2A8,4);
TASK_PP(16'hB2A9,4);
TASK_PP(16'hB2AA,4);
TASK_PP(16'hB2AB,4);
TASK_PP(16'hB2AC,4);
TASK_PP(16'hB2AD,4);
TASK_PP(16'hB2AE,4);
TASK_PP(16'hB2AF,4);
TASK_PP(16'hB2B0,4);
TASK_PP(16'hB2B1,4);
TASK_PP(16'hB2B2,4);
TASK_PP(16'hB2B3,4);
TASK_PP(16'hB2B4,4);
TASK_PP(16'hB2B5,4);
TASK_PP(16'hB2B6,4);
TASK_PP(16'hB2B7,4);
TASK_PP(16'hB2B8,4);
TASK_PP(16'hB2B9,4);
TASK_PP(16'hB2BA,4);
TASK_PP(16'hB2BB,4);
TASK_PP(16'hB2BC,4);
TASK_PP(16'hB2BD,4);
TASK_PP(16'hB2BE,4);
TASK_PP(16'hB2BF,4);
TASK_PP(16'hB2C0,4);
TASK_PP(16'hB2C1,4);
TASK_PP(16'hB2C2,4);
TASK_PP(16'hB2C3,4);
TASK_PP(16'hB2C4,4);
TASK_PP(16'hB2C5,4);
TASK_PP(16'hB2C6,4);
TASK_PP(16'hB2C7,4);
TASK_PP(16'hB2C8,4);
TASK_PP(16'hB2C9,4);
TASK_PP(16'hB2CA,4);
TASK_PP(16'hB2CB,4);
TASK_PP(16'hB2CC,4);
TASK_PP(16'hB2CD,4);
TASK_PP(16'hB2CE,4);
TASK_PP(16'hB2CF,4);
TASK_PP(16'hB2D0,4);
TASK_PP(16'hB2D1,4);
TASK_PP(16'hB2D2,4);
TASK_PP(16'hB2D3,4);
TASK_PP(16'hB2D4,4);
TASK_PP(16'hB2D5,4);
TASK_PP(16'hB2D6,4);
TASK_PP(16'hB2D7,4);
TASK_PP(16'hB2D8,4);
TASK_PP(16'hB2D9,4);
TASK_PP(16'hB2DA,4);
TASK_PP(16'hB2DB,4);
TASK_PP(16'hB2DC,4);
TASK_PP(16'hB2DD,4);
TASK_PP(16'hB2DE,4);
TASK_PP(16'hB2DF,4);
TASK_PP(16'hB2E0,4);
TASK_PP(16'hB2E1,4);
TASK_PP(16'hB2E2,4);
TASK_PP(16'hB2E3,4);
TASK_PP(16'hB2E4,4);
TASK_PP(16'hB2E5,4);
TASK_PP(16'hB2E6,4);
TASK_PP(16'hB2E7,4);
TASK_PP(16'hB2E8,4);
TASK_PP(16'hB2E9,4);
TASK_PP(16'hB2EA,4);
TASK_PP(16'hB2EB,4);
TASK_PP(16'hB2EC,4);
TASK_PP(16'hB2ED,4);
TASK_PP(16'hB2EE,4);
TASK_PP(16'hB2EF,4);
TASK_PP(16'hB2F0,4);
TASK_PP(16'hB2F1,4);
TASK_PP(16'hB2F2,4);
TASK_PP(16'hB2F3,4);
TASK_PP(16'hB2F4,4);
TASK_PP(16'hB2F5,4);
TASK_PP(16'hB2F6,4);
TASK_PP(16'hB2F7,4);
TASK_PP(16'hB2F8,4);
TASK_PP(16'hB2F9,4);
TASK_PP(16'hB2FA,4);
TASK_PP(16'hB2FB,4);
TASK_PP(16'hB2FC,4);
TASK_PP(16'hB2FD,4);
TASK_PP(16'hB2FE,4);
TASK_PP(16'hB2FF,4);
TASK_PP(16'hB300,4);
TASK_PP(16'hB301,4);
TASK_PP(16'hB302,4);
TASK_PP(16'hB303,4);
TASK_PP(16'hB304,4);
TASK_PP(16'hB305,4);
TASK_PP(16'hB306,4);
TASK_PP(16'hB307,4);
TASK_PP(16'hB308,4);
TASK_PP(16'hB309,4);
TASK_PP(16'hB30A,4);
TASK_PP(16'hB30B,4);
TASK_PP(16'hB30C,4);
TASK_PP(16'hB30D,4);
TASK_PP(16'hB30E,4);
TASK_PP(16'hB30F,4);
TASK_PP(16'hB310,4);
TASK_PP(16'hB311,4);
TASK_PP(16'hB312,4);
TASK_PP(16'hB313,4);
TASK_PP(16'hB314,4);
TASK_PP(16'hB315,4);
TASK_PP(16'hB316,4);
TASK_PP(16'hB317,4);
TASK_PP(16'hB318,4);
TASK_PP(16'hB319,4);
TASK_PP(16'hB31A,4);
TASK_PP(16'hB31B,4);
TASK_PP(16'hB31C,4);
TASK_PP(16'hB31D,4);
TASK_PP(16'hB31E,4);
TASK_PP(16'hB31F,4);
TASK_PP(16'hB320,4);
TASK_PP(16'hB321,4);
TASK_PP(16'hB322,4);
TASK_PP(16'hB323,4);
TASK_PP(16'hB324,4);
TASK_PP(16'hB325,4);
TASK_PP(16'hB326,4);
TASK_PP(16'hB327,4);
TASK_PP(16'hB328,4);
TASK_PP(16'hB329,4);
TASK_PP(16'hB32A,4);
TASK_PP(16'hB32B,4);
TASK_PP(16'hB32C,4);
TASK_PP(16'hB32D,4);
TASK_PP(16'hB32E,4);
TASK_PP(16'hB32F,4);
TASK_PP(16'hB330,4);
TASK_PP(16'hB331,4);
TASK_PP(16'hB332,4);
TASK_PP(16'hB333,4);
TASK_PP(16'hB334,4);
TASK_PP(16'hB335,4);
TASK_PP(16'hB336,4);
TASK_PP(16'hB337,4);
TASK_PP(16'hB338,4);
TASK_PP(16'hB339,4);
TASK_PP(16'hB33A,4);
TASK_PP(16'hB33B,4);
TASK_PP(16'hB33C,4);
TASK_PP(16'hB33D,4);
TASK_PP(16'hB33E,4);
TASK_PP(16'hB33F,4);
TASK_PP(16'hB340,4);
TASK_PP(16'hB341,4);
TASK_PP(16'hB342,4);
TASK_PP(16'hB343,4);
TASK_PP(16'hB344,4);
TASK_PP(16'hB345,4);
TASK_PP(16'hB346,4);
TASK_PP(16'hB347,4);
TASK_PP(16'hB348,4);
TASK_PP(16'hB349,4);
TASK_PP(16'hB34A,4);
TASK_PP(16'hB34B,4);
TASK_PP(16'hB34C,4);
TASK_PP(16'hB34D,4);
TASK_PP(16'hB34E,4);
TASK_PP(16'hB34F,4);
TASK_PP(16'hB350,4);
TASK_PP(16'hB351,4);
TASK_PP(16'hB352,4);
TASK_PP(16'hB353,4);
TASK_PP(16'hB354,4);
TASK_PP(16'hB355,4);
TASK_PP(16'hB356,4);
TASK_PP(16'hB357,4);
TASK_PP(16'hB358,4);
TASK_PP(16'hB359,4);
TASK_PP(16'hB35A,4);
TASK_PP(16'hB35B,4);
TASK_PP(16'hB35C,4);
TASK_PP(16'hB35D,4);
TASK_PP(16'hB35E,4);
TASK_PP(16'hB35F,4);
TASK_PP(16'hB360,4);
TASK_PP(16'hB361,4);
TASK_PP(16'hB362,4);
TASK_PP(16'hB363,4);
TASK_PP(16'hB364,4);
TASK_PP(16'hB365,4);
TASK_PP(16'hB366,4);
TASK_PP(16'hB367,4);
TASK_PP(16'hB368,4);
TASK_PP(16'hB369,4);
TASK_PP(16'hB36A,4);
TASK_PP(16'hB36B,4);
TASK_PP(16'hB36C,4);
TASK_PP(16'hB36D,4);
TASK_PP(16'hB36E,4);
TASK_PP(16'hB36F,4);
TASK_PP(16'hB370,4);
TASK_PP(16'hB371,4);
TASK_PP(16'hB372,4);
TASK_PP(16'hB373,4);
TASK_PP(16'hB374,4);
TASK_PP(16'hB375,4);
TASK_PP(16'hB376,4);
TASK_PP(16'hB377,4);
TASK_PP(16'hB378,4);
TASK_PP(16'hB379,4);
TASK_PP(16'hB37A,4);
TASK_PP(16'hB37B,4);
TASK_PP(16'hB37C,4);
TASK_PP(16'hB37D,4);
TASK_PP(16'hB37E,4);
TASK_PP(16'hB37F,4);
TASK_PP(16'hB380,4);
TASK_PP(16'hB381,4);
TASK_PP(16'hB382,4);
TASK_PP(16'hB383,4);
TASK_PP(16'hB384,4);
TASK_PP(16'hB385,4);
TASK_PP(16'hB386,4);
TASK_PP(16'hB387,4);
TASK_PP(16'hB388,4);
TASK_PP(16'hB389,4);
TASK_PP(16'hB38A,4);
TASK_PP(16'hB38B,4);
TASK_PP(16'hB38C,4);
TASK_PP(16'hB38D,4);
TASK_PP(16'hB38E,4);
TASK_PP(16'hB38F,4);
TASK_PP(16'hB390,4);
TASK_PP(16'hB391,4);
TASK_PP(16'hB392,4);
TASK_PP(16'hB393,4);
TASK_PP(16'hB394,4);
TASK_PP(16'hB395,4);
TASK_PP(16'hB396,4);
TASK_PP(16'hB397,4);
TASK_PP(16'hB398,4);
TASK_PP(16'hB399,4);
TASK_PP(16'hB39A,4);
TASK_PP(16'hB39B,4);
TASK_PP(16'hB39C,4);
TASK_PP(16'hB39D,4);
TASK_PP(16'hB39E,4);
TASK_PP(16'hB39F,4);
TASK_PP(16'hB3A0,4);
TASK_PP(16'hB3A1,4);
TASK_PP(16'hB3A2,4);
TASK_PP(16'hB3A3,4);
TASK_PP(16'hB3A4,4);
TASK_PP(16'hB3A5,4);
TASK_PP(16'hB3A6,4);
TASK_PP(16'hB3A7,4);
TASK_PP(16'hB3A8,4);
TASK_PP(16'hB3A9,4);
TASK_PP(16'hB3AA,4);
TASK_PP(16'hB3AB,4);
TASK_PP(16'hB3AC,4);
TASK_PP(16'hB3AD,4);
TASK_PP(16'hB3AE,4);
TASK_PP(16'hB3AF,4);
TASK_PP(16'hB3B0,4);
TASK_PP(16'hB3B1,4);
TASK_PP(16'hB3B2,4);
TASK_PP(16'hB3B3,4);
TASK_PP(16'hB3B4,4);
TASK_PP(16'hB3B5,4);
TASK_PP(16'hB3B6,4);
TASK_PP(16'hB3B7,4);
TASK_PP(16'hB3B8,4);
TASK_PP(16'hB3B9,4);
TASK_PP(16'hB3BA,4);
TASK_PP(16'hB3BB,4);
TASK_PP(16'hB3BC,4);
TASK_PP(16'hB3BD,4);
TASK_PP(16'hB3BE,4);
TASK_PP(16'hB3BF,4);
TASK_PP(16'hB3C0,4);
TASK_PP(16'hB3C1,4);
TASK_PP(16'hB3C2,4);
TASK_PP(16'hB3C3,4);
TASK_PP(16'hB3C4,4);
TASK_PP(16'hB3C5,4);
TASK_PP(16'hB3C6,4);
TASK_PP(16'hB3C7,4);
TASK_PP(16'hB3C8,4);
TASK_PP(16'hB3C9,4);
TASK_PP(16'hB3CA,4);
TASK_PP(16'hB3CB,4);
TASK_PP(16'hB3CC,4);
TASK_PP(16'hB3CD,4);
TASK_PP(16'hB3CE,4);
TASK_PP(16'hB3CF,4);
TASK_PP(16'hB3D0,4);
TASK_PP(16'hB3D1,4);
TASK_PP(16'hB3D2,4);
TASK_PP(16'hB3D3,4);
TASK_PP(16'hB3D4,4);
TASK_PP(16'hB3D5,4);
TASK_PP(16'hB3D6,4);
TASK_PP(16'hB3D7,4);
TASK_PP(16'hB3D8,4);
TASK_PP(16'hB3D9,4);
TASK_PP(16'hB3DA,4);
TASK_PP(16'hB3DB,4);
TASK_PP(16'hB3DC,4);
TASK_PP(16'hB3DD,4);
TASK_PP(16'hB3DE,4);
TASK_PP(16'hB3DF,4);
TASK_PP(16'hB3E0,4);
TASK_PP(16'hB3E1,4);
TASK_PP(16'hB3E2,4);
TASK_PP(16'hB3E3,4);
TASK_PP(16'hB3E4,4);
TASK_PP(16'hB3E5,4);
TASK_PP(16'hB3E6,4);
TASK_PP(16'hB3E7,4);
TASK_PP(16'hB3E8,4);
TASK_PP(16'hB3E9,4);
TASK_PP(16'hB3EA,4);
TASK_PP(16'hB3EB,4);
TASK_PP(16'hB3EC,4);
TASK_PP(16'hB3ED,4);
TASK_PP(16'hB3EE,4);
TASK_PP(16'hB3EF,4);
TASK_PP(16'hB3F0,4);
TASK_PP(16'hB3F1,4);
TASK_PP(16'hB3F2,4);
TASK_PP(16'hB3F3,4);
TASK_PP(16'hB3F4,4);
TASK_PP(16'hB3F5,4);
TASK_PP(16'hB3F6,4);
TASK_PP(16'hB3F7,4);
TASK_PP(16'hB3F8,4);
TASK_PP(16'hB3F9,4);
TASK_PP(16'hB3FA,4);
TASK_PP(16'hB3FB,4);
TASK_PP(16'hB3FC,4);
TASK_PP(16'hB3FD,4);
TASK_PP(16'hB3FE,4);
TASK_PP(16'hB3FF,4);
TASK_PP(16'hB400,4);
TASK_PP(16'hB401,4);
TASK_PP(16'hB402,4);
TASK_PP(16'hB403,4);
TASK_PP(16'hB404,4);
TASK_PP(16'hB405,4);
TASK_PP(16'hB406,4);
TASK_PP(16'hB407,4);
TASK_PP(16'hB408,4);
TASK_PP(16'hB409,4);
TASK_PP(16'hB40A,4);
TASK_PP(16'hB40B,4);
TASK_PP(16'hB40C,4);
TASK_PP(16'hB40D,4);
TASK_PP(16'hB40E,4);
TASK_PP(16'hB40F,4);
TASK_PP(16'hB410,4);
TASK_PP(16'hB411,4);
TASK_PP(16'hB412,4);
TASK_PP(16'hB413,4);
TASK_PP(16'hB414,4);
TASK_PP(16'hB415,4);
TASK_PP(16'hB416,4);
TASK_PP(16'hB417,4);
TASK_PP(16'hB418,4);
TASK_PP(16'hB419,4);
TASK_PP(16'hB41A,4);
TASK_PP(16'hB41B,4);
TASK_PP(16'hB41C,4);
TASK_PP(16'hB41D,4);
TASK_PP(16'hB41E,4);
TASK_PP(16'hB41F,4);
TASK_PP(16'hB420,4);
TASK_PP(16'hB421,4);
TASK_PP(16'hB422,4);
TASK_PP(16'hB423,4);
TASK_PP(16'hB424,4);
TASK_PP(16'hB425,4);
TASK_PP(16'hB426,4);
TASK_PP(16'hB427,4);
TASK_PP(16'hB428,4);
TASK_PP(16'hB429,4);
TASK_PP(16'hB42A,4);
TASK_PP(16'hB42B,4);
TASK_PP(16'hB42C,4);
TASK_PP(16'hB42D,4);
TASK_PP(16'hB42E,4);
TASK_PP(16'hB42F,4);
TASK_PP(16'hB430,4);
TASK_PP(16'hB431,4);
TASK_PP(16'hB432,4);
TASK_PP(16'hB433,4);
TASK_PP(16'hB434,4);
TASK_PP(16'hB435,4);
TASK_PP(16'hB436,4);
TASK_PP(16'hB437,4);
TASK_PP(16'hB438,4);
TASK_PP(16'hB439,4);
TASK_PP(16'hB43A,4);
TASK_PP(16'hB43B,4);
TASK_PP(16'hB43C,4);
TASK_PP(16'hB43D,4);
TASK_PP(16'hB43E,4);
TASK_PP(16'hB43F,4);
TASK_PP(16'hB440,4);
TASK_PP(16'hB441,4);
TASK_PP(16'hB442,4);
TASK_PP(16'hB443,4);
TASK_PP(16'hB444,4);
TASK_PP(16'hB445,4);
TASK_PP(16'hB446,4);
TASK_PP(16'hB447,4);
TASK_PP(16'hB448,4);
TASK_PP(16'hB449,4);
TASK_PP(16'hB44A,4);
TASK_PP(16'hB44B,4);
TASK_PP(16'hB44C,4);
TASK_PP(16'hB44D,4);
TASK_PP(16'hB44E,4);
TASK_PP(16'hB44F,4);
TASK_PP(16'hB450,4);
TASK_PP(16'hB451,4);
TASK_PP(16'hB452,4);
TASK_PP(16'hB453,4);
TASK_PP(16'hB454,4);
TASK_PP(16'hB455,4);
TASK_PP(16'hB456,4);
TASK_PP(16'hB457,4);
TASK_PP(16'hB458,4);
TASK_PP(16'hB459,4);
TASK_PP(16'hB45A,4);
TASK_PP(16'hB45B,4);
TASK_PP(16'hB45C,4);
TASK_PP(16'hB45D,4);
TASK_PP(16'hB45E,4);
TASK_PP(16'hB45F,4);
TASK_PP(16'hB460,4);
TASK_PP(16'hB461,4);
TASK_PP(16'hB462,4);
TASK_PP(16'hB463,4);
TASK_PP(16'hB464,4);
TASK_PP(16'hB465,4);
TASK_PP(16'hB466,4);
TASK_PP(16'hB467,4);
TASK_PP(16'hB468,4);
TASK_PP(16'hB469,4);
TASK_PP(16'hB46A,4);
TASK_PP(16'hB46B,4);
TASK_PP(16'hB46C,4);
TASK_PP(16'hB46D,4);
TASK_PP(16'hB46E,4);
TASK_PP(16'hB46F,4);
TASK_PP(16'hB470,4);
TASK_PP(16'hB471,4);
TASK_PP(16'hB472,4);
TASK_PP(16'hB473,4);
TASK_PP(16'hB474,4);
TASK_PP(16'hB475,4);
TASK_PP(16'hB476,4);
TASK_PP(16'hB477,4);
TASK_PP(16'hB478,4);
TASK_PP(16'hB479,4);
TASK_PP(16'hB47A,4);
TASK_PP(16'hB47B,4);
TASK_PP(16'hB47C,4);
TASK_PP(16'hB47D,4);
TASK_PP(16'hB47E,4);
TASK_PP(16'hB47F,4);
TASK_PP(16'hB480,4);
TASK_PP(16'hB481,4);
TASK_PP(16'hB482,4);
TASK_PP(16'hB483,4);
TASK_PP(16'hB484,4);
TASK_PP(16'hB485,4);
TASK_PP(16'hB486,4);
TASK_PP(16'hB487,4);
TASK_PP(16'hB488,4);
TASK_PP(16'hB489,4);
TASK_PP(16'hB48A,4);
TASK_PP(16'hB48B,4);
TASK_PP(16'hB48C,4);
TASK_PP(16'hB48D,4);
TASK_PP(16'hB48E,4);
TASK_PP(16'hB48F,4);
TASK_PP(16'hB490,4);
TASK_PP(16'hB491,4);
TASK_PP(16'hB492,4);
TASK_PP(16'hB493,4);
TASK_PP(16'hB494,4);
TASK_PP(16'hB495,4);
TASK_PP(16'hB496,4);
TASK_PP(16'hB497,4);
TASK_PP(16'hB498,4);
TASK_PP(16'hB499,4);
TASK_PP(16'hB49A,4);
TASK_PP(16'hB49B,4);
TASK_PP(16'hB49C,4);
TASK_PP(16'hB49D,4);
TASK_PP(16'hB49E,4);
TASK_PP(16'hB49F,4);
TASK_PP(16'hB4A0,4);
TASK_PP(16'hB4A1,4);
TASK_PP(16'hB4A2,4);
TASK_PP(16'hB4A3,4);
TASK_PP(16'hB4A4,4);
TASK_PP(16'hB4A5,4);
TASK_PP(16'hB4A6,4);
TASK_PP(16'hB4A7,4);
TASK_PP(16'hB4A8,4);
TASK_PP(16'hB4A9,4);
TASK_PP(16'hB4AA,4);
TASK_PP(16'hB4AB,4);
TASK_PP(16'hB4AC,4);
TASK_PP(16'hB4AD,4);
TASK_PP(16'hB4AE,4);
TASK_PP(16'hB4AF,4);
TASK_PP(16'hB4B0,4);
TASK_PP(16'hB4B1,4);
TASK_PP(16'hB4B2,4);
TASK_PP(16'hB4B3,4);
TASK_PP(16'hB4B4,4);
TASK_PP(16'hB4B5,4);
TASK_PP(16'hB4B6,4);
TASK_PP(16'hB4B7,4);
TASK_PP(16'hB4B8,4);
TASK_PP(16'hB4B9,4);
TASK_PP(16'hB4BA,4);
TASK_PP(16'hB4BB,4);
TASK_PP(16'hB4BC,4);
TASK_PP(16'hB4BD,4);
TASK_PP(16'hB4BE,4);
TASK_PP(16'hB4BF,4);
TASK_PP(16'hB4C0,4);
TASK_PP(16'hB4C1,4);
TASK_PP(16'hB4C2,4);
TASK_PP(16'hB4C3,4);
TASK_PP(16'hB4C4,4);
TASK_PP(16'hB4C5,4);
TASK_PP(16'hB4C6,4);
TASK_PP(16'hB4C7,4);
TASK_PP(16'hB4C8,4);
TASK_PP(16'hB4C9,4);
TASK_PP(16'hB4CA,4);
TASK_PP(16'hB4CB,4);
TASK_PP(16'hB4CC,4);
TASK_PP(16'hB4CD,4);
TASK_PP(16'hB4CE,4);
TASK_PP(16'hB4CF,4);
TASK_PP(16'hB4D0,4);
TASK_PP(16'hB4D1,4);
TASK_PP(16'hB4D2,4);
TASK_PP(16'hB4D3,4);
TASK_PP(16'hB4D4,4);
TASK_PP(16'hB4D5,4);
TASK_PP(16'hB4D6,4);
TASK_PP(16'hB4D7,4);
TASK_PP(16'hB4D8,4);
TASK_PP(16'hB4D9,4);
TASK_PP(16'hB4DA,4);
TASK_PP(16'hB4DB,4);
TASK_PP(16'hB4DC,4);
TASK_PP(16'hB4DD,4);
TASK_PP(16'hB4DE,4);
TASK_PP(16'hB4DF,4);
TASK_PP(16'hB4E0,4);
TASK_PP(16'hB4E1,4);
TASK_PP(16'hB4E2,4);
TASK_PP(16'hB4E3,4);
TASK_PP(16'hB4E4,4);
TASK_PP(16'hB4E5,4);
TASK_PP(16'hB4E6,4);
TASK_PP(16'hB4E7,4);
TASK_PP(16'hB4E8,4);
TASK_PP(16'hB4E9,4);
TASK_PP(16'hB4EA,4);
TASK_PP(16'hB4EB,4);
TASK_PP(16'hB4EC,4);
TASK_PP(16'hB4ED,4);
TASK_PP(16'hB4EE,4);
TASK_PP(16'hB4EF,4);
TASK_PP(16'hB4F0,4);
TASK_PP(16'hB4F1,4);
TASK_PP(16'hB4F2,4);
TASK_PP(16'hB4F3,4);
TASK_PP(16'hB4F4,4);
TASK_PP(16'hB4F5,4);
TASK_PP(16'hB4F6,4);
TASK_PP(16'hB4F7,4);
TASK_PP(16'hB4F8,4);
TASK_PP(16'hB4F9,4);
TASK_PP(16'hB4FA,4);
TASK_PP(16'hB4FB,4);
TASK_PP(16'hB4FC,4);
TASK_PP(16'hB4FD,4);
TASK_PP(16'hB4FE,4);
TASK_PP(16'hB4FF,4);
TASK_PP(16'hB500,4);
TASK_PP(16'hB501,4);
TASK_PP(16'hB502,4);
TASK_PP(16'hB503,4);
TASK_PP(16'hB504,4);
TASK_PP(16'hB505,4);
TASK_PP(16'hB506,4);
TASK_PP(16'hB507,4);
TASK_PP(16'hB508,4);
TASK_PP(16'hB509,4);
TASK_PP(16'hB50A,4);
TASK_PP(16'hB50B,4);
TASK_PP(16'hB50C,4);
TASK_PP(16'hB50D,4);
TASK_PP(16'hB50E,4);
TASK_PP(16'hB50F,4);
TASK_PP(16'hB510,4);
TASK_PP(16'hB511,4);
TASK_PP(16'hB512,4);
TASK_PP(16'hB513,4);
TASK_PP(16'hB514,4);
TASK_PP(16'hB515,4);
TASK_PP(16'hB516,4);
TASK_PP(16'hB517,4);
TASK_PP(16'hB518,4);
TASK_PP(16'hB519,4);
TASK_PP(16'hB51A,4);
TASK_PP(16'hB51B,4);
TASK_PP(16'hB51C,4);
TASK_PP(16'hB51D,4);
TASK_PP(16'hB51E,4);
TASK_PP(16'hB51F,4);
TASK_PP(16'hB520,4);
TASK_PP(16'hB521,4);
TASK_PP(16'hB522,4);
TASK_PP(16'hB523,4);
TASK_PP(16'hB524,4);
TASK_PP(16'hB525,4);
TASK_PP(16'hB526,4);
TASK_PP(16'hB527,4);
TASK_PP(16'hB528,4);
TASK_PP(16'hB529,4);
TASK_PP(16'hB52A,4);
TASK_PP(16'hB52B,4);
TASK_PP(16'hB52C,4);
TASK_PP(16'hB52D,4);
TASK_PP(16'hB52E,4);
TASK_PP(16'hB52F,4);
TASK_PP(16'hB530,4);
TASK_PP(16'hB531,4);
TASK_PP(16'hB532,4);
TASK_PP(16'hB533,4);
TASK_PP(16'hB534,4);
TASK_PP(16'hB535,4);
TASK_PP(16'hB536,4);
TASK_PP(16'hB537,4);
TASK_PP(16'hB538,4);
TASK_PP(16'hB539,4);
TASK_PP(16'hB53A,4);
TASK_PP(16'hB53B,4);
TASK_PP(16'hB53C,4);
TASK_PP(16'hB53D,4);
TASK_PP(16'hB53E,4);
TASK_PP(16'hB53F,4);
TASK_PP(16'hB540,4);
TASK_PP(16'hB541,4);
TASK_PP(16'hB542,4);
TASK_PP(16'hB543,4);
TASK_PP(16'hB544,4);
TASK_PP(16'hB545,4);
TASK_PP(16'hB546,4);
TASK_PP(16'hB547,4);
TASK_PP(16'hB548,4);
TASK_PP(16'hB549,4);
TASK_PP(16'hB54A,4);
TASK_PP(16'hB54B,4);
TASK_PP(16'hB54C,4);
TASK_PP(16'hB54D,4);
TASK_PP(16'hB54E,4);
TASK_PP(16'hB54F,4);
TASK_PP(16'hB550,4);
TASK_PP(16'hB551,4);
TASK_PP(16'hB552,4);
TASK_PP(16'hB553,4);
TASK_PP(16'hB554,4);
TASK_PP(16'hB555,4);
TASK_PP(16'hB556,4);
TASK_PP(16'hB557,4);
TASK_PP(16'hB558,4);
TASK_PP(16'hB559,4);
TASK_PP(16'hB55A,4);
TASK_PP(16'hB55B,4);
TASK_PP(16'hB55C,4);
TASK_PP(16'hB55D,4);
TASK_PP(16'hB55E,4);
TASK_PP(16'hB55F,4);
TASK_PP(16'hB560,4);
TASK_PP(16'hB561,4);
TASK_PP(16'hB562,4);
TASK_PP(16'hB563,4);
TASK_PP(16'hB564,4);
TASK_PP(16'hB565,4);
TASK_PP(16'hB566,4);
TASK_PP(16'hB567,4);
TASK_PP(16'hB568,4);
TASK_PP(16'hB569,4);
TASK_PP(16'hB56A,4);
TASK_PP(16'hB56B,4);
TASK_PP(16'hB56C,4);
TASK_PP(16'hB56D,4);
TASK_PP(16'hB56E,4);
TASK_PP(16'hB56F,4);
TASK_PP(16'hB570,4);
TASK_PP(16'hB571,4);
TASK_PP(16'hB572,4);
TASK_PP(16'hB573,4);
TASK_PP(16'hB574,4);
TASK_PP(16'hB575,4);
TASK_PP(16'hB576,4);
TASK_PP(16'hB577,4);
TASK_PP(16'hB578,4);
TASK_PP(16'hB579,4);
TASK_PP(16'hB57A,4);
TASK_PP(16'hB57B,4);
TASK_PP(16'hB57C,4);
TASK_PP(16'hB57D,4);
TASK_PP(16'hB57E,4);
TASK_PP(16'hB57F,4);
TASK_PP(16'hB580,4);
TASK_PP(16'hB581,4);
TASK_PP(16'hB582,4);
TASK_PP(16'hB583,4);
TASK_PP(16'hB584,4);
TASK_PP(16'hB585,4);
TASK_PP(16'hB586,4);
TASK_PP(16'hB587,4);
TASK_PP(16'hB588,4);
TASK_PP(16'hB589,4);
TASK_PP(16'hB58A,4);
TASK_PP(16'hB58B,4);
TASK_PP(16'hB58C,4);
TASK_PP(16'hB58D,4);
TASK_PP(16'hB58E,4);
TASK_PP(16'hB58F,4);
TASK_PP(16'hB590,4);
TASK_PP(16'hB591,4);
TASK_PP(16'hB592,4);
TASK_PP(16'hB593,4);
TASK_PP(16'hB594,4);
TASK_PP(16'hB595,4);
TASK_PP(16'hB596,4);
TASK_PP(16'hB597,4);
TASK_PP(16'hB598,4);
TASK_PP(16'hB599,4);
TASK_PP(16'hB59A,4);
TASK_PP(16'hB59B,4);
TASK_PP(16'hB59C,4);
TASK_PP(16'hB59D,4);
TASK_PP(16'hB59E,4);
TASK_PP(16'hB59F,4);
TASK_PP(16'hB5A0,4);
TASK_PP(16'hB5A1,4);
TASK_PP(16'hB5A2,4);
TASK_PP(16'hB5A3,4);
TASK_PP(16'hB5A4,4);
TASK_PP(16'hB5A5,4);
TASK_PP(16'hB5A6,4);
TASK_PP(16'hB5A7,4);
TASK_PP(16'hB5A8,4);
TASK_PP(16'hB5A9,4);
TASK_PP(16'hB5AA,4);
TASK_PP(16'hB5AB,4);
TASK_PP(16'hB5AC,4);
TASK_PP(16'hB5AD,4);
TASK_PP(16'hB5AE,4);
TASK_PP(16'hB5AF,4);
TASK_PP(16'hB5B0,4);
TASK_PP(16'hB5B1,4);
TASK_PP(16'hB5B2,4);
TASK_PP(16'hB5B3,4);
TASK_PP(16'hB5B4,4);
TASK_PP(16'hB5B5,4);
TASK_PP(16'hB5B6,4);
TASK_PP(16'hB5B7,4);
TASK_PP(16'hB5B8,4);
TASK_PP(16'hB5B9,4);
TASK_PP(16'hB5BA,4);
TASK_PP(16'hB5BB,4);
TASK_PP(16'hB5BC,4);
TASK_PP(16'hB5BD,4);
TASK_PP(16'hB5BE,4);
TASK_PP(16'hB5BF,4);
TASK_PP(16'hB5C0,4);
TASK_PP(16'hB5C1,4);
TASK_PP(16'hB5C2,4);
TASK_PP(16'hB5C3,4);
TASK_PP(16'hB5C4,4);
TASK_PP(16'hB5C5,4);
TASK_PP(16'hB5C6,4);
TASK_PP(16'hB5C7,4);
TASK_PP(16'hB5C8,4);
TASK_PP(16'hB5C9,4);
TASK_PP(16'hB5CA,4);
TASK_PP(16'hB5CB,4);
TASK_PP(16'hB5CC,4);
TASK_PP(16'hB5CD,4);
TASK_PP(16'hB5CE,4);
TASK_PP(16'hB5CF,4);
TASK_PP(16'hB5D0,4);
TASK_PP(16'hB5D1,4);
TASK_PP(16'hB5D2,4);
TASK_PP(16'hB5D3,4);
TASK_PP(16'hB5D4,4);
TASK_PP(16'hB5D5,4);
TASK_PP(16'hB5D6,4);
TASK_PP(16'hB5D7,4);
TASK_PP(16'hB5D8,4);
TASK_PP(16'hB5D9,4);
TASK_PP(16'hB5DA,4);
TASK_PP(16'hB5DB,4);
TASK_PP(16'hB5DC,4);
TASK_PP(16'hB5DD,4);
TASK_PP(16'hB5DE,4);
TASK_PP(16'hB5DF,4);
TASK_PP(16'hB5E0,4);
TASK_PP(16'hB5E1,4);
TASK_PP(16'hB5E2,4);
TASK_PP(16'hB5E3,4);
TASK_PP(16'hB5E4,4);
TASK_PP(16'hB5E5,4);
TASK_PP(16'hB5E6,4);
TASK_PP(16'hB5E7,4);
TASK_PP(16'hB5E8,4);
TASK_PP(16'hB5E9,4);
TASK_PP(16'hB5EA,4);
TASK_PP(16'hB5EB,4);
TASK_PP(16'hB5EC,4);
TASK_PP(16'hB5ED,4);
TASK_PP(16'hB5EE,4);
TASK_PP(16'hB5EF,4);
TASK_PP(16'hB5F0,4);
TASK_PP(16'hB5F1,4);
TASK_PP(16'hB5F2,4);
TASK_PP(16'hB5F3,4);
TASK_PP(16'hB5F4,4);
TASK_PP(16'hB5F5,4);
TASK_PP(16'hB5F6,4);
TASK_PP(16'hB5F7,4);
TASK_PP(16'hB5F8,4);
TASK_PP(16'hB5F9,4);
TASK_PP(16'hB5FA,4);
TASK_PP(16'hB5FB,4);
TASK_PP(16'hB5FC,4);
TASK_PP(16'hB5FD,4);
TASK_PP(16'hB5FE,4);
TASK_PP(16'hB5FF,4);
TASK_PP(16'hB600,4);
TASK_PP(16'hB601,4);
TASK_PP(16'hB602,4);
TASK_PP(16'hB603,4);
TASK_PP(16'hB604,4);
TASK_PP(16'hB605,4);
TASK_PP(16'hB606,4);
TASK_PP(16'hB607,4);
TASK_PP(16'hB608,4);
TASK_PP(16'hB609,4);
TASK_PP(16'hB60A,4);
TASK_PP(16'hB60B,4);
TASK_PP(16'hB60C,4);
TASK_PP(16'hB60D,4);
TASK_PP(16'hB60E,4);
TASK_PP(16'hB60F,4);
TASK_PP(16'hB610,4);
TASK_PP(16'hB611,4);
TASK_PP(16'hB612,4);
TASK_PP(16'hB613,4);
TASK_PP(16'hB614,4);
TASK_PP(16'hB615,4);
TASK_PP(16'hB616,4);
TASK_PP(16'hB617,4);
TASK_PP(16'hB618,4);
TASK_PP(16'hB619,4);
TASK_PP(16'hB61A,4);
TASK_PP(16'hB61B,4);
TASK_PP(16'hB61C,4);
TASK_PP(16'hB61D,4);
TASK_PP(16'hB61E,4);
TASK_PP(16'hB61F,4);
TASK_PP(16'hB620,4);
TASK_PP(16'hB621,4);
TASK_PP(16'hB622,4);
TASK_PP(16'hB623,4);
TASK_PP(16'hB624,4);
TASK_PP(16'hB625,4);
TASK_PP(16'hB626,4);
TASK_PP(16'hB627,4);
TASK_PP(16'hB628,4);
TASK_PP(16'hB629,4);
TASK_PP(16'hB62A,4);
TASK_PP(16'hB62B,4);
TASK_PP(16'hB62C,4);
TASK_PP(16'hB62D,4);
TASK_PP(16'hB62E,4);
TASK_PP(16'hB62F,4);
TASK_PP(16'hB630,4);
TASK_PP(16'hB631,4);
TASK_PP(16'hB632,4);
TASK_PP(16'hB633,4);
TASK_PP(16'hB634,4);
TASK_PP(16'hB635,4);
TASK_PP(16'hB636,4);
TASK_PP(16'hB637,4);
TASK_PP(16'hB638,4);
TASK_PP(16'hB639,4);
TASK_PP(16'hB63A,4);
TASK_PP(16'hB63B,4);
TASK_PP(16'hB63C,4);
TASK_PP(16'hB63D,4);
TASK_PP(16'hB63E,4);
TASK_PP(16'hB63F,4);
TASK_PP(16'hB640,4);
TASK_PP(16'hB641,4);
TASK_PP(16'hB642,4);
TASK_PP(16'hB643,4);
TASK_PP(16'hB644,4);
TASK_PP(16'hB645,4);
TASK_PP(16'hB646,4);
TASK_PP(16'hB647,4);
TASK_PP(16'hB648,4);
TASK_PP(16'hB649,4);
TASK_PP(16'hB64A,4);
TASK_PP(16'hB64B,4);
TASK_PP(16'hB64C,4);
TASK_PP(16'hB64D,4);
TASK_PP(16'hB64E,4);
TASK_PP(16'hB64F,4);
TASK_PP(16'hB650,4);
TASK_PP(16'hB651,4);
TASK_PP(16'hB652,4);
TASK_PP(16'hB653,4);
TASK_PP(16'hB654,4);
TASK_PP(16'hB655,4);
TASK_PP(16'hB656,4);
TASK_PP(16'hB657,4);
TASK_PP(16'hB658,4);
TASK_PP(16'hB659,4);
TASK_PP(16'hB65A,4);
TASK_PP(16'hB65B,4);
TASK_PP(16'hB65C,4);
TASK_PP(16'hB65D,4);
TASK_PP(16'hB65E,4);
TASK_PP(16'hB65F,4);
TASK_PP(16'hB660,4);
TASK_PP(16'hB661,4);
TASK_PP(16'hB662,4);
TASK_PP(16'hB663,4);
TASK_PP(16'hB664,4);
TASK_PP(16'hB665,4);
TASK_PP(16'hB666,4);
TASK_PP(16'hB667,4);
TASK_PP(16'hB668,4);
TASK_PP(16'hB669,4);
TASK_PP(16'hB66A,4);
TASK_PP(16'hB66B,4);
TASK_PP(16'hB66C,4);
TASK_PP(16'hB66D,4);
TASK_PP(16'hB66E,4);
TASK_PP(16'hB66F,4);
TASK_PP(16'hB670,4);
TASK_PP(16'hB671,4);
TASK_PP(16'hB672,4);
TASK_PP(16'hB673,4);
TASK_PP(16'hB674,4);
TASK_PP(16'hB675,4);
TASK_PP(16'hB676,4);
TASK_PP(16'hB677,4);
TASK_PP(16'hB678,4);
TASK_PP(16'hB679,4);
TASK_PP(16'hB67A,4);
TASK_PP(16'hB67B,4);
TASK_PP(16'hB67C,4);
TASK_PP(16'hB67D,4);
TASK_PP(16'hB67E,4);
TASK_PP(16'hB67F,4);
TASK_PP(16'hB680,4);
TASK_PP(16'hB681,4);
TASK_PP(16'hB682,4);
TASK_PP(16'hB683,4);
TASK_PP(16'hB684,4);
TASK_PP(16'hB685,4);
TASK_PP(16'hB686,4);
TASK_PP(16'hB687,4);
TASK_PP(16'hB688,4);
TASK_PP(16'hB689,4);
TASK_PP(16'hB68A,4);
TASK_PP(16'hB68B,4);
TASK_PP(16'hB68C,4);
TASK_PP(16'hB68D,4);
TASK_PP(16'hB68E,4);
TASK_PP(16'hB68F,4);
TASK_PP(16'hB690,4);
TASK_PP(16'hB691,4);
TASK_PP(16'hB692,4);
TASK_PP(16'hB693,4);
TASK_PP(16'hB694,4);
TASK_PP(16'hB695,4);
TASK_PP(16'hB696,4);
TASK_PP(16'hB697,4);
TASK_PP(16'hB698,4);
TASK_PP(16'hB699,4);
TASK_PP(16'hB69A,4);
TASK_PP(16'hB69B,4);
TASK_PP(16'hB69C,4);
TASK_PP(16'hB69D,4);
TASK_PP(16'hB69E,4);
TASK_PP(16'hB69F,4);
TASK_PP(16'hB6A0,4);
TASK_PP(16'hB6A1,4);
TASK_PP(16'hB6A2,4);
TASK_PP(16'hB6A3,4);
TASK_PP(16'hB6A4,4);
TASK_PP(16'hB6A5,4);
TASK_PP(16'hB6A6,4);
TASK_PP(16'hB6A7,4);
TASK_PP(16'hB6A8,4);
TASK_PP(16'hB6A9,4);
TASK_PP(16'hB6AA,4);
TASK_PP(16'hB6AB,4);
TASK_PP(16'hB6AC,4);
TASK_PP(16'hB6AD,4);
TASK_PP(16'hB6AE,4);
TASK_PP(16'hB6AF,4);
TASK_PP(16'hB6B0,4);
TASK_PP(16'hB6B1,4);
TASK_PP(16'hB6B2,4);
TASK_PP(16'hB6B3,4);
TASK_PP(16'hB6B4,4);
TASK_PP(16'hB6B5,4);
TASK_PP(16'hB6B6,4);
TASK_PP(16'hB6B7,4);
TASK_PP(16'hB6B8,4);
TASK_PP(16'hB6B9,4);
TASK_PP(16'hB6BA,4);
TASK_PP(16'hB6BB,4);
TASK_PP(16'hB6BC,4);
TASK_PP(16'hB6BD,4);
TASK_PP(16'hB6BE,4);
TASK_PP(16'hB6BF,4);
TASK_PP(16'hB6C0,4);
TASK_PP(16'hB6C1,4);
TASK_PP(16'hB6C2,4);
TASK_PP(16'hB6C3,4);
TASK_PP(16'hB6C4,4);
TASK_PP(16'hB6C5,4);
TASK_PP(16'hB6C6,4);
TASK_PP(16'hB6C7,4);
TASK_PP(16'hB6C8,4);
TASK_PP(16'hB6C9,4);
TASK_PP(16'hB6CA,4);
TASK_PP(16'hB6CB,4);
TASK_PP(16'hB6CC,4);
TASK_PP(16'hB6CD,4);
TASK_PP(16'hB6CE,4);
TASK_PP(16'hB6CF,4);
TASK_PP(16'hB6D0,4);
TASK_PP(16'hB6D1,4);
TASK_PP(16'hB6D2,4);
TASK_PP(16'hB6D3,4);
TASK_PP(16'hB6D4,4);
TASK_PP(16'hB6D5,4);
TASK_PP(16'hB6D6,4);
TASK_PP(16'hB6D7,4);
TASK_PP(16'hB6D8,4);
TASK_PP(16'hB6D9,4);
TASK_PP(16'hB6DA,4);
TASK_PP(16'hB6DB,4);
TASK_PP(16'hB6DC,4);
TASK_PP(16'hB6DD,4);
TASK_PP(16'hB6DE,4);
TASK_PP(16'hB6DF,4);
TASK_PP(16'hB6E0,4);
TASK_PP(16'hB6E1,4);
TASK_PP(16'hB6E2,4);
TASK_PP(16'hB6E3,4);
TASK_PP(16'hB6E4,4);
TASK_PP(16'hB6E5,4);
TASK_PP(16'hB6E6,4);
TASK_PP(16'hB6E7,4);
TASK_PP(16'hB6E8,4);
TASK_PP(16'hB6E9,4);
TASK_PP(16'hB6EA,4);
TASK_PP(16'hB6EB,4);
TASK_PP(16'hB6EC,4);
TASK_PP(16'hB6ED,4);
TASK_PP(16'hB6EE,4);
TASK_PP(16'hB6EF,4);
TASK_PP(16'hB6F0,4);
TASK_PP(16'hB6F1,4);
TASK_PP(16'hB6F2,4);
TASK_PP(16'hB6F3,4);
TASK_PP(16'hB6F4,4);
TASK_PP(16'hB6F5,4);
TASK_PP(16'hB6F6,4);
TASK_PP(16'hB6F7,4);
TASK_PP(16'hB6F8,4);
TASK_PP(16'hB6F9,4);
TASK_PP(16'hB6FA,4);
TASK_PP(16'hB6FB,4);
TASK_PP(16'hB6FC,4);
TASK_PP(16'hB6FD,4);
TASK_PP(16'hB6FE,4);
TASK_PP(16'hB6FF,4);
TASK_PP(16'hB700,4);
TASK_PP(16'hB701,4);
TASK_PP(16'hB702,4);
TASK_PP(16'hB703,4);
TASK_PP(16'hB704,4);
TASK_PP(16'hB705,4);
TASK_PP(16'hB706,4);
TASK_PP(16'hB707,4);
TASK_PP(16'hB708,4);
TASK_PP(16'hB709,4);
TASK_PP(16'hB70A,4);
TASK_PP(16'hB70B,4);
TASK_PP(16'hB70C,4);
TASK_PP(16'hB70D,4);
TASK_PP(16'hB70E,4);
TASK_PP(16'hB70F,4);
TASK_PP(16'hB710,4);
TASK_PP(16'hB711,4);
TASK_PP(16'hB712,4);
TASK_PP(16'hB713,4);
TASK_PP(16'hB714,4);
TASK_PP(16'hB715,4);
TASK_PP(16'hB716,4);
TASK_PP(16'hB717,4);
TASK_PP(16'hB718,4);
TASK_PP(16'hB719,4);
TASK_PP(16'hB71A,4);
TASK_PP(16'hB71B,4);
TASK_PP(16'hB71C,4);
TASK_PP(16'hB71D,4);
TASK_PP(16'hB71E,4);
TASK_PP(16'hB71F,4);
TASK_PP(16'hB720,4);
TASK_PP(16'hB721,4);
TASK_PP(16'hB722,4);
TASK_PP(16'hB723,4);
TASK_PP(16'hB724,4);
TASK_PP(16'hB725,4);
TASK_PP(16'hB726,4);
TASK_PP(16'hB727,4);
TASK_PP(16'hB728,4);
TASK_PP(16'hB729,4);
TASK_PP(16'hB72A,4);
TASK_PP(16'hB72B,4);
TASK_PP(16'hB72C,4);
TASK_PP(16'hB72D,4);
TASK_PP(16'hB72E,4);
TASK_PP(16'hB72F,4);
TASK_PP(16'hB730,4);
TASK_PP(16'hB731,4);
TASK_PP(16'hB732,4);
TASK_PP(16'hB733,4);
TASK_PP(16'hB734,4);
TASK_PP(16'hB735,4);
TASK_PP(16'hB736,4);
TASK_PP(16'hB737,4);
TASK_PP(16'hB738,4);
TASK_PP(16'hB739,4);
TASK_PP(16'hB73A,4);
TASK_PP(16'hB73B,4);
TASK_PP(16'hB73C,4);
TASK_PP(16'hB73D,4);
TASK_PP(16'hB73E,4);
TASK_PP(16'hB73F,4);
TASK_PP(16'hB740,4);
TASK_PP(16'hB741,4);
TASK_PP(16'hB742,4);
TASK_PP(16'hB743,4);
TASK_PP(16'hB744,4);
TASK_PP(16'hB745,4);
TASK_PP(16'hB746,4);
TASK_PP(16'hB747,4);
TASK_PP(16'hB748,4);
TASK_PP(16'hB749,4);
TASK_PP(16'hB74A,4);
TASK_PP(16'hB74B,4);
TASK_PP(16'hB74C,4);
TASK_PP(16'hB74D,4);
TASK_PP(16'hB74E,4);
TASK_PP(16'hB74F,4);
TASK_PP(16'hB750,4);
TASK_PP(16'hB751,4);
TASK_PP(16'hB752,4);
TASK_PP(16'hB753,4);
TASK_PP(16'hB754,4);
TASK_PP(16'hB755,4);
TASK_PP(16'hB756,4);
TASK_PP(16'hB757,4);
TASK_PP(16'hB758,4);
TASK_PP(16'hB759,4);
TASK_PP(16'hB75A,4);
TASK_PP(16'hB75B,4);
TASK_PP(16'hB75C,4);
TASK_PP(16'hB75D,4);
TASK_PP(16'hB75E,4);
TASK_PP(16'hB75F,4);
TASK_PP(16'hB760,4);
TASK_PP(16'hB761,4);
TASK_PP(16'hB762,4);
TASK_PP(16'hB763,4);
TASK_PP(16'hB764,4);
TASK_PP(16'hB765,4);
TASK_PP(16'hB766,4);
TASK_PP(16'hB767,4);
TASK_PP(16'hB768,4);
TASK_PP(16'hB769,4);
TASK_PP(16'hB76A,4);
TASK_PP(16'hB76B,4);
TASK_PP(16'hB76C,4);
TASK_PP(16'hB76D,4);
TASK_PP(16'hB76E,4);
TASK_PP(16'hB76F,4);
TASK_PP(16'hB770,4);
TASK_PP(16'hB771,4);
TASK_PP(16'hB772,4);
TASK_PP(16'hB773,4);
TASK_PP(16'hB774,4);
TASK_PP(16'hB775,4);
TASK_PP(16'hB776,4);
TASK_PP(16'hB777,4);
TASK_PP(16'hB778,4);
TASK_PP(16'hB779,4);
TASK_PP(16'hB77A,4);
TASK_PP(16'hB77B,4);
TASK_PP(16'hB77C,4);
TASK_PP(16'hB77D,4);
TASK_PP(16'hB77E,4);
TASK_PP(16'hB77F,4);
TASK_PP(16'hB780,4);
TASK_PP(16'hB781,4);
TASK_PP(16'hB782,4);
TASK_PP(16'hB783,4);
TASK_PP(16'hB784,4);
TASK_PP(16'hB785,4);
TASK_PP(16'hB786,4);
TASK_PP(16'hB787,4);
TASK_PP(16'hB788,4);
TASK_PP(16'hB789,4);
TASK_PP(16'hB78A,4);
TASK_PP(16'hB78B,4);
TASK_PP(16'hB78C,4);
TASK_PP(16'hB78D,4);
TASK_PP(16'hB78E,4);
TASK_PP(16'hB78F,4);
TASK_PP(16'hB790,4);
TASK_PP(16'hB791,4);
TASK_PP(16'hB792,4);
TASK_PP(16'hB793,4);
TASK_PP(16'hB794,4);
TASK_PP(16'hB795,4);
TASK_PP(16'hB796,4);
TASK_PP(16'hB797,4);
TASK_PP(16'hB798,4);
TASK_PP(16'hB799,4);
TASK_PP(16'hB79A,4);
TASK_PP(16'hB79B,4);
TASK_PP(16'hB79C,4);
TASK_PP(16'hB79D,4);
TASK_PP(16'hB79E,4);
TASK_PP(16'hB79F,4);
TASK_PP(16'hB7A0,4);
TASK_PP(16'hB7A1,4);
TASK_PP(16'hB7A2,4);
TASK_PP(16'hB7A3,4);
TASK_PP(16'hB7A4,4);
TASK_PP(16'hB7A5,4);
TASK_PP(16'hB7A6,4);
TASK_PP(16'hB7A7,4);
TASK_PP(16'hB7A8,4);
TASK_PP(16'hB7A9,4);
TASK_PP(16'hB7AA,4);
TASK_PP(16'hB7AB,4);
TASK_PP(16'hB7AC,4);
TASK_PP(16'hB7AD,4);
TASK_PP(16'hB7AE,4);
TASK_PP(16'hB7AF,4);
TASK_PP(16'hB7B0,4);
TASK_PP(16'hB7B1,4);
TASK_PP(16'hB7B2,4);
TASK_PP(16'hB7B3,4);
TASK_PP(16'hB7B4,4);
TASK_PP(16'hB7B5,4);
TASK_PP(16'hB7B6,4);
TASK_PP(16'hB7B7,4);
TASK_PP(16'hB7B8,4);
TASK_PP(16'hB7B9,4);
TASK_PP(16'hB7BA,4);
TASK_PP(16'hB7BB,4);
TASK_PP(16'hB7BC,4);
TASK_PP(16'hB7BD,4);
TASK_PP(16'hB7BE,4);
TASK_PP(16'hB7BF,4);
TASK_PP(16'hB7C0,4);
TASK_PP(16'hB7C1,4);
TASK_PP(16'hB7C2,4);
TASK_PP(16'hB7C3,4);
TASK_PP(16'hB7C4,4);
TASK_PP(16'hB7C5,4);
TASK_PP(16'hB7C6,4);
TASK_PP(16'hB7C7,4);
TASK_PP(16'hB7C8,4);
TASK_PP(16'hB7C9,4);
TASK_PP(16'hB7CA,4);
TASK_PP(16'hB7CB,4);
TASK_PP(16'hB7CC,4);
TASK_PP(16'hB7CD,4);
TASK_PP(16'hB7CE,4);
TASK_PP(16'hB7CF,4);
TASK_PP(16'hB7D0,4);
TASK_PP(16'hB7D1,4);
TASK_PP(16'hB7D2,4);
TASK_PP(16'hB7D3,4);
TASK_PP(16'hB7D4,4);
TASK_PP(16'hB7D5,4);
TASK_PP(16'hB7D6,4);
TASK_PP(16'hB7D7,4);
TASK_PP(16'hB7D8,4);
TASK_PP(16'hB7D9,4);
TASK_PP(16'hB7DA,4);
TASK_PP(16'hB7DB,4);
TASK_PP(16'hB7DC,4);
TASK_PP(16'hB7DD,4);
TASK_PP(16'hB7DE,4);
TASK_PP(16'hB7DF,4);
TASK_PP(16'hB7E0,4);
TASK_PP(16'hB7E1,4);
TASK_PP(16'hB7E2,4);
TASK_PP(16'hB7E3,4);
TASK_PP(16'hB7E4,4);
TASK_PP(16'hB7E5,4);
TASK_PP(16'hB7E6,4);
TASK_PP(16'hB7E7,4);
TASK_PP(16'hB7E8,4);
TASK_PP(16'hB7E9,4);
TASK_PP(16'hB7EA,4);
TASK_PP(16'hB7EB,4);
TASK_PP(16'hB7EC,4);
TASK_PP(16'hB7ED,4);
TASK_PP(16'hB7EE,4);
TASK_PP(16'hB7EF,4);
TASK_PP(16'hB7F0,4);
TASK_PP(16'hB7F1,4);
TASK_PP(16'hB7F2,4);
TASK_PP(16'hB7F3,4);
TASK_PP(16'hB7F4,4);
TASK_PP(16'hB7F5,4);
TASK_PP(16'hB7F6,4);
TASK_PP(16'hB7F7,4);
TASK_PP(16'hB7F8,4);
TASK_PP(16'hB7F9,4);
TASK_PP(16'hB7FA,4);
TASK_PP(16'hB7FB,4);
TASK_PP(16'hB7FC,4);
TASK_PP(16'hB7FD,4);
TASK_PP(16'hB7FE,4);
TASK_PP(16'hB7FF,4);
TASK_PP(16'hB800,4);
TASK_PP(16'hB801,4);
TASK_PP(16'hB802,4);
TASK_PP(16'hB803,4);
TASK_PP(16'hB804,4);
TASK_PP(16'hB805,4);
TASK_PP(16'hB806,4);
TASK_PP(16'hB807,4);
TASK_PP(16'hB808,4);
TASK_PP(16'hB809,4);
TASK_PP(16'hB80A,4);
TASK_PP(16'hB80B,4);
TASK_PP(16'hB80C,4);
TASK_PP(16'hB80D,4);
TASK_PP(16'hB80E,4);
TASK_PP(16'hB80F,4);
TASK_PP(16'hB810,4);
TASK_PP(16'hB811,4);
TASK_PP(16'hB812,4);
TASK_PP(16'hB813,4);
TASK_PP(16'hB814,4);
TASK_PP(16'hB815,4);
TASK_PP(16'hB816,4);
TASK_PP(16'hB817,4);
TASK_PP(16'hB818,4);
TASK_PP(16'hB819,4);
TASK_PP(16'hB81A,4);
TASK_PP(16'hB81B,4);
TASK_PP(16'hB81C,4);
TASK_PP(16'hB81D,4);
TASK_PP(16'hB81E,4);
TASK_PP(16'hB81F,4);
TASK_PP(16'hB820,4);
TASK_PP(16'hB821,4);
TASK_PP(16'hB822,4);
TASK_PP(16'hB823,4);
TASK_PP(16'hB824,4);
TASK_PP(16'hB825,4);
TASK_PP(16'hB826,4);
TASK_PP(16'hB827,4);
TASK_PP(16'hB828,4);
TASK_PP(16'hB829,4);
TASK_PP(16'hB82A,4);
TASK_PP(16'hB82B,4);
TASK_PP(16'hB82C,4);
TASK_PP(16'hB82D,4);
TASK_PP(16'hB82E,4);
TASK_PP(16'hB82F,4);
TASK_PP(16'hB830,4);
TASK_PP(16'hB831,4);
TASK_PP(16'hB832,4);
TASK_PP(16'hB833,4);
TASK_PP(16'hB834,4);
TASK_PP(16'hB835,4);
TASK_PP(16'hB836,4);
TASK_PP(16'hB837,4);
TASK_PP(16'hB838,4);
TASK_PP(16'hB839,4);
TASK_PP(16'hB83A,4);
TASK_PP(16'hB83B,4);
TASK_PP(16'hB83C,4);
TASK_PP(16'hB83D,4);
TASK_PP(16'hB83E,4);
TASK_PP(16'hB83F,4);
TASK_PP(16'hB840,4);
TASK_PP(16'hB841,4);
TASK_PP(16'hB842,4);
TASK_PP(16'hB843,4);
TASK_PP(16'hB844,4);
TASK_PP(16'hB845,4);
TASK_PP(16'hB846,4);
TASK_PP(16'hB847,4);
TASK_PP(16'hB848,4);
TASK_PP(16'hB849,4);
TASK_PP(16'hB84A,4);
TASK_PP(16'hB84B,4);
TASK_PP(16'hB84C,4);
TASK_PP(16'hB84D,4);
TASK_PP(16'hB84E,4);
TASK_PP(16'hB84F,4);
TASK_PP(16'hB850,4);
TASK_PP(16'hB851,4);
TASK_PP(16'hB852,4);
TASK_PP(16'hB853,4);
TASK_PP(16'hB854,4);
TASK_PP(16'hB855,4);
TASK_PP(16'hB856,4);
TASK_PP(16'hB857,4);
TASK_PP(16'hB858,4);
TASK_PP(16'hB859,4);
TASK_PP(16'hB85A,4);
TASK_PP(16'hB85B,4);
TASK_PP(16'hB85C,4);
TASK_PP(16'hB85D,4);
TASK_PP(16'hB85E,4);
TASK_PP(16'hB85F,4);
TASK_PP(16'hB860,4);
TASK_PP(16'hB861,4);
TASK_PP(16'hB862,4);
TASK_PP(16'hB863,4);
TASK_PP(16'hB864,4);
TASK_PP(16'hB865,4);
TASK_PP(16'hB866,4);
TASK_PP(16'hB867,4);
TASK_PP(16'hB868,4);
TASK_PP(16'hB869,4);
TASK_PP(16'hB86A,4);
TASK_PP(16'hB86B,4);
TASK_PP(16'hB86C,4);
TASK_PP(16'hB86D,4);
TASK_PP(16'hB86E,4);
TASK_PP(16'hB86F,4);
TASK_PP(16'hB870,4);
TASK_PP(16'hB871,4);
TASK_PP(16'hB872,4);
TASK_PP(16'hB873,4);
TASK_PP(16'hB874,4);
TASK_PP(16'hB875,4);
TASK_PP(16'hB876,4);
TASK_PP(16'hB877,4);
TASK_PP(16'hB878,4);
TASK_PP(16'hB879,4);
TASK_PP(16'hB87A,4);
TASK_PP(16'hB87B,4);
TASK_PP(16'hB87C,4);
TASK_PP(16'hB87D,4);
TASK_PP(16'hB87E,4);
TASK_PP(16'hB87F,4);
TASK_PP(16'hB880,4);
TASK_PP(16'hB881,4);
TASK_PP(16'hB882,4);
TASK_PP(16'hB883,4);
TASK_PP(16'hB884,4);
TASK_PP(16'hB885,4);
TASK_PP(16'hB886,4);
TASK_PP(16'hB887,4);
TASK_PP(16'hB888,4);
TASK_PP(16'hB889,4);
TASK_PP(16'hB88A,4);
TASK_PP(16'hB88B,4);
TASK_PP(16'hB88C,4);
TASK_PP(16'hB88D,4);
TASK_PP(16'hB88E,4);
TASK_PP(16'hB88F,4);
TASK_PP(16'hB890,4);
TASK_PP(16'hB891,4);
TASK_PP(16'hB892,4);
TASK_PP(16'hB893,4);
TASK_PP(16'hB894,4);
TASK_PP(16'hB895,4);
TASK_PP(16'hB896,4);
TASK_PP(16'hB897,4);
TASK_PP(16'hB898,4);
TASK_PP(16'hB899,4);
TASK_PP(16'hB89A,4);
TASK_PP(16'hB89B,4);
TASK_PP(16'hB89C,4);
TASK_PP(16'hB89D,4);
TASK_PP(16'hB89E,4);
TASK_PP(16'hB89F,4);
TASK_PP(16'hB8A0,4);
TASK_PP(16'hB8A1,4);
TASK_PP(16'hB8A2,4);
TASK_PP(16'hB8A3,4);
TASK_PP(16'hB8A4,4);
TASK_PP(16'hB8A5,4);
TASK_PP(16'hB8A6,4);
TASK_PP(16'hB8A7,4);
TASK_PP(16'hB8A8,4);
TASK_PP(16'hB8A9,4);
TASK_PP(16'hB8AA,4);
TASK_PP(16'hB8AB,4);
TASK_PP(16'hB8AC,4);
TASK_PP(16'hB8AD,4);
TASK_PP(16'hB8AE,4);
TASK_PP(16'hB8AF,4);
TASK_PP(16'hB8B0,4);
TASK_PP(16'hB8B1,4);
TASK_PP(16'hB8B2,4);
TASK_PP(16'hB8B3,4);
TASK_PP(16'hB8B4,4);
TASK_PP(16'hB8B5,4);
TASK_PP(16'hB8B6,4);
TASK_PP(16'hB8B7,4);
TASK_PP(16'hB8B8,4);
TASK_PP(16'hB8B9,4);
TASK_PP(16'hB8BA,4);
TASK_PP(16'hB8BB,4);
TASK_PP(16'hB8BC,4);
TASK_PP(16'hB8BD,4);
TASK_PP(16'hB8BE,4);
TASK_PP(16'hB8BF,4);
TASK_PP(16'hB8C0,4);
TASK_PP(16'hB8C1,4);
TASK_PP(16'hB8C2,4);
TASK_PP(16'hB8C3,4);
TASK_PP(16'hB8C4,4);
TASK_PP(16'hB8C5,4);
TASK_PP(16'hB8C6,4);
TASK_PP(16'hB8C7,4);
TASK_PP(16'hB8C8,4);
TASK_PP(16'hB8C9,4);
TASK_PP(16'hB8CA,4);
TASK_PP(16'hB8CB,4);
TASK_PP(16'hB8CC,4);
TASK_PP(16'hB8CD,4);
TASK_PP(16'hB8CE,4);
TASK_PP(16'hB8CF,4);
TASK_PP(16'hB8D0,4);
TASK_PP(16'hB8D1,4);
TASK_PP(16'hB8D2,4);
TASK_PP(16'hB8D3,4);
TASK_PP(16'hB8D4,4);
TASK_PP(16'hB8D5,4);
TASK_PP(16'hB8D6,4);
TASK_PP(16'hB8D7,4);
TASK_PP(16'hB8D8,4);
TASK_PP(16'hB8D9,4);
TASK_PP(16'hB8DA,4);
TASK_PP(16'hB8DB,4);
TASK_PP(16'hB8DC,4);
TASK_PP(16'hB8DD,4);
TASK_PP(16'hB8DE,4);
TASK_PP(16'hB8DF,4);
TASK_PP(16'hB8E0,4);
TASK_PP(16'hB8E1,4);
TASK_PP(16'hB8E2,4);
TASK_PP(16'hB8E3,4);
TASK_PP(16'hB8E4,4);
TASK_PP(16'hB8E5,4);
TASK_PP(16'hB8E6,4);
TASK_PP(16'hB8E7,4);
TASK_PP(16'hB8E8,4);
TASK_PP(16'hB8E9,4);
TASK_PP(16'hB8EA,4);
TASK_PP(16'hB8EB,4);
TASK_PP(16'hB8EC,4);
TASK_PP(16'hB8ED,4);
TASK_PP(16'hB8EE,4);
TASK_PP(16'hB8EF,4);
TASK_PP(16'hB8F0,4);
TASK_PP(16'hB8F1,4);
TASK_PP(16'hB8F2,4);
TASK_PP(16'hB8F3,4);
TASK_PP(16'hB8F4,4);
TASK_PP(16'hB8F5,4);
TASK_PP(16'hB8F6,4);
TASK_PP(16'hB8F7,4);
TASK_PP(16'hB8F8,4);
TASK_PP(16'hB8F9,4);
TASK_PP(16'hB8FA,4);
TASK_PP(16'hB8FB,4);
TASK_PP(16'hB8FC,4);
TASK_PP(16'hB8FD,4);
TASK_PP(16'hB8FE,4);
TASK_PP(16'hB8FF,4);
TASK_PP(16'hB900,4);
TASK_PP(16'hB901,4);
TASK_PP(16'hB902,4);
TASK_PP(16'hB903,4);
TASK_PP(16'hB904,4);
TASK_PP(16'hB905,4);
TASK_PP(16'hB906,4);
TASK_PP(16'hB907,4);
TASK_PP(16'hB908,4);
TASK_PP(16'hB909,4);
TASK_PP(16'hB90A,4);
TASK_PP(16'hB90B,4);
TASK_PP(16'hB90C,4);
TASK_PP(16'hB90D,4);
TASK_PP(16'hB90E,4);
TASK_PP(16'hB90F,4);
TASK_PP(16'hB910,4);
TASK_PP(16'hB911,4);
TASK_PP(16'hB912,4);
TASK_PP(16'hB913,4);
TASK_PP(16'hB914,4);
TASK_PP(16'hB915,4);
TASK_PP(16'hB916,4);
TASK_PP(16'hB917,4);
TASK_PP(16'hB918,4);
TASK_PP(16'hB919,4);
TASK_PP(16'hB91A,4);
TASK_PP(16'hB91B,4);
TASK_PP(16'hB91C,4);
TASK_PP(16'hB91D,4);
TASK_PP(16'hB91E,4);
TASK_PP(16'hB91F,4);
TASK_PP(16'hB920,4);
TASK_PP(16'hB921,4);
TASK_PP(16'hB922,4);
TASK_PP(16'hB923,4);
TASK_PP(16'hB924,4);
TASK_PP(16'hB925,4);
TASK_PP(16'hB926,4);
TASK_PP(16'hB927,4);
TASK_PP(16'hB928,4);
TASK_PP(16'hB929,4);
TASK_PP(16'hB92A,4);
TASK_PP(16'hB92B,4);
TASK_PP(16'hB92C,4);
TASK_PP(16'hB92D,4);
TASK_PP(16'hB92E,4);
TASK_PP(16'hB92F,4);
TASK_PP(16'hB930,4);
TASK_PP(16'hB931,4);
TASK_PP(16'hB932,4);
TASK_PP(16'hB933,4);
TASK_PP(16'hB934,4);
TASK_PP(16'hB935,4);
TASK_PP(16'hB936,4);
TASK_PP(16'hB937,4);
TASK_PP(16'hB938,4);
TASK_PP(16'hB939,4);
TASK_PP(16'hB93A,4);
TASK_PP(16'hB93B,4);
TASK_PP(16'hB93C,4);
TASK_PP(16'hB93D,4);
TASK_PP(16'hB93E,4);
TASK_PP(16'hB93F,4);
TASK_PP(16'hB940,4);
TASK_PP(16'hB941,4);
TASK_PP(16'hB942,4);
TASK_PP(16'hB943,4);
TASK_PP(16'hB944,4);
TASK_PP(16'hB945,4);
TASK_PP(16'hB946,4);
TASK_PP(16'hB947,4);
TASK_PP(16'hB948,4);
TASK_PP(16'hB949,4);
TASK_PP(16'hB94A,4);
TASK_PP(16'hB94B,4);
TASK_PP(16'hB94C,4);
TASK_PP(16'hB94D,4);
TASK_PP(16'hB94E,4);
TASK_PP(16'hB94F,4);
TASK_PP(16'hB950,4);
TASK_PP(16'hB951,4);
TASK_PP(16'hB952,4);
TASK_PP(16'hB953,4);
TASK_PP(16'hB954,4);
TASK_PP(16'hB955,4);
TASK_PP(16'hB956,4);
TASK_PP(16'hB957,4);
TASK_PP(16'hB958,4);
TASK_PP(16'hB959,4);
TASK_PP(16'hB95A,4);
TASK_PP(16'hB95B,4);
TASK_PP(16'hB95C,4);
TASK_PP(16'hB95D,4);
TASK_PP(16'hB95E,4);
TASK_PP(16'hB95F,4);
TASK_PP(16'hB960,4);
TASK_PP(16'hB961,4);
TASK_PP(16'hB962,4);
TASK_PP(16'hB963,4);
TASK_PP(16'hB964,4);
TASK_PP(16'hB965,4);
TASK_PP(16'hB966,4);
TASK_PP(16'hB967,4);
TASK_PP(16'hB968,4);
TASK_PP(16'hB969,4);
TASK_PP(16'hB96A,4);
TASK_PP(16'hB96B,4);
TASK_PP(16'hB96C,4);
TASK_PP(16'hB96D,4);
TASK_PP(16'hB96E,4);
TASK_PP(16'hB96F,4);
TASK_PP(16'hB970,4);
TASK_PP(16'hB971,4);
TASK_PP(16'hB972,4);
TASK_PP(16'hB973,4);
TASK_PP(16'hB974,4);
TASK_PP(16'hB975,4);
TASK_PP(16'hB976,4);
TASK_PP(16'hB977,4);
TASK_PP(16'hB978,4);
TASK_PP(16'hB979,4);
TASK_PP(16'hB97A,4);
TASK_PP(16'hB97B,4);
TASK_PP(16'hB97C,4);
TASK_PP(16'hB97D,4);
TASK_PP(16'hB97E,4);
TASK_PP(16'hB97F,4);
TASK_PP(16'hB980,4);
TASK_PP(16'hB981,4);
TASK_PP(16'hB982,4);
TASK_PP(16'hB983,4);
TASK_PP(16'hB984,4);
TASK_PP(16'hB985,4);
TASK_PP(16'hB986,4);
TASK_PP(16'hB987,4);
TASK_PP(16'hB988,4);
TASK_PP(16'hB989,4);
TASK_PP(16'hB98A,4);
TASK_PP(16'hB98B,4);
TASK_PP(16'hB98C,4);
TASK_PP(16'hB98D,4);
TASK_PP(16'hB98E,4);
TASK_PP(16'hB98F,4);
TASK_PP(16'hB990,4);
TASK_PP(16'hB991,4);
TASK_PP(16'hB992,4);
TASK_PP(16'hB993,4);
TASK_PP(16'hB994,4);
TASK_PP(16'hB995,4);
TASK_PP(16'hB996,4);
TASK_PP(16'hB997,4);
TASK_PP(16'hB998,4);
TASK_PP(16'hB999,4);
TASK_PP(16'hB99A,4);
TASK_PP(16'hB99B,4);
TASK_PP(16'hB99C,4);
TASK_PP(16'hB99D,4);
TASK_PP(16'hB99E,4);
TASK_PP(16'hB99F,4);
TASK_PP(16'hB9A0,4);
TASK_PP(16'hB9A1,4);
TASK_PP(16'hB9A2,4);
TASK_PP(16'hB9A3,4);
TASK_PP(16'hB9A4,4);
TASK_PP(16'hB9A5,4);
TASK_PP(16'hB9A6,4);
TASK_PP(16'hB9A7,4);
TASK_PP(16'hB9A8,4);
TASK_PP(16'hB9A9,4);
TASK_PP(16'hB9AA,4);
TASK_PP(16'hB9AB,4);
TASK_PP(16'hB9AC,4);
TASK_PP(16'hB9AD,4);
TASK_PP(16'hB9AE,4);
TASK_PP(16'hB9AF,4);
TASK_PP(16'hB9B0,4);
TASK_PP(16'hB9B1,4);
TASK_PP(16'hB9B2,4);
TASK_PP(16'hB9B3,4);
TASK_PP(16'hB9B4,4);
TASK_PP(16'hB9B5,4);
TASK_PP(16'hB9B6,4);
TASK_PP(16'hB9B7,4);
TASK_PP(16'hB9B8,4);
TASK_PP(16'hB9B9,4);
TASK_PP(16'hB9BA,4);
TASK_PP(16'hB9BB,4);
TASK_PP(16'hB9BC,4);
TASK_PP(16'hB9BD,4);
TASK_PP(16'hB9BE,4);
TASK_PP(16'hB9BF,4);
TASK_PP(16'hB9C0,4);
TASK_PP(16'hB9C1,4);
TASK_PP(16'hB9C2,4);
TASK_PP(16'hB9C3,4);
TASK_PP(16'hB9C4,4);
TASK_PP(16'hB9C5,4);
TASK_PP(16'hB9C6,4);
TASK_PP(16'hB9C7,4);
TASK_PP(16'hB9C8,4);
TASK_PP(16'hB9C9,4);
TASK_PP(16'hB9CA,4);
TASK_PP(16'hB9CB,4);
TASK_PP(16'hB9CC,4);
TASK_PP(16'hB9CD,4);
TASK_PP(16'hB9CE,4);
TASK_PP(16'hB9CF,4);
TASK_PP(16'hB9D0,4);
TASK_PP(16'hB9D1,4);
TASK_PP(16'hB9D2,4);
TASK_PP(16'hB9D3,4);
TASK_PP(16'hB9D4,4);
TASK_PP(16'hB9D5,4);
TASK_PP(16'hB9D6,4);
TASK_PP(16'hB9D7,4);
TASK_PP(16'hB9D8,4);
TASK_PP(16'hB9D9,4);
TASK_PP(16'hB9DA,4);
TASK_PP(16'hB9DB,4);
TASK_PP(16'hB9DC,4);
TASK_PP(16'hB9DD,4);
TASK_PP(16'hB9DE,4);
TASK_PP(16'hB9DF,4);
TASK_PP(16'hB9E0,4);
TASK_PP(16'hB9E1,4);
TASK_PP(16'hB9E2,4);
TASK_PP(16'hB9E3,4);
TASK_PP(16'hB9E4,4);
TASK_PP(16'hB9E5,4);
TASK_PP(16'hB9E6,4);
TASK_PP(16'hB9E7,4);
TASK_PP(16'hB9E8,4);
TASK_PP(16'hB9E9,4);
TASK_PP(16'hB9EA,4);
TASK_PP(16'hB9EB,4);
TASK_PP(16'hB9EC,4);
TASK_PP(16'hB9ED,4);
TASK_PP(16'hB9EE,4);
TASK_PP(16'hB9EF,4);
TASK_PP(16'hB9F0,4);
TASK_PP(16'hB9F1,4);
TASK_PP(16'hB9F2,4);
TASK_PP(16'hB9F3,4);
TASK_PP(16'hB9F4,4);
TASK_PP(16'hB9F5,4);
TASK_PP(16'hB9F6,4);
TASK_PP(16'hB9F7,4);
TASK_PP(16'hB9F8,4);
TASK_PP(16'hB9F9,4);
TASK_PP(16'hB9FA,4);
TASK_PP(16'hB9FB,4);
TASK_PP(16'hB9FC,4);
TASK_PP(16'hB9FD,4);
TASK_PP(16'hB9FE,4);
TASK_PP(16'hB9FF,4);
TASK_PP(16'hBA00,4);
TASK_PP(16'hBA01,4);
TASK_PP(16'hBA02,4);
TASK_PP(16'hBA03,4);
TASK_PP(16'hBA04,4);
TASK_PP(16'hBA05,4);
TASK_PP(16'hBA06,4);
TASK_PP(16'hBA07,4);
TASK_PP(16'hBA08,4);
TASK_PP(16'hBA09,4);
TASK_PP(16'hBA0A,4);
TASK_PP(16'hBA0B,4);
TASK_PP(16'hBA0C,4);
TASK_PP(16'hBA0D,4);
TASK_PP(16'hBA0E,4);
TASK_PP(16'hBA0F,4);
TASK_PP(16'hBA10,4);
TASK_PP(16'hBA11,4);
TASK_PP(16'hBA12,4);
TASK_PP(16'hBA13,4);
TASK_PP(16'hBA14,4);
TASK_PP(16'hBA15,4);
TASK_PP(16'hBA16,4);
TASK_PP(16'hBA17,4);
TASK_PP(16'hBA18,4);
TASK_PP(16'hBA19,4);
TASK_PP(16'hBA1A,4);
TASK_PP(16'hBA1B,4);
TASK_PP(16'hBA1C,4);
TASK_PP(16'hBA1D,4);
TASK_PP(16'hBA1E,4);
TASK_PP(16'hBA1F,4);
TASK_PP(16'hBA20,4);
TASK_PP(16'hBA21,4);
TASK_PP(16'hBA22,4);
TASK_PP(16'hBA23,4);
TASK_PP(16'hBA24,4);
TASK_PP(16'hBA25,4);
TASK_PP(16'hBA26,4);
TASK_PP(16'hBA27,4);
TASK_PP(16'hBA28,4);
TASK_PP(16'hBA29,4);
TASK_PP(16'hBA2A,4);
TASK_PP(16'hBA2B,4);
TASK_PP(16'hBA2C,4);
TASK_PP(16'hBA2D,4);
TASK_PP(16'hBA2E,4);
TASK_PP(16'hBA2F,4);
TASK_PP(16'hBA30,4);
TASK_PP(16'hBA31,4);
TASK_PP(16'hBA32,4);
TASK_PP(16'hBA33,4);
TASK_PP(16'hBA34,4);
TASK_PP(16'hBA35,4);
TASK_PP(16'hBA36,4);
TASK_PP(16'hBA37,4);
TASK_PP(16'hBA38,4);
TASK_PP(16'hBA39,4);
TASK_PP(16'hBA3A,4);
TASK_PP(16'hBA3B,4);
TASK_PP(16'hBA3C,4);
TASK_PP(16'hBA3D,4);
TASK_PP(16'hBA3E,4);
TASK_PP(16'hBA3F,4);
TASK_PP(16'hBA40,4);
TASK_PP(16'hBA41,4);
TASK_PP(16'hBA42,4);
TASK_PP(16'hBA43,4);
TASK_PP(16'hBA44,4);
TASK_PP(16'hBA45,4);
TASK_PP(16'hBA46,4);
TASK_PP(16'hBA47,4);
TASK_PP(16'hBA48,4);
TASK_PP(16'hBA49,4);
TASK_PP(16'hBA4A,4);
TASK_PP(16'hBA4B,4);
TASK_PP(16'hBA4C,4);
TASK_PP(16'hBA4D,4);
TASK_PP(16'hBA4E,4);
TASK_PP(16'hBA4F,4);
TASK_PP(16'hBA50,4);
TASK_PP(16'hBA51,4);
TASK_PP(16'hBA52,4);
TASK_PP(16'hBA53,4);
TASK_PP(16'hBA54,4);
TASK_PP(16'hBA55,4);
TASK_PP(16'hBA56,4);
TASK_PP(16'hBA57,4);
TASK_PP(16'hBA58,4);
TASK_PP(16'hBA59,4);
TASK_PP(16'hBA5A,4);
TASK_PP(16'hBA5B,4);
TASK_PP(16'hBA5C,4);
TASK_PP(16'hBA5D,4);
TASK_PP(16'hBA5E,4);
TASK_PP(16'hBA5F,4);
TASK_PP(16'hBA60,4);
TASK_PP(16'hBA61,4);
TASK_PP(16'hBA62,4);
TASK_PP(16'hBA63,4);
TASK_PP(16'hBA64,4);
TASK_PP(16'hBA65,4);
TASK_PP(16'hBA66,4);
TASK_PP(16'hBA67,4);
TASK_PP(16'hBA68,4);
TASK_PP(16'hBA69,4);
TASK_PP(16'hBA6A,4);
TASK_PP(16'hBA6B,4);
TASK_PP(16'hBA6C,4);
TASK_PP(16'hBA6D,4);
TASK_PP(16'hBA6E,4);
TASK_PP(16'hBA6F,4);
TASK_PP(16'hBA70,4);
TASK_PP(16'hBA71,4);
TASK_PP(16'hBA72,4);
TASK_PP(16'hBA73,4);
TASK_PP(16'hBA74,4);
TASK_PP(16'hBA75,4);
TASK_PP(16'hBA76,4);
TASK_PP(16'hBA77,4);
TASK_PP(16'hBA78,4);
TASK_PP(16'hBA79,4);
TASK_PP(16'hBA7A,4);
TASK_PP(16'hBA7B,4);
TASK_PP(16'hBA7C,4);
TASK_PP(16'hBA7D,4);
TASK_PP(16'hBA7E,4);
TASK_PP(16'hBA7F,4);
TASK_PP(16'hBA80,4);
TASK_PP(16'hBA81,4);
TASK_PP(16'hBA82,4);
TASK_PP(16'hBA83,4);
TASK_PP(16'hBA84,4);
TASK_PP(16'hBA85,4);
TASK_PP(16'hBA86,4);
TASK_PP(16'hBA87,4);
TASK_PP(16'hBA88,4);
TASK_PP(16'hBA89,4);
TASK_PP(16'hBA8A,4);
TASK_PP(16'hBA8B,4);
TASK_PP(16'hBA8C,4);
TASK_PP(16'hBA8D,4);
TASK_PP(16'hBA8E,4);
TASK_PP(16'hBA8F,4);
TASK_PP(16'hBA90,4);
TASK_PP(16'hBA91,4);
TASK_PP(16'hBA92,4);
TASK_PP(16'hBA93,4);
TASK_PP(16'hBA94,4);
TASK_PP(16'hBA95,4);
TASK_PP(16'hBA96,4);
TASK_PP(16'hBA97,4);
TASK_PP(16'hBA98,4);
TASK_PP(16'hBA99,4);
TASK_PP(16'hBA9A,4);
TASK_PP(16'hBA9B,4);
TASK_PP(16'hBA9C,4);
TASK_PP(16'hBA9D,4);
TASK_PP(16'hBA9E,4);
TASK_PP(16'hBA9F,4);
TASK_PP(16'hBAA0,4);
TASK_PP(16'hBAA1,4);
TASK_PP(16'hBAA2,4);
TASK_PP(16'hBAA3,4);
TASK_PP(16'hBAA4,4);
TASK_PP(16'hBAA5,4);
TASK_PP(16'hBAA6,4);
TASK_PP(16'hBAA7,4);
TASK_PP(16'hBAA8,4);
TASK_PP(16'hBAA9,4);
TASK_PP(16'hBAAA,4);
TASK_PP(16'hBAAB,4);
TASK_PP(16'hBAAC,4);
TASK_PP(16'hBAAD,4);
TASK_PP(16'hBAAE,4);
TASK_PP(16'hBAAF,4);
TASK_PP(16'hBAB0,4);
TASK_PP(16'hBAB1,4);
TASK_PP(16'hBAB2,4);
TASK_PP(16'hBAB3,4);
TASK_PP(16'hBAB4,4);
TASK_PP(16'hBAB5,4);
TASK_PP(16'hBAB6,4);
TASK_PP(16'hBAB7,4);
TASK_PP(16'hBAB8,4);
TASK_PP(16'hBAB9,4);
TASK_PP(16'hBABA,4);
TASK_PP(16'hBABB,4);
TASK_PP(16'hBABC,4);
TASK_PP(16'hBABD,4);
TASK_PP(16'hBABE,4);
TASK_PP(16'hBABF,4);
TASK_PP(16'hBAC0,4);
TASK_PP(16'hBAC1,4);
TASK_PP(16'hBAC2,4);
TASK_PP(16'hBAC3,4);
TASK_PP(16'hBAC4,4);
TASK_PP(16'hBAC5,4);
TASK_PP(16'hBAC6,4);
TASK_PP(16'hBAC7,4);
TASK_PP(16'hBAC8,4);
TASK_PP(16'hBAC9,4);
TASK_PP(16'hBACA,4);
TASK_PP(16'hBACB,4);
TASK_PP(16'hBACC,4);
TASK_PP(16'hBACD,4);
TASK_PP(16'hBACE,4);
TASK_PP(16'hBACF,4);
TASK_PP(16'hBAD0,4);
TASK_PP(16'hBAD1,4);
TASK_PP(16'hBAD2,4);
TASK_PP(16'hBAD3,4);
TASK_PP(16'hBAD4,4);
TASK_PP(16'hBAD5,4);
TASK_PP(16'hBAD6,4);
TASK_PP(16'hBAD7,4);
TASK_PP(16'hBAD8,4);
TASK_PP(16'hBAD9,4);
TASK_PP(16'hBADA,4);
TASK_PP(16'hBADB,4);
TASK_PP(16'hBADC,4);
TASK_PP(16'hBADD,4);
TASK_PP(16'hBADE,4);
TASK_PP(16'hBADF,4);
TASK_PP(16'hBAE0,4);
TASK_PP(16'hBAE1,4);
TASK_PP(16'hBAE2,4);
TASK_PP(16'hBAE3,4);
TASK_PP(16'hBAE4,4);
TASK_PP(16'hBAE5,4);
TASK_PP(16'hBAE6,4);
TASK_PP(16'hBAE7,4);
TASK_PP(16'hBAE8,4);
TASK_PP(16'hBAE9,4);
TASK_PP(16'hBAEA,4);
TASK_PP(16'hBAEB,4);
TASK_PP(16'hBAEC,4);
TASK_PP(16'hBAED,4);
TASK_PP(16'hBAEE,4);
TASK_PP(16'hBAEF,4);
TASK_PP(16'hBAF0,4);
TASK_PP(16'hBAF1,4);
TASK_PP(16'hBAF2,4);
TASK_PP(16'hBAF3,4);
TASK_PP(16'hBAF4,4);
TASK_PP(16'hBAF5,4);
TASK_PP(16'hBAF6,4);
TASK_PP(16'hBAF7,4);
TASK_PP(16'hBAF8,4);
TASK_PP(16'hBAF9,4);
TASK_PP(16'hBAFA,4);
TASK_PP(16'hBAFB,4);
TASK_PP(16'hBAFC,4);
TASK_PP(16'hBAFD,4);
TASK_PP(16'hBAFE,4);
TASK_PP(16'hBAFF,4);
TASK_PP(16'hBB00,4);
TASK_PP(16'hBB01,4);
TASK_PP(16'hBB02,4);
TASK_PP(16'hBB03,4);
TASK_PP(16'hBB04,4);
TASK_PP(16'hBB05,4);
TASK_PP(16'hBB06,4);
TASK_PP(16'hBB07,4);
TASK_PP(16'hBB08,4);
TASK_PP(16'hBB09,4);
TASK_PP(16'hBB0A,4);
TASK_PP(16'hBB0B,4);
TASK_PP(16'hBB0C,4);
TASK_PP(16'hBB0D,4);
TASK_PP(16'hBB0E,4);
TASK_PP(16'hBB0F,4);
TASK_PP(16'hBB10,4);
TASK_PP(16'hBB11,4);
TASK_PP(16'hBB12,4);
TASK_PP(16'hBB13,4);
TASK_PP(16'hBB14,4);
TASK_PP(16'hBB15,4);
TASK_PP(16'hBB16,4);
TASK_PP(16'hBB17,4);
TASK_PP(16'hBB18,4);
TASK_PP(16'hBB19,4);
TASK_PP(16'hBB1A,4);
TASK_PP(16'hBB1B,4);
TASK_PP(16'hBB1C,4);
TASK_PP(16'hBB1D,4);
TASK_PP(16'hBB1E,4);
TASK_PP(16'hBB1F,4);
TASK_PP(16'hBB20,4);
TASK_PP(16'hBB21,4);
TASK_PP(16'hBB22,4);
TASK_PP(16'hBB23,4);
TASK_PP(16'hBB24,4);
TASK_PP(16'hBB25,4);
TASK_PP(16'hBB26,4);
TASK_PP(16'hBB27,4);
TASK_PP(16'hBB28,4);
TASK_PP(16'hBB29,4);
TASK_PP(16'hBB2A,4);
TASK_PP(16'hBB2B,4);
TASK_PP(16'hBB2C,4);
TASK_PP(16'hBB2D,4);
TASK_PP(16'hBB2E,4);
TASK_PP(16'hBB2F,4);
TASK_PP(16'hBB30,4);
TASK_PP(16'hBB31,4);
TASK_PP(16'hBB32,4);
TASK_PP(16'hBB33,4);
TASK_PP(16'hBB34,4);
TASK_PP(16'hBB35,4);
TASK_PP(16'hBB36,4);
TASK_PP(16'hBB37,4);
TASK_PP(16'hBB38,4);
TASK_PP(16'hBB39,4);
TASK_PP(16'hBB3A,4);
TASK_PP(16'hBB3B,4);
TASK_PP(16'hBB3C,4);
TASK_PP(16'hBB3D,4);
TASK_PP(16'hBB3E,4);
TASK_PP(16'hBB3F,4);
TASK_PP(16'hBB40,4);
TASK_PP(16'hBB41,4);
TASK_PP(16'hBB42,4);
TASK_PP(16'hBB43,4);
TASK_PP(16'hBB44,4);
TASK_PP(16'hBB45,4);
TASK_PP(16'hBB46,4);
TASK_PP(16'hBB47,4);
TASK_PP(16'hBB48,4);
TASK_PP(16'hBB49,4);
TASK_PP(16'hBB4A,4);
TASK_PP(16'hBB4B,4);
TASK_PP(16'hBB4C,4);
TASK_PP(16'hBB4D,4);
TASK_PP(16'hBB4E,4);
TASK_PP(16'hBB4F,4);
TASK_PP(16'hBB50,4);
TASK_PP(16'hBB51,4);
TASK_PP(16'hBB52,4);
TASK_PP(16'hBB53,4);
TASK_PP(16'hBB54,4);
TASK_PP(16'hBB55,4);
TASK_PP(16'hBB56,4);
TASK_PP(16'hBB57,4);
TASK_PP(16'hBB58,4);
TASK_PP(16'hBB59,4);
TASK_PP(16'hBB5A,4);
TASK_PP(16'hBB5B,4);
TASK_PP(16'hBB5C,4);
TASK_PP(16'hBB5D,4);
TASK_PP(16'hBB5E,4);
TASK_PP(16'hBB5F,4);
TASK_PP(16'hBB60,4);
TASK_PP(16'hBB61,4);
TASK_PP(16'hBB62,4);
TASK_PP(16'hBB63,4);
TASK_PP(16'hBB64,4);
TASK_PP(16'hBB65,4);
TASK_PP(16'hBB66,4);
TASK_PP(16'hBB67,4);
TASK_PP(16'hBB68,4);
TASK_PP(16'hBB69,4);
TASK_PP(16'hBB6A,4);
TASK_PP(16'hBB6B,4);
TASK_PP(16'hBB6C,4);
TASK_PP(16'hBB6D,4);
TASK_PP(16'hBB6E,4);
TASK_PP(16'hBB6F,4);
TASK_PP(16'hBB70,4);
TASK_PP(16'hBB71,4);
TASK_PP(16'hBB72,4);
TASK_PP(16'hBB73,4);
TASK_PP(16'hBB74,4);
TASK_PP(16'hBB75,4);
TASK_PP(16'hBB76,4);
TASK_PP(16'hBB77,4);
TASK_PP(16'hBB78,4);
TASK_PP(16'hBB79,4);
TASK_PP(16'hBB7A,4);
TASK_PP(16'hBB7B,4);
TASK_PP(16'hBB7C,4);
TASK_PP(16'hBB7D,4);
TASK_PP(16'hBB7E,4);
TASK_PP(16'hBB7F,4);
TASK_PP(16'hBB80,4);
TASK_PP(16'hBB81,4);
TASK_PP(16'hBB82,4);
TASK_PP(16'hBB83,4);
TASK_PP(16'hBB84,4);
TASK_PP(16'hBB85,4);
TASK_PP(16'hBB86,4);
TASK_PP(16'hBB87,4);
TASK_PP(16'hBB88,4);
TASK_PP(16'hBB89,4);
TASK_PP(16'hBB8A,4);
TASK_PP(16'hBB8B,4);
TASK_PP(16'hBB8C,4);
TASK_PP(16'hBB8D,4);
TASK_PP(16'hBB8E,4);
TASK_PP(16'hBB8F,4);
TASK_PP(16'hBB90,4);
TASK_PP(16'hBB91,4);
TASK_PP(16'hBB92,4);
TASK_PP(16'hBB93,4);
TASK_PP(16'hBB94,4);
TASK_PP(16'hBB95,4);
TASK_PP(16'hBB96,4);
TASK_PP(16'hBB97,4);
TASK_PP(16'hBB98,4);
TASK_PP(16'hBB99,4);
TASK_PP(16'hBB9A,4);
TASK_PP(16'hBB9B,4);
TASK_PP(16'hBB9C,4);
TASK_PP(16'hBB9D,4);
TASK_PP(16'hBB9E,4);
TASK_PP(16'hBB9F,4);
TASK_PP(16'hBBA0,4);
TASK_PP(16'hBBA1,4);
TASK_PP(16'hBBA2,4);
TASK_PP(16'hBBA3,4);
TASK_PP(16'hBBA4,4);
TASK_PP(16'hBBA5,4);
TASK_PP(16'hBBA6,4);
TASK_PP(16'hBBA7,4);
TASK_PP(16'hBBA8,4);
TASK_PP(16'hBBA9,4);
TASK_PP(16'hBBAA,4);
TASK_PP(16'hBBAB,4);
TASK_PP(16'hBBAC,4);
TASK_PP(16'hBBAD,4);
TASK_PP(16'hBBAE,4);
TASK_PP(16'hBBAF,4);
TASK_PP(16'hBBB0,4);
TASK_PP(16'hBBB1,4);
TASK_PP(16'hBBB2,4);
TASK_PP(16'hBBB3,4);
TASK_PP(16'hBBB4,4);
TASK_PP(16'hBBB5,4);
TASK_PP(16'hBBB6,4);
TASK_PP(16'hBBB7,4);
TASK_PP(16'hBBB8,4);
TASK_PP(16'hBBB9,4);
TASK_PP(16'hBBBA,4);
TASK_PP(16'hBBBB,4);
TASK_PP(16'hBBBC,4);
TASK_PP(16'hBBBD,4);
TASK_PP(16'hBBBE,4);
TASK_PP(16'hBBBF,4);
TASK_PP(16'hBBC0,4);
TASK_PP(16'hBBC1,4);
TASK_PP(16'hBBC2,4);
TASK_PP(16'hBBC3,4);
TASK_PP(16'hBBC4,4);
TASK_PP(16'hBBC5,4);
TASK_PP(16'hBBC6,4);
TASK_PP(16'hBBC7,4);
TASK_PP(16'hBBC8,4);
TASK_PP(16'hBBC9,4);
TASK_PP(16'hBBCA,4);
TASK_PP(16'hBBCB,4);
TASK_PP(16'hBBCC,4);
TASK_PP(16'hBBCD,4);
TASK_PP(16'hBBCE,4);
TASK_PP(16'hBBCF,4);
TASK_PP(16'hBBD0,4);
TASK_PP(16'hBBD1,4);
TASK_PP(16'hBBD2,4);
TASK_PP(16'hBBD3,4);
TASK_PP(16'hBBD4,4);
TASK_PP(16'hBBD5,4);
TASK_PP(16'hBBD6,4);
TASK_PP(16'hBBD7,4);
TASK_PP(16'hBBD8,4);
TASK_PP(16'hBBD9,4);
TASK_PP(16'hBBDA,4);
TASK_PP(16'hBBDB,4);
TASK_PP(16'hBBDC,4);
TASK_PP(16'hBBDD,4);
TASK_PP(16'hBBDE,4);
TASK_PP(16'hBBDF,4);
TASK_PP(16'hBBE0,4);
TASK_PP(16'hBBE1,4);
TASK_PP(16'hBBE2,4);
TASK_PP(16'hBBE3,4);
TASK_PP(16'hBBE4,4);
TASK_PP(16'hBBE5,4);
TASK_PP(16'hBBE6,4);
TASK_PP(16'hBBE7,4);
TASK_PP(16'hBBE8,4);
TASK_PP(16'hBBE9,4);
TASK_PP(16'hBBEA,4);
TASK_PP(16'hBBEB,4);
TASK_PP(16'hBBEC,4);
TASK_PP(16'hBBED,4);
TASK_PP(16'hBBEE,4);
TASK_PP(16'hBBEF,4);
TASK_PP(16'hBBF0,4);
TASK_PP(16'hBBF1,4);
TASK_PP(16'hBBF2,4);
TASK_PP(16'hBBF3,4);
TASK_PP(16'hBBF4,4);
TASK_PP(16'hBBF5,4);
TASK_PP(16'hBBF6,4);
TASK_PP(16'hBBF7,4);
TASK_PP(16'hBBF8,4);
TASK_PP(16'hBBF9,4);
TASK_PP(16'hBBFA,4);
TASK_PP(16'hBBFB,4);
TASK_PP(16'hBBFC,4);
TASK_PP(16'hBBFD,4);
TASK_PP(16'hBBFE,4);
TASK_PP(16'hBBFF,4);
TASK_PP(16'hBC00,4);
TASK_PP(16'hBC01,4);
TASK_PP(16'hBC02,4);
TASK_PP(16'hBC03,4);
TASK_PP(16'hBC04,4);
TASK_PP(16'hBC05,4);
TASK_PP(16'hBC06,4);
TASK_PP(16'hBC07,4);
TASK_PP(16'hBC08,4);
TASK_PP(16'hBC09,4);
TASK_PP(16'hBC0A,4);
TASK_PP(16'hBC0B,4);
TASK_PP(16'hBC0C,4);
TASK_PP(16'hBC0D,4);
TASK_PP(16'hBC0E,4);
TASK_PP(16'hBC0F,4);
TASK_PP(16'hBC10,4);
TASK_PP(16'hBC11,4);
TASK_PP(16'hBC12,4);
TASK_PP(16'hBC13,4);
TASK_PP(16'hBC14,4);
TASK_PP(16'hBC15,4);
TASK_PP(16'hBC16,4);
TASK_PP(16'hBC17,4);
TASK_PP(16'hBC18,4);
TASK_PP(16'hBC19,4);
TASK_PP(16'hBC1A,4);
TASK_PP(16'hBC1B,4);
TASK_PP(16'hBC1C,4);
TASK_PP(16'hBC1D,4);
TASK_PP(16'hBC1E,4);
TASK_PP(16'hBC1F,4);
TASK_PP(16'hBC20,4);
TASK_PP(16'hBC21,4);
TASK_PP(16'hBC22,4);
TASK_PP(16'hBC23,4);
TASK_PP(16'hBC24,4);
TASK_PP(16'hBC25,4);
TASK_PP(16'hBC26,4);
TASK_PP(16'hBC27,4);
TASK_PP(16'hBC28,4);
TASK_PP(16'hBC29,4);
TASK_PP(16'hBC2A,4);
TASK_PP(16'hBC2B,4);
TASK_PP(16'hBC2C,4);
TASK_PP(16'hBC2D,4);
TASK_PP(16'hBC2E,4);
TASK_PP(16'hBC2F,4);
TASK_PP(16'hBC30,4);
TASK_PP(16'hBC31,4);
TASK_PP(16'hBC32,4);
TASK_PP(16'hBC33,4);
TASK_PP(16'hBC34,4);
TASK_PP(16'hBC35,4);
TASK_PP(16'hBC36,4);
TASK_PP(16'hBC37,4);
TASK_PP(16'hBC38,4);
TASK_PP(16'hBC39,4);
TASK_PP(16'hBC3A,4);
TASK_PP(16'hBC3B,4);
TASK_PP(16'hBC3C,4);
TASK_PP(16'hBC3D,4);
TASK_PP(16'hBC3E,4);
TASK_PP(16'hBC3F,4);
TASK_PP(16'hBC40,4);
TASK_PP(16'hBC41,4);
TASK_PP(16'hBC42,4);
TASK_PP(16'hBC43,4);
TASK_PP(16'hBC44,4);
TASK_PP(16'hBC45,4);
TASK_PP(16'hBC46,4);
TASK_PP(16'hBC47,4);
TASK_PP(16'hBC48,4);
TASK_PP(16'hBC49,4);
TASK_PP(16'hBC4A,4);
TASK_PP(16'hBC4B,4);
TASK_PP(16'hBC4C,4);
TASK_PP(16'hBC4D,4);
TASK_PP(16'hBC4E,4);
TASK_PP(16'hBC4F,4);
TASK_PP(16'hBC50,4);
TASK_PP(16'hBC51,4);
TASK_PP(16'hBC52,4);
TASK_PP(16'hBC53,4);
TASK_PP(16'hBC54,4);
TASK_PP(16'hBC55,4);
TASK_PP(16'hBC56,4);
TASK_PP(16'hBC57,4);
TASK_PP(16'hBC58,4);
TASK_PP(16'hBC59,4);
TASK_PP(16'hBC5A,4);
TASK_PP(16'hBC5B,4);
TASK_PP(16'hBC5C,4);
TASK_PP(16'hBC5D,4);
TASK_PP(16'hBC5E,4);
TASK_PP(16'hBC5F,4);
TASK_PP(16'hBC60,4);
TASK_PP(16'hBC61,4);
TASK_PP(16'hBC62,4);
TASK_PP(16'hBC63,4);
TASK_PP(16'hBC64,4);
TASK_PP(16'hBC65,4);
TASK_PP(16'hBC66,4);
TASK_PP(16'hBC67,4);
TASK_PP(16'hBC68,4);
TASK_PP(16'hBC69,4);
TASK_PP(16'hBC6A,4);
TASK_PP(16'hBC6B,4);
TASK_PP(16'hBC6C,4);
TASK_PP(16'hBC6D,4);
TASK_PP(16'hBC6E,4);
TASK_PP(16'hBC6F,4);
TASK_PP(16'hBC70,4);
TASK_PP(16'hBC71,4);
TASK_PP(16'hBC72,4);
TASK_PP(16'hBC73,4);
TASK_PP(16'hBC74,4);
TASK_PP(16'hBC75,4);
TASK_PP(16'hBC76,4);
TASK_PP(16'hBC77,4);
TASK_PP(16'hBC78,4);
TASK_PP(16'hBC79,4);
TASK_PP(16'hBC7A,4);
TASK_PP(16'hBC7B,4);
TASK_PP(16'hBC7C,4);
TASK_PP(16'hBC7D,4);
TASK_PP(16'hBC7E,4);
TASK_PP(16'hBC7F,4);
TASK_PP(16'hBC80,4);
TASK_PP(16'hBC81,4);
TASK_PP(16'hBC82,4);
TASK_PP(16'hBC83,4);
TASK_PP(16'hBC84,4);
TASK_PP(16'hBC85,4);
TASK_PP(16'hBC86,4);
TASK_PP(16'hBC87,4);
TASK_PP(16'hBC88,4);
TASK_PP(16'hBC89,4);
TASK_PP(16'hBC8A,4);
TASK_PP(16'hBC8B,4);
TASK_PP(16'hBC8C,4);
TASK_PP(16'hBC8D,4);
TASK_PP(16'hBC8E,4);
TASK_PP(16'hBC8F,4);
TASK_PP(16'hBC90,4);
TASK_PP(16'hBC91,4);
TASK_PP(16'hBC92,4);
TASK_PP(16'hBC93,4);
TASK_PP(16'hBC94,4);
TASK_PP(16'hBC95,4);
TASK_PP(16'hBC96,4);
TASK_PP(16'hBC97,4);
TASK_PP(16'hBC98,4);
TASK_PP(16'hBC99,4);
TASK_PP(16'hBC9A,4);
TASK_PP(16'hBC9B,4);
TASK_PP(16'hBC9C,4);
TASK_PP(16'hBC9D,4);
TASK_PP(16'hBC9E,4);
TASK_PP(16'hBC9F,4);
TASK_PP(16'hBCA0,4);
TASK_PP(16'hBCA1,4);
TASK_PP(16'hBCA2,4);
TASK_PP(16'hBCA3,4);
TASK_PP(16'hBCA4,4);
TASK_PP(16'hBCA5,4);
TASK_PP(16'hBCA6,4);
TASK_PP(16'hBCA7,4);
TASK_PP(16'hBCA8,4);
TASK_PP(16'hBCA9,4);
TASK_PP(16'hBCAA,4);
TASK_PP(16'hBCAB,4);
TASK_PP(16'hBCAC,4);
TASK_PP(16'hBCAD,4);
TASK_PP(16'hBCAE,4);
TASK_PP(16'hBCAF,4);
TASK_PP(16'hBCB0,4);
TASK_PP(16'hBCB1,4);
TASK_PP(16'hBCB2,4);
TASK_PP(16'hBCB3,4);
TASK_PP(16'hBCB4,4);
TASK_PP(16'hBCB5,4);
TASK_PP(16'hBCB6,4);
TASK_PP(16'hBCB7,4);
TASK_PP(16'hBCB8,4);
TASK_PP(16'hBCB9,4);
TASK_PP(16'hBCBA,4);
TASK_PP(16'hBCBB,4);
TASK_PP(16'hBCBC,4);
TASK_PP(16'hBCBD,4);
TASK_PP(16'hBCBE,4);
TASK_PP(16'hBCBF,4);
TASK_PP(16'hBCC0,4);
TASK_PP(16'hBCC1,4);
TASK_PP(16'hBCC2,4);
TASK_PP(16'hBCC3,4);
TASK_PP(16'hBCC4,4);
TASK_PP(16'hBCC5,4);
TASK_PP(16'hBCC6,4);
TASK_PP(16'hBCC7,4);
TASK_PP(16'hBCC8,4);
TASK_PP(16'hBCC9,4);
TASK_PP(16'hBCCA,4);
TASK_PP(16'hBCCB,4);
TASK_PP(16'hBCCC,4);
TASK_PP(16'hBCCD,4);
TASK_PP(16'hBCCE,4);
TASK_PP(16'hBCCF,4);
TASK_PP(16'hBCD0,4);
TASK_PP(16'hBCD1,4);
TASK_PP(16'hBCD2,4);
TASK_PP(16'hBCD3,4);
TASK_PP(16'hBCD4,4);
TASK_PP(16'hBCD5,4);
TASK_PP(16'hBCD6,4);
TASK_PP(16'hBCD7,4);
TASK_PP(16'hBCD8,4);
TASK_PP(16'hBCD9,4);
TASK_PP(16'hBCDA,4);
TASK_PP(16'hBCDB,4);
TASK_PP(16'hBCDC,4);
TASK_PP(16'hBCDD,4);
TASK_PP(16'hBCDE,4);
TASK_PP(16'hBCDF,4);
TASK_PP(16'hBCE0,4);
TASK_PP(16'hBCE1,4);
TASK_PP(16'hBCE2,4);
TASK_PP(16'hBCE3,4);
TASK_PP(16'hBCE4,4);
TASK_PP(16'hBCE5,4);
TASK_PP(16'hBCE6,4);
TASK_PP(16'hBCE7,4);
TASK_PP(16'hBCE8,4);
TASK_PP(16'hBCE9,4);
TASK_PP(16'hBCEA,4);
TASK_PP(16'hBCEB,4);
TASK_PP(16'hBCEC,4);
TASK_PP(16'hBCED,4);
TASK_PP(16'hBCEE,4);
TASK_PP(16'hBCEF,4);
TASK_PP(16'hBCF0,4);
TASK_PP(16'hBCF1,4);
TASK_PP(16'hBCF2,4);
TASK_PP(16'hBCF3,4);
TASK_PP(16'hBCF4,4);
TASK_PP(16'hBCF5,4);
TASK_PP(16'hBCF6,4);
TASK_PP(16'hBCF7,4);
TASK_PP(16'hBCF8,4);
TASK_PP(16'hBCF9,4);
TASK_PP(16'hBCFA,4);
TASK_PP(16'hBCFB,4);
TASK_PP(16'hBCFC,4);
TASK_PP(16'hBCFD,4);
TASK_PP(16'hBCFE,4);
TASK_PP(16'hBCFF,4);
TASK_PP(16'hBD00,4);
TASK_PP(16'hBD01,4);
TASK_PP(16'hBD02,4);
TASK_PP(16'hBD03,4);
TASK_PP(16'hBD04,4);
TASK_PP(16'hBD05,4);
TASK_PP(16'hBD06,4);
TASK_PP(16'hBD07,4);
TASK_PP(16'hBD08,4);
TASK_PP(16'hBD09,4);
TASK_PP(16'hBD0A,4);
TASK_PP(16'hBD0B,4);
TASK_PP(16'hBD0C,4);
TASK_PP(16'hBD0D,4);
TASK_PP(16'hBD0E,4);
TASK_PP(16'hBD0F,4);
TASK_PP(16'hBD10,4);
TASK_PP(16'hBD11,4);
TASK_PP(16'hBD12,4);
TASK_PP(16'hBD13,4);
TASK_PP(16'hBD14,4);
TASK_PP(16'hBD15,4);
TASK_PP(16'hBD16,4);
TASK_PP(16'hBD17,4);
TASK_PP(16'hBD18,4);
TASK_PP(16'hBD19,4);
TASK_PP(16'hBD1A,4);
TASK_PP(16'hBD1B,4);
TASK_PP(16'hBD1C,4);
TASK_PP(16'hBD1D,4);
TASK_PP(16'hBD1E,4);
TASK_PP(16'hBD1F,4);
TASK_PP(16'hBD20,4);
TASK_PP(16'hBD21,4);
TASK_PP(16'hBD22,4);
TASK_PP(16'hBD23,4);
TASK_PP(16'hBD24,4);
TASK_PP(16'hBD25,4);
TASK_PP(16'hBD26,4);
TASK_PP(16'hBD27,4);
TASK_PP(16'hBD28,4);
TASK_PP(16'hBD29,4);
TASK_PP(16'hBD2A,4);
TASK_PP(16'hBD2B,4);
TASK_PP(16'hBD2C,4);
TASK_PP(16'hBD2D,4);
TASK_PP(16'hBD2E,4);
TASK_PP(16'hBD2F,4);
TASK_PP(16'hBD30,4);
TASK_PP(16'hBD31,4);
TASK_PP(16'hBD32,4);
TASK_PP(16'hBD33,4);
TASK_PP(16'hBD34,4);
TASK_PP(16'hBD35,4);
TASK_PP(16'hBD36,4);
TASK_PP(16'hBD37,4);
TASK_PP(16'hBD38,4);
TASK_PP(16'hBD39,4);
TASK_PP(16'hBD3A,4);
TASK_PP(16'hBD3B,4);
TASK_PP(16'hBD3C,4);
TASK_PP(16'hBD3D,4);
TASK_PP(16'hBD3E,4);
TASK_PP(16'hBD3F,4);
TASK_PP(16'hBD40,4);
TASK_PP(16'hBD41,4);
TASK_PP(16'hBD42,4);
TASK_PP(16'hBD43,4);
TASK_PP(16'hBD44,4);
TASK_PP(16'hBD45,4);
TASK_PP(16'hBD46,4);
TASK_PP(16'hBD47,4);
TASK_PP(16'hBD48,4);
TASK_PP(16'hBD49,4);
TASK_PP(16'hBD4A,4);
TASK_PP(16'hBD4B,4);
TASK_PP(16'hBD4C,4);
TASK_PP(16'hBD4D,4);
TASK_PP(16'hBD4E,4);
TASK_PP(16'hBD4F,4);
TASK_PP(16'hBD50,4);
TASK_PP(16'hBD51,4);
TASK_PP(16'hBD52,4);
TASK_PP(16'hBD53,4);
TASK_PP(16'hBD54,4);
TASK_PP(16'hBD55,4);
TASK_PP(16'hBD56,4);
TASK_PP(16'hBD57,4);
TASK_PP(16'hBD58,4);
TASK_PP(16'hBD59,4);
TASK_PP(16'hBD5A,4);
TASK_PP(16'hBD5B,4);
TASK_PP(16'hBD5C,4);
TASK_PP(16'hBD5D,4);
TASK_PP(16'hBD5E,4);
TASK_PP(16'hBD5F,4);
TASK_PP(16'hBD60,4);
TASK_PP(16'hBD61,4);
TASK_PP(16'hBD62,4);
TASK_PP(16'hBD63,4);
TASK_PP(16'hBD64,4);
TASK_PP(16'hBD65,4);
TASK_PP(16'hBD66,4);
TASK_PP(16'hBD67,4);
TASK_PP(16'hBD68,4);
TASK_PP(16'hBD69,4);
TASK_PP(16'hBD6A,4);
TASK_PP(16'hBD6B,4);
TASK_PP(16'hBD6C,4);
TASK_PP(16'hBD6D,4);
TASK_PP(16'hBD6E,4);
TASK_PP(16'hBD6F,4);
TASK_PP(16'hBD70,4);
TASK_PP(16'hBD71,4);
TASK_PP(16'hBD72,4);
TASK_PP(16'hBD73,4);
TASK_PP(16'hBD74,4);
TASK_PP(16'hBD75,4);
TASK_PP(16'hBD76,4);
TASK_PP(16'hBD77,4);
TASK_PP(16'hBD78,4);
TASK_PP(16'hBD79,4);
TASK_PP(16'hBD7A,4);
TASK_PP(16'hBD7B,4);
TASK_PP(16'hBD7C,4);
TASK_PP(16'hBD7D,4);
TASK_PP(16'hBD7E,4);
TASK_PP(16'hBD7F,4);
TASK_PP(16'hBD80,4);
TASK_PP(16'hBD81,4);
TASK_PP(16'hBD82,4);
TASK_PP(16'hBD83,4);
TASK_PP(16'hBD84,4);
TASK_PP(16'hBD85,4);
TASK_PP(16'hBD86,4);
TASK_PP(16'hBD87,4);
TASK_PP(16'hBD88,4);
TASK_PP(16'hBD89,4);
TASK_PP(16'hBD8A,4);
TASK_PP(16'hBD8B,4);
TASK_PP(16'hBD8C,4);
TASK_PP(16'hBD8D,4);
TASK_PP(16'hBD8E,4);
TASK_PP(16'hBD8F,4);
TASK_PP(16'hBD90,4);
TASK_PP(16'hBD91,4);
TASK_PP(16'hBD92,4);
TASK_PP(16'hBD93,4);
TASK_PP(16'hBD94,4);
TASK_PP(16'hBD95,4);
TASK_PP(16'hBD96,4);
TASK_PP(16'hBD97,4);
TASK_PP(16'hBD98,4);
TASK_PP(16'hBD99,4);
TASK_PP(16'hBD9A,4);
TASK_PP(16'hBD9B,4);
TASK_PP(16'hBD9C,4);
TASK_PP(16'hBD9D,4);
TASK_PP(16'hBD9E,4);
TASK_PP(16'hBD9F,4);
TASK_PP(16'hBDA0,4);
TASK_PP(16'hBDA1,4);
TASK_PP(16'hBDA2,4);
TASK_PP(16'hBDA3,4);
TASK_PP(16'hBDA4,4);
TASK_PP(16'hBDA5,4);
TASK_PP(16'hBDA6,4);
TASK_PP(16'hBDA7,4);
TASK_PP(16'hBDA8,4);
TASK_PP(16'hBDA9,4);
TASK_PP(16'hBDAA,4);
TASK_PP(16'hBDAB,4);
TASK_PP(16'hBDAC,4);
TASK_PP(16'hBDAD,4);
TASK_PP(16'hBDAE,4);
TASK_PP(16'hBDAF,4);
TASK_PP(16'hBDB0,4);
TASK_PP(16'hBDB1,4);
TASK_PP(16'hBDB2,4);
TASK_PP(16'hBDB3,4);
TASK_PP(16'hBDB4,4);
TASK_PP(16'hBDB5,4);
TASK_PP(16'hBDB6,4);
TASK_PP(16'hBDB7,4);
TASK_PP(16'hBDB8,4);
TASK_PP(16'hBDB9,4);
TASK_PP(16'hBDBA,4);
TASK_PP(16'hBDBB,4);
TASK_PP(16'hBDBC,4);
TASK_PP(16'hBDBD,4);
TASK_PP(16'hBDBE,4);
TASK_PP(16'hBDBF,4);
TASK_PP(16'hBDC0,4);
TASK_PP(16'hBDC1,4);
TASK_PP(16'hBDC2,4);
TASK_PP(16'hBDC3,4);
TASK_PP(16'hBDC4,4);
TASK_PP(16'hBDC5,4);
TASK_PP(16'hBDC6,4);
TASK_PP(16'hBDC7,4);
TASK_PP(16'hBDC8,4);
TASK_PP(16'hBDC9,4);
TASK_PP(16'hBDCA,4);
TASK_PP(16'hBDCB,4);
TASK_PP(16'hBDCC,4);
TASK_PP(16'hBDCD,4);
TASK_PP(16'hBDCE,4);
TASK_PP(16'hBDCF,4);
TASK_PP(16'hBDD0,4);
TASK_PP(16'hBDD1,4);
TASK_PP(16'hBDD2,4);
TASK_PP(16'hBDD3,4);
TASK_PP(16'hBDD4,4);
TASK_PP(16'hBDD5,4);
TASK_PP(16'hBDD6,4);
TASK_PP(16'hBDD7,4);
TASK_PP(16'hBDD8,4);
TASK_PP(16'hBDD9,4);
TASK_PP(16'hBDDA,4);
TASK_PP(16'hBDDB,4);
TASK_PP(16'hBDDC,4);
TASK_PP(16'hBDDD,4);
TASK_PP(16'hBDDE,4);
TASK_PP(16'hBDDF,4);
TASK_PP(16'hBDE0,4);
TASK_PP(16'hBDE1,4);
TASK_PP(16'hBDE2,4);
TASK_PP(16'hBDE3,4);
TASK_PP(16'hBDE4,4);
TASK_PP(16'hBDE5,4);
TASK_PP(16'hBDE6,4);
TASK_PP(16'hBDE7,4);
TASK_PP(16'hBDE8,4);
TASK_PP(16'hBDE9,4);
TASK_PP(16'hBDEA,4);
TASK_PP(16'hBDEB,4);
TASK_PP(16'hBDEC,4);
TASK_PP(16'hBDED,4);
TASK_PP(16'hBDEE,4);
TASK_PP(16'hBDEF,4);
TASK_PP(16'hBDF0,4);
TASK_PP(16'hBDF1,4);
TASK_PP(16'hBDF2,4);
TASK_PP(16'hBDF3,4);
TASK_PP(16'hBDF4,4);
TASK_PP(16'hBDF5,4);
TASK_PP(16'hBDF6,4);
TASK_PP(16'hBDF7,4);
TASK_PP(16'hBDF8,4);
TASK_PP(16'hBDF9,4);
TASK_PP(16'hBDFA,4);
TASK_PP(16'hBDFB,4);
TASK_PP(16'hBDFC,4);
TASK_PP(16'hBDFD,4);
TASK_PP(16'hBDFE,4);
TASK_PP(16'hBDFF,4);
TASK_PP(16'hBE00,4);
TASK_PP(16'hBE01,4);
TASK_PP(16'hBE02,4);
TASK_PP(16'hBE03,4);
TASK_PP(16'hBE04,4);
TASK_PP(16'hBE05,4);
TASK_PP(16'hBE06,4);
TASK_PP(16'hBE07,4);
TASK_PP(16'hBE08,4);
TASK_PP(16'hBE09,4);
TASK_PP(16'hBE0A,4);
TASK_PP(16'hBE0B,4);
TASK_PP(16'hBE0C,4);
TASK_PP(16'hBE0D,4);
TASK_PP(16'hBE0E,4);
TASK_PP(16'hBE0F,4);
TASK_PP(16'hBE10,4);
TASK_PP(16'hBE11,4);
TASK_PP(16'hBE12,4);
TASK_PP(16'hBE13,4);
TASK_PP(16'hBE14,4);
TASK_PP(16'hBE15,4);
TASK_PP(16'hBE16,4);
TASK_PP(16'hBE17,4);
TASK_PP(16'hBE18,4);
TASK_PP(16'hBE19,4);
TASK_PP(16'hBE1A,4);
TASK_PP(16'hBE1B,4);
TASK_PP(16'hBE1C,4);
TASK_PP(16'hBE1D,4);
TASK_PP(16'hBE1E,4);
TASK_PP(16'hBE1F,4);
TASK_PP(16'hBE20,4);
TASK_PP(16'hBE21,4);
TASK_PP(16'hBE22,4);
TASK_PP(16'hBE23,4);
TASK_PP(16'hBE24,4);
TASK_PP(16'hBE25,4);
TASK_PP(16'hBE26,4);
TASK_PP(16'hBE27,4);
TASK_PP(16'hBE28,4);
TASK_PP(16'hBE29,4);
TASK_PP(16'hBE2A,4);
TASK_PP(16'hBE2B,4);
TASK_PP(16'hBE2C,4);
TASK_PP(16'hBE2D,4);
TASK_PP(16'hBE2E,4);
TASK_PP(16'hBE2F,4);
TASK_PP(16'hBE30,4);
TASK_PP(16'hBE31,4);
TASK_PP(16'hBE32,4);
TASK_PP(16'hBE33,4);
TASK_PP(16'hBE34,4);
TASK_PP(16'hBE35,4);
TASK_PP(16'hBE36,4);
TASK_PP(16'hBE37,4);
TASK_PP(16'hBE38,4);
TASK_PP(16'hBE39,4);
TASK_PP(16'hBE3A,4);
TASK_PP(16'hBE3B,4);
TASK_PP(16'hBE3C,4);
TASK_PP(16'hBE3D,4);
TASK_PP(16'hBE3E,4);
TASK_PP(16'hBE3F,4);
TASK_PP(16'hBE40,4);
TASK_PP(16'hBE41,4);
TASK_PP(16'hBE42,4);
TASK_PP(16'hBE43,4);
TASK_PP(16'hBE44,4);
TASK_PP(16'hBE45,4);
TASK_PP(16'hBE46,4);
TASK_PP(16'hBE47,4);
TASK_PP(16'hBE48,4);
TASK_PP(16'hBE49,4);
TASK_PP(16'hBE4A,4);
TASK_PP(16'hBE4B,4);
TASK_PP(16'hBE4C,4);
TASK_PP(16'hBE4D,4);
TASK_PP(16'hBE4E,4);
TASK_PP(16'hBE4F,4);
TASK_PP(16'hBE50,4);
TASK_PP(16'hBE51,4);
TASK_PP(16'hBE52,4);
TASK_PP(16'hBE53,4);
TASK_PP(16'hBE54,4);
TASK_PP(16'hBE55,4);
TASK_PP(16'hBE56,4);
TASK_PP(16'hBE57,4);
TASK_PP(16'hBE58,4);
TASK_PP(16'hBE59,4);
TASK_PP(16'hBE5A,4);
TASK_PP(16'hBE5B,4);
TASK_PP(16'hBE5C,4);
TASK_PP(16'hBE5D,4);
TASK_PP(16'hBE5E,4);
TASK_PP(16'hBE5F,4);
TASK_PP(16'hBE60,4);
TASK_PP(16'hBE61,4);
TASK_PP(16'hBE62,4);
TASK_PP(16'hBE63,4);
TASK_PP(16'hBE64,4);
TASK_PP(16'hBE65,4);
TASK_PP(16'hBE66,4);
TASK_PP(16'hBE67,4);
TASK_PP(16'hBE68,4);
TASK_PP(16'hBE69,4);
TASK_PP(16'hBE6A,4);
TASK_PP(16'hBE6B,4);
TASK_PP(16'hBE6C,4);
TASK_PP(16'hBE6D,4);
TASK_PP(16'hBE6E,4);
TASK_PP(16'hBE6F,4);
TASK_PP(16'hBE70,4);
TASK_PP(16'hBE71,4);
TASK_PP(16'hBE72,4);
TASK_PP(16'hBE73,4);
TASK_PP(16'hBE74,4);
TASK_PP(16'hBE75,4);
TASK_PP(16'hBE76,4);
TASK_PP(16'hBE77,4);
TASK_PP(16'hBE78,4);
TASK_PP(16'hBE79,4);
TASK_PP(16'hBE7A,4);
TASK_PP(16'hBE7B,4);
TASK_PP(16'hBE7C,4);
TASK_PP(16'hBE7D,4);
TASK_PP(16'hBE7E,4);
TASK_PP(16'hBE7F,4);
TASK_PP(16'hBE80,4);
TASK_PP(16'hBE81,4);
TASK_PP(16'hBE82,4);
TASK_PP(16'hBE83,4);
TASK_PP(16'hBE84,4);
TASK_PP(16'hBE85,4);
TASK_PP(16'hBE86,4);
TASK_PP(16'hBE87,4);
TASK_PP(16'hBE88,4);
TASK_PP(16'hBE89,4);
TASK_PP(16'hBE8A,4);
TASK_PP(16'hBE8B,4);
TASK_PP(16'hBE8C,4);
TASK_PP(16'hBE8D,4);
TASK_PP(16'hBE8E,4);
TASK_PP(16'hBE8F,4);
TASK_PP(16'hBE90,4);
TASK_PP(16'hBE91,4);
TASK_PP(16'hBE92,4);
TASK_PP(16'hBE93,4);
TASK_PP(16'hBE94,4);
TASK_PP(16'hBE95,4);
TASK_PP(16'hBE96,4);
TASK_PP(16'hBE97,4);
TASK_PP(16'hBE98,4);
TASK_PP(16'hBE99,4);
TASK_PP(16'hBE9A,4);
TASK_PP(16'hBE9B,4);
TASK_PP(16'hBE9C,4);
TASK_PP(16'hBE9D,4);
TASK_PP(16'hBE9E,4);
TASK_PP(16'hBE9F,4);
TASK_PP(16'hBEA0,4);
TASK_PP(16'hBEA1,4);
TASK_PP(16'hBEA2,4);
TASK_PP(16'hBEA3,4);
TASK_PP(16'hBEA4,4);
TASK_PP(16'hBEA5,4);
TASK_PP(16'hBEA6,4);
TASK_PP(16'hBEA7,4);
TASK_PP(16'hBEA8,4);
TASK_PP(16'hBEA9,4);
TASK_PP(16'hBEAA,4);
TASK_PP(16'hBEAB,4);
TASK_PP(16'hBEAC,4);
TASK_PP(16'hBEAD,4);
TASK_PP(16'hBEAE,4);
TASK_PP(16'hBEAF,4);
TASK_PP(16'hBEB0,4);
TASK_PP(16'hBEB1,4);
TASK_PP(16'hBEB2,4);
TASK_PP(16'hBEB3,4);
TASK_PP(16'hBEB4,4);
TASK_PP(16'hBEB5,4);
TASK_PP(16'hBEB6,4);
TASK_PP(16'hBEB7,4);
TASK_PP(16'hBEB8,4);
TASK_PP(16'hBEB9,4);
TASK_PP(16'hBEBA,4);
TASK_PP(16'hBEBB,4);
TASK_PP(16'hBEBC,4);
TASK_PP(16'hBEBD,4);
TASK_PP(16'hBEBE,4);
TASK_PP(16'hBEBF,4);
TASK_PP(16'hBEC0,4);
TASK_PP(16'hBEC1,4);
TASK_PP(16'hBEC2,4);
TASK_PP(16'hBEC3,4);
TASK_PP(16'hBEC4,4);
TASK_PP(16'hBEC5,4);
TASK_PP(16'hBEC6,4);
TASK_PP(16'hBEC7,4);
TASK_PP(16'hBEC8,4);
TASK_PP(16'hBEC9,4);
TASK_PP(16'hBECA,4);
TASK_PP(16'hBECB,4);
TASK_PP(16'hBECC,4);
TASK_PP(16'hBECD,4);
TASK_PP(16'hBECE,4);
TASK_PP(16'hBECF,4);
TASK_PP(16'hBED0,4);
TASK_PP(16'hBED1,4);
TASK_PP(16'hBED2,4);
TASK_PP(16'hBED3,4);
TASK_PP(16'hBED4,4);
TASK_PP(16'hBED5,4);
TASK_PP(16'hBED6,4);
TASK_PP(16'hBED7,4);
TASK_PP(16'hBED8,4);
TASK_PP(16'hBED9,4);
TASK_PP(16'hBEDA,4);
TASK_PP(16'hBEDB,4);
TASK_PP(16'hBEDC,4);
TASK_PP(16'hBEDD,4);
TASK_PP(16'hBEDE,4);
TASK_PP(16'hBEDF,4);
TASK_PP(16'hBEE0,4);
TASK_PP(16'hBEE1,4);
TASK_PP(16'hBEE2,4);
TASK_PP(16'hBEE3,4);
TASK_PP(16'hBEE4,4);
TASK_PP(16'hBEE5,4);
TASK_PP(16'hBEE6,4);
TASK_PP(16'hBEE7,4);
TASK_PP(16'hBEE8,4);
TASK_PP(16'hBEE9,4);
TASK_PP(16'hBEEA,4);
TASK_PP(16'hBEEB,4);
TASK_PP(16'hBEEC,4);
TASK_PP(16'hBEED,4);
TASK_PP(16'hBEEE,4);
TASK_PP(16'hBEEF,4);
TASK_PP(16'hBEF0,4);
TASK_PP(16'hBEF1,4);
TASK_PP(16'hBEF2,4);
TASK_PP(16'hBEF3,4);
TASK_PP(16'hBEF4,4);
TASK_PP(16'hBEF5,4);
TASK_PP(16'hBEF6,4);
TASK_PP(16'hBEF7,4);
TASK_PP(16'hBEF8,4);
TASK_PP(16'hBEF9,4);
TASK_PP(16'hBEFA,4);
TASK_PP(16'hBEFB,4);
TASK_PP(16'hBEFC,4);
TASK_PP(16'hBEFD,4);
TASK_PP(16'hBEFE,4);
TASK_PP(16'hBEFF,4);
TASK_PP(16'hBF00,4);
TASK_PP(16'hBF01,4);
TASK_PP(16'hBF02,4);
TASK_PP(16'hBF03,4);
TASK_PP(16'hBF04,4);
TASK_PP(16'hBF05,4);
TASK_PP(16'hBF06,4);
TASK_PP(16'hBF07,4);
TASK_PP(16'hBF08,4);
TASK_PP(16'hBF09,4);
TASK_PP(16'hBF0A,4);
TASK_PP(16'hBF0B,4);
TASK_PP(16'hBF0C,4);
TASK_PP(16'hBF0D,4);
TASK_PP(16'hBF0E,4);
TASK_PP(16'hBF0F,4);
TASK_PP(16'hBF10,4);
TASK_PP(16'hBF11,4);
TASK_PP(16'hBF12,4);
TASK_PP(16'hBF13,4);
TASK_PP(16'hBF14,4);
TASK_PP(16'hBF15,4);
TASK_PP(16'hBF16,4);
TASK_PP(16'hBF17,4);
TASK_PP(16'hBF18,4);
TASK_PP(16'hBF19,4);
TASK_PP(16'hBF1A,4);
TASK_PP(16'hBF1B,4);
TASK_PP(16'hBF1C,4);
TASK_PP(16'hBF1D,4);
TASK_PP(16'hBF1E,4);
TASK_PP(16'hBF1F,4);
TASK_PP(16'hBF20,4);
TASK_PP(16'hBF21,4);
TASK_PP(16'hBF22,4);
TASK_PP(16'hBF23,4);
TASK_PP(16'hBF24,4);
TASK_PP(16'hBF25,4);
TASK_PP(16'hBF26,4);
TASK_PP(16'hBF27,4);
TASK_PP(16'hBF28,4);
TASK_PP(16'hBF29,4);
TASK_PP(16'hBF2A,4);
TASK_PP(16'hBF2B,4);
TASK_PP(16'hBF2C,4);
TASK_PP(16'hBF2D,4);
TASK_PP(16'hBF2E,4);
TASK_PP(16'hBF2F,4);
TASK_PP(16'hBF30,4);
TASK_PP(16'hBF31,4);
TASK_PP(16'hBF32,4);
TASK_PP(16'hBF33,4);
TASK_PP(16'hBF34,4);
TASK_PP(16'hBF35,4);
TASK_PP(16'hBF36,4);
TASK_PP(16'hBF37,4);
TASK_PP(16'hBF38,4);
TASK_PP(16'hBF39,4);
TASK_PP(16'hBF3A,4);
TASK_PP(16'hBF3B,4);
TASK_PP(16'hBF3C,4);
TASK_PP(16'hBF3D,4);
TASK_PP(16'hBF3E,4);
TASK_PP(16'hBF3F,4);
TASK_PP(16'hBF40,4);
TASK_PP(16'hBF41,4);
TASK_PP(16'hBF42,4);
TASK_PP(16'hBF43,4);
TASK_PP(16'hBF44,4);
TASK_PP(16'hBF45,4);
TASK_PP(16'hBF46,4);
TASK_PP(16'hBF47,4);
TASK_PP(16'hBF48,4);
TASK_PP(16'hBF49,4);
TASK_PP(16'hBF4A,4);
TASK_PP(16'hBF4B,4);
TASK_PP(16'hBF4C,4);
TASK_PP(16'hBF4D,4);
TASK_PP(16'hBF4E,4);
TASK_PP(16'hBF4F,4);
TASK_PP(16'hBF50,4);
TASK_PP(16'hBF51,4);
TASK_PP(16'hBF52,4);
TASK_PP(16'hBF53,4);
TASK_PP(16'hBF54,4);
TASK_PP(16'hBF55,4);
TASK_PP(16'hBF56,4);
TASK_PP(16'hBF57,4);
TASK_PP(16'hBF58,4);
TASK_PP(16'hBF59,4);
TASK_PP(16'hBF5A,4);
TASK_PP(16'hBF5B,4);
TASK_PP(16'hBF5C,4);
TASK_PP(16'hBF5D,4);
TASK_PP(16'hBF5E,4);
TASK_PP(16'hBF5F,4);
TASK_PP(16'hBF60,4);
TASK_PP(16'hBF61,4);
TASK_PP(16'hBF62,4);
TASK_PP(16'hBF63,4);
TASK_PP(16'hBF64,4);
TASK_PP(16'hBF65,4);
TASK_PP(16'hBF66,4);
TASK_PP(16'hBF67,4);
TASK_PP(16'hBF68,4);
TASK_PP(16'hBF69,4);
TASK_PP(16'hBF6A,4);
TASK_PP(16'hBF6B,4);
TASK_PP(16'hBF6C,4);
TASK_PP(16'hBF6D,4);
TASK_PP(16'hBF6E,4);
TASK_PP(16'hBF6F,4);
TASK_PP(16'hBF70,4);
TASK_PP(16'hBF71,4);
TASK_PP(16'hBF72,4);
TASK_PP(16'hBF73,4);
TASK_PP(16'hBF74,4);
TASK_PP(16'hBF75,4);
TASK_PP(16'hBF76,4);
TASK_PP(16'hBF77,4);
TASK_PP(16'hBF78,4);
TASK_PP(16'hBF79,4);
TASK_PP(16'hBF7A,4);
TASK_PP(16'hBF7B,4);
TASK_PP(16'hBF7C,4);
TASK_PP(16'hBF7D,4);
TASK_PP(16'hBF7E,4);
TASK_PP(16'hBF7F,4);
TASK_PP(16'hBF80,4);
TASK_PP(16'hBF81,4);
TASK_PP(16'hBF82,4);
TASK_PP(16'hBF83,4);
TASK_PP(16'hBF84,4);
TASK_PP(16'hBF85,4);
TASK_PP(16'hBF86,4);
TASK_PP(16'hBF87,4);
TASK_PP(16'hBF88,4);
TASK_PP(16'hBF89,4);
TASK_PP(16'hBF8A,4);
TASK_PP(16'hBF8B,4);
TASK_PP(16'hBF8C,4);
TASK_PP(16'hBF8D,4);
TASK_PP(16'hBF8E,4);
TASK_PP(16'hBF8F,4);
TASK_PP(16'hBF90,4);
TASK_PP(16'hBF91,4);
TASK_PP(16'hBF92,4);
TASK_PP(16'hBF93,4);
TASK_PP(16'hBF94,4);
TASK_PP(16'hBF95,4);
TASK_PP(16'hBF96,4);
TASK_PP(16'hBF97,4);
TASK_PP(16'hBF98,4);
TASK_PP(16'hBF99,4);
TASK_PP(16'hBF9A,4);
TASK_PP(16'hBF9B,4);
TASK_PP(16'hBF9C,4);
TASK_PP(16'hBF9D,4);
TASK_PP(16'hBF9E,4);
TASK_PP(16'hBF9F,4);
TASK_PP(16'hBFA0,4);
TASK_PP(16'hBFA1,4);
TASK_PP(16'hBFA2,4);
TASK_PP(16'hBFA3,4);
TASK_PP(16'hBFA4,4);
TASK_PP(16'hBFA5,4);
TASK_PP(16'hBFA6,4);
TASK_PP(16'hBFA7,4);
TASK_PP(16'hBFA8,4);
TASK_PP(16'hBFA9,4);
TASK_PP(16'hBFAA,4);
TASK_PP(16'hBFAB,4);
TASK_PP(16'hBFAC,4);
TASK_PP(16'hBFAD,4);
TASK_PP(16'hBFAE,4);
TASK_PP(16'hBFAF,4);
TASK_PP(16'hBFB0,4);
TASK_PP(16'hBFB1,4);
TASK_PP(16'hBFB2,4);
TASK_PP(16'hBFB3,4);
TASK_PP(16'hBFB4,4);
TASK_PP(16'hBFB5,4);
TASK_PP(16'hBFB6,4);
TASK_PP(16'hBFB7,4);
TASK_PP(16'hBFB8,4);
TASK_PP(16'hBFB9,4);
TASK_PP(16'hBFBA,4);
TASK_PP(16'hBFBB,4);
TASK_PP(16'hBFBC,4);
TASK_PP(16'hBFBD,4);
TASK_PP(16'hBFBE,4);
TASK_PP(16'hBFBF,4);
TASK_PP(16'hBFC0,4);
TASK_PP(16'hBFC1,4);
TASK_PP(16'hBFC2,4);
TASK_PP(16'hBFC3,4);
TASK_PP(16'hBFC4,4);
TASK_PP(16'hBFC5,4);
TASK_PP(16'hBFC6,4);
TASK_PP(16'hBFC7,4);
TASK_PP(16'hBFC8,4);
TASK_PP(16'hBFC9,4);
TASK_PP(16'hBFCA,4);
TASK_PP(16'hBFCB,4);
TASK_PP(16'hBFCC,4);
TASK_PP(16'hBFCD,4);
TASK_PP(16'hBFCE,4);
TASK_PP(16'hBFCF,4);
TASK_PP(16'hBFD0,4);
TASK_PP(16'hBFD1,4);
TASK_PP(16'hBFD2,4);
TASK_PP(16'hBFD3,4);
TASK_PP(16'hBFD4,4);
TASK_PP(16'hBFD5,4);
TASK_PP(16'hBFD6,4);
TASK_PP(16'hBFD7,4);
TASK_PP(16'hBFD8,4);
TASK_PP(16'hBFD9,4);
TASK_PP(16'hBFDA,4);
TASK_PP(16'hBFDB,4);
TASK_PP(16'hBFDC,4);
TASK_PP(16'hBFDD,4);
TASK_PP(16'hBFDE,4);
TASK_PP(16'hBFDF,4);
TASK_PP(16'hBFE0,4);
TASK_PP(16'hBFE1,4);
TASK_PP(16'hBFE2,4);
TASK_PP(16'hBFE3,4);
TASK_PP(16'hBFE4,4);
TASK_PP(16'hBFE5,4);
TASK_PP(16'hBFE6,4);
TASK_PP(16'hBFE7,4);
TASK_PP(16'hBFE8,4);
TASK_PP(16'hBFE9,4);
TASK_PP(16'hBFEA,4);
TASK_PP(16'hBFEB,4);
TASK_PP(16'hBFEC,4);
TASK_PP(16'hBFED,4);
TASK_PP(16'hBFEE,4);
TASK_PP(16'hBFEF,4);
TASK_PP(16'hBFF0,4);
TASK_PP(16'hBFF1,4);
TASK_PP(16'hBFF2,4);
TASK_PP(16'hBFF3,4);
TASK_PP(16'hBFF4,4);
TASK_PP(16'hBFF5,4);
TASK_PP(16'hBFF6,4);
TASK_PP(16'hBFF7,4);
TASK_PP(16'hBFF8,4);
TASK_PP(16'hBFF9,4);
TASK_PP(16'hBFFA,4);
TASK_PP(16'hBFFB,4);
TASK_PP(16'hBFFC,4);
TASK_PP(16'hBFFD,4);
TASK_PP(16'hBFFE,4);
TASK_PP(16'hBFFF,4);
TASK_PP(16'hC000,4);
TASK_PP(16'hC001,4);
TASK_PP(16'hC002,4);
TASK_PP(16'hC003,4);
TASK_PP(16'hC004,4);
TASK_PP(16'hC005,4);
TASK_PP(16'hC006,4);
TASK_PP(16'hC007,4);
TASK_PP(16'hC008,4);
TASK_PP(16'hC009,4);
TASK_PP(16'hC00A,4);
TASK_PP(16'hC00B,4);
TASK_PP(16'hC00C,4);
TASK_PP(16'hC00D,4);
TASK_PP(16'hC00E,4);
TASK_PP(16'hC00F,4);
TASK_PP(16'hC010,4);
TASK_PP(16'hC011,4);
TASK_PP(16'hC012,4);
TASK_PP(16'hC013,4);
TASK_PP(16'hC014,4);
TASK_PP(16'hC015,4);
TASK_PP(16'hC016,4);
TASK_PP(16'hC017,4);
TASK_PP(16'hC018,4);
TASK_PP(16'hC019,4);
TASK_PP(16'hC01A,4);
TASK_PP(16'hC01B,4);
TASK_PP(16'hC01C,4);
TASK_PP(16'hC01D,4);
TASK_PP(16'hC01E,4);
TASK_PP(16'hC01F,4);
TASK_PP(16'hC020,4);
TASK_PP(16'hC021,4);
TASK_PP(16'hC022,4);
TASK_PP(16'hC023,4);
TASK_PP(16'hC024,4);
TASK_PP(16'hC025,4);
TASK_PP(16'hC026,4);
TASK_PP(16'hC027,4);
TASK_PP(16'hC028,4);
TASK_PP(16'hC029,4);
TASK_PP(16'hC02A,4);
TASK_PP(16'hC02B,4);
TASK_PP(16'hC02C,4);
TASK_PP(16'hC02D,4);
TASK_PP(16'hC02E,4);
TASK_PP(16'hC02F,4);
TASK_PP(16'hC030,4);
TASK_PP(16'hC031,4);
TASK_PP(16'hC032,4);
TASK_PP(16'hC033,4);
TASK_PP(16'hC034,4);
TASK_PP(16'hC035,4);
TASK_PP(16'hC036,4);
TASK_PP(16'hC037,4);
TASK_PP(16'hC038,4);
TASK_PP(16'hC039,4);
TASK_PP(16'hC03A,4);
TASK_PP(16'hC03B,4);
TASK_PP(16'hC03C,4);
TASK_PP(16'hC03D,4);
TASK_PP(16'hC03E,4);
TASK_PP(16'hC03F,4);
TASK_PP(16'hC040,4);
TASK_PP(16'hC041,4);
TASK_PP(16'hC042,4);
TASK_PP(16'hC043,4);
TASK_PP(16'hC044,4);
TASK_PP(16'hC045,4);
TASK_PP(16'hC046,4);
TASK_PP(16'hC047,4);
TASK_PP(16'hC048,4);
TASK_PP(16'hC049,4);
TASK_PP(16'hC04A,4);
TASK_PP(16'hC04B,4);
TASK_PP(16'hC04C,4);
TASK_PP(16'hC04D,4);
TASK_PP(16'hC04E,4);
TASK_PP(16'hC04F,4);
TASK_PP(16'hC050,4);
TASK_PP(16'hC051,4);
TASK_PP(16'hC052,4);
TASK_PP(16'hC053,4);
TASK_PP(16'hC054,4);
TASK_PP(16'hC055,4);
TASK_PP(16'hC056,4);
TASK_PP(16'hC057,4);
TASK_PP(16'hC058,4);
TASK_PP(16'hC059,4);
TASK_PP(16'hC05A,4);
TASK_PP(16'hC05B,4);
TASK_PP(16'hC05C,4);
TASK_PP(16'hC05D,4);
TASK_PP(16'hC05E,4);
TASK_PP(16'hC05F,4);
TASK_PP(16'hC060,4);
TASK_PP(16'hC061,4);
TASK_PP(16'hC062,4);
TASK_PP(16'hC063,4);
TASK_PP(16'hC064,4);
TASK_PP(16'hC065,4);
TASK_PP(16'hC066,4);
TASK_PP(16'hC067,4);
TASK_PP(16'hC068,4);
TASK_PP(16'hC069,4);
TASK_PP(16'hC06A,4);
TASK_PP(16'hC06B,4);
TASK_PP(16'hC06C,4);
TASK_PP(16'hC06D,4);
TASK_PP(16'hC06E,4);
TASK_PP(16'hC06F,4);
TASK_PP(16'hC070,4);
TASK_PP(16'hC071,4);
TASK_PP(16'hC072,4);
TASK_PP(16'hC073,4);
TASK_PP(16'hC074,4);
TASK_PP(16'hC075,4);
TASK_PP(16'hC076,4);
TASK_PP(16'hC077,4);
TASK_PP(16'hC078,4);
TASK_PP(16'hC079,4);
TASK_PP(16'hC07A,4);
TASK_PP(16'hC07B,4);
TASK_PP(16'hC07C,4);
TASK_PP(16'hC07D,4);
TASK_PP(16'hC07E,4);
TASK_PP(16'hC07F,4);
TASK_PP(16'hC080,4);
TASK_PP(16'hC081,4);
TASK_PP(16'hC082,4);
TASK_PP(16'hC083,4);
TASK_PP(16'hC084,4);
TASK_PP(16'hC085,4);
TASK_PP(16'hC086,4);
TASK_PP(16'hC087,4);
TASK_PP(16'hC088,4);
TASK_PP(16'hC089,4);
TASK_PP(16'hC08A,4);
TASK_PP(16'hC08B,4);
TASK_PP(16'hC08C,4);
TASK_PP(16'hC08D,4);
TASK_PP(16'hC08E,4);
TASK_PP(16'hC08F,4);
TASK_PP(16'hC090,4);
TASK_PP(16'hC091,4);
TASK_PP(16'hC092,4);
TASK_PP(16'hC093,4);
TASK_PP(16'hC094,4);
TASK_PP(16'hC095,4);
TASK_PP(16'hC096,4);
TASK_PP(16'hC097,4);
TASK_PP(16'hC098,4);
TASK_PP(16'hC099,4);
TASK_PP(16'hC09A,4);
TASK_PP(16'hC09B,4);
TASK_PP(16'hC09C,4);
TASK_PP(16'hC09D,4);
TASK_PP(16'hC09E,4);
TASK_PP(16'hC09F,4);
TASK_PP(16'hC0A0,4);
TASK_PP(16'hC0A1,4);
TASK_PP(16'hC0A2,4);
TASK_PP(16'hC0A3,4);
TASK_PP(16'hC0A4,4);
TASK_PP(16'hC0A5,4);
TASK_PP(16'hC0A6,4);
TASK_PP(16'hC0A7,4);
TASK_PP(16'hC0A8,4);
TASK_PP(16'hC0A9,4);
TASK_PP(16'hC0AA,4);
TASK_PP(16'hC0AB,4);
TASK_PP(16'hC0AC,4);
TASK_PP(16'hC0AD,4);
TASK_PP(16'hC0AE,4);
TASK_PP(16'hC0AF,4);
TASK_PP(16'hC0B0,4);
TASK_PP(16'hC0B1,4);
TASK_PP(16'hC0B2,4);
TASK_PP(16'hC0B3,4);
TASK_PP(16'hC0B4,4);
TASK_PP(16'hC0B5,4);
TASK_PP(16'hC0B6,4);
TASK_PP(16'hC0B7,4);
TASK_PP(16'hC0B8,4);
TASK_PP(16'hC0B9,4);
TASK_PP(16'hC0BA,4);
TASK_PP(16'hC0BB,4);
TASK_PP(16'hC0BC,4);
TASK_PP(16'hC0BD,4);
TASK_PP(16'hC0BE,4);
TASK_PP(16'hC0BF,4);
TASK_PP(16'hC0C0,4);
TASK_PP(16'hC0C1,4);
TASK_PP(16'hC0C2,4);
TASK_PP(16'hC0C3,4);
TASK_PP(16'hC0C4,4);
TASK_PP(16'hC0C5,4);
TASK_PP(16'hC0C6,4);
TASK_PP(16'hC0C7,4);
TASK_PP(16'hC0C8,4);
TASK_PP(16'hC0C9,4);
TASK_PP(16'hC0CA,4);
TASK_PP(16'hC0CB,4);
TASK_PP(16'hC0CC,4);
TASK_PP(16'hC0CD,4);
TASK_PP(16'hC0CE,4);
TASK_PP(16'hC0CF,4);
TASK_PP(16'hC0D0,4);
TASK_PP(16'hC0D1,4);
TASK_PP(16'hC0D2,4);
TASK_PP(16'hC0D3,4);
TASK_PP(16'hC0D4,4);
TASK_PP(16'hC0D5,4);
TASK_PP(16'hC0D6,4);
TASK_PP(16'hC0D7,4);
TASK_PP(16'hC0D8,4);
TASK_PP(16'hC0D9,4);
TASK_PP(16'hC0DA,4);
TASK_PP(16'hC0DB,4);
TASK_PP(16'hC0DC,4);
TASK_PP(16'hC0DD,4);
TASK_PP(16'hC0DE,4);
TASK_PP(16'hC0DF,4);
TASK_PP(16'hC0E0,4);
TASK_PP(16'hC0E1,4);
TASK_PP(16'hC0E2,4);
TASK_PP(16'hC0E3,4);
TASK_PP(16'hC0E4,4);
TASK_PP(16'hC0E5,4);
TASK_PP(16'hC0E6,4);
TASK_PP(16'hC0E7,4);
TASK_PP(16'hC0E8,4);
TASK_PP(16'hC0E9,4);
TASK_PP(16'hC0EA,4);
TASK_PP(16'hC0EB,4);
TASK_PP(16'hC0EC,4);
TASK_PP(16'hC0ED,4);
TASK_PP(16'hC0EE,4);
TASK_PP(16'hC0EF,4);
TASK_PP(16'hC0F0,4);
TASK_PP(16'hC0F1,4);
TASK_PP(16'hC0F2,4);
TASK_PP(16'hC0F3,4);
TASK_PP(16'hC0F4,4);
TASK_PP(16'hC0F5,4);
TASK_PP(16'hC0F6,4);
TASK_PP(16'hC0F7,4);
TASK_PP(16'hC0F8,4);
TASK_PP(16'hC0F9,4);
TASK_PP(16'hC0FA,4);
TASK_PP(16'hC0FB,4);
TASK_PP(16'hC0FC,4);
TASK_PP(16'hC0FD,4);
TASK_PP(16'hC0FE,4);
TASK_PP(16'hC0FF,4);
TASK_PP(16'hC100,4);
TASK_PP(16'hC101,4);
TASK_PP(16'hC102,4);
TASK_PP(16'hC103,4);
TASK_PP(16'hC104,4);
TASK_PP(16'hC105,4);
TASK_PP(16'hC106,4);
TASK_PP(16'hC107,4);
TASK_PP(16'hC108,4);
TASK_PP(16'hC109,4);
TASK_PP(16'hC10A,4);
TASK_PP(16'hC10B,4);
TASK_PP(16'hC10C,4);
TASK_PP(16'hC10D,4);
TASK_PP(16'hC10E,4);
TASK_PP(16'hC10F,4);
TASK_PP(16'hC110,4);
TASK_PP(16'hC111,4);
TASK_PP(16'hC112,4);
TASK_PP(16'hC113,4);
TASK_PP(16'hC114,4);
TASK_PP(16'hC115,4);
TASK_PP(16'hC116,4);
TASK_PP(16'hC117,4);
TASK_PP(16'hC118,4);
TASK_PP(16'hC119,4);
TASK_PP(16'hC11A,4);
TASK_PP(16'hC11B,4);
TASK_PP(16'hC11C,4);
TASK_PP(16'hC11D,4);
TASK_PP(16'hC11E,4);
TASK_PP(16'hC11F,4);
TASK_PP(16'hC120,4);
TASK_PP(16'hC121,4);
TASK_PP(16'hC122,4);
TASK_PP(16'hC123,4);
TASK_PP(16'hC124,4);
TASK_PP(16'hC125,4);
TASK_PP(16'hC126,4);
TASK_PP(16'hC127,4);
TASK_PP(16'hC128,4);
TASK_PP(16'hC129,4);
TASK_PP(16'hC12A,4);
TASK_PP(16'hC12B,4);
TASK_PP(16'hC12C,4);
TASK_PP(16'hC12D,4);
TASK_PP(16'hC12E,4);
TASK_PP(16'hC12F,4);
TASK_PP(16'hC130,4);
TASK_PP(16'hC131,4);
TASK_PP(16'hC132,4);
TASK_PP(16'hC133,4);
TASK_PP(16'hC134,4);
TASK_PP(16'hC135,4);
TASK_PP(16'hC136,4);
TASK_PP(16'hC137,4);
TASK_PP(16'hC138,4);
TASK_PP(16'hC139,4);
TASK_PP(16'hC13A,4);
TASK_PP(16'hC13B,4);
TASK_PP(16'hC13C,4);
TASK_PP(16'hC13D,4);
TASK_PP(16'hC13E,4);
TASK_PP(16'hC13F,4);
TASK_PP(16'hC140,4);
TASK_PP(16'hC141,4);
TASK_PP(16'hC142,4);
TASK_PP(16'hC143,4);
TASK_PP(16'hC144,4);
TASK_PP(16'hC145,4);
TASK_PP(16'hC146,4);
TASK_PP(16'hC147,4);
TASK_PP(16'hC148,4);
TASK_PP(16'hC149,4);
TASK_PP(16'hC14A,4);
TASK_PP(16'hC14B,4);
TASK_PP(16'hC14C,4);
TASK_PP(16'hC14D,4);
TASK_PP(16'hC14E,4);
TASK_PP(16'hC14F,4);
TASK_PP(16'hC150,4);
TASK_PP(16'hC151,4);
TASK_PP(16'hC152,4);
TASK_PP(16'hC153,4);
TASK_PP(16'hC154,4);
TASK_PP(16'hC155,4);
TASK_PP(16'hC156,4);
TASK_PP(16'hC157,4);
TASK_PP(16'hC158,4);
TASK_PP(16'hC159,4);
TASK_PP(16'hC15A,4);
TASK_PP(16'hC15B,4);
TASK_PP(16'hC15C,4);
TASK_PP(16'hC15D,4);
TASK_PP(16'hC15E,4);
TASK_PP(16'hC15F,4);
TASK_PP(16'hC160,4);
TASK_PP(16'hC161,4);
TASK_PP(16'hC162,4);
TASK_PP(16'hC163,4);
TASK_PP(16'hC164,4);
TASK_PP(16'hC165,4);
TASK_PP(16'hC166,4);
TASK_PP(16'hC167,4);
TASK_PP(16'hC168,4);
TASK_PP(16'hC169,4);
TASK_PP(16'hC16A,4);
TASK_PP(16'hC16B,4);
TASK_PP(16'hC16C,4);
TASK_PP(16'hC16D,4);
TASK_PP(16'hC16E,4);
TASK_PP(16'hC16F,4);
TASK_PP(16'hC170,4);
TASK_PP(16'hC171,4);
TASK_PP(16'hC172,4);
TASK_PP(16'hC173,4);
TASK_PP(16'hC174,4);
TASK_PP(16'hC175,4);
TASK_PP(16'hC176,4);
TASK_PP(16'hC177,4);
TASK_PP(16'hC178,4);
TASK_PP(16'hC179,4);
TASK_PP(16'hC17A,4);
TASK_PP(16'hC17B,4);
TASK_PP(16'hC17C,4);
TASK_PP(16'hC17D,4);
TASK_PP(16'hC17E,4);
TASK_PP(16'hC17F,4);
TASK_PP(16'hC180,4);
TASK_PP(16'hC181,4);
TASK_PP(16'hC182,4);
TASK_PP(16'hC183,4);
TASK_PP(16'hC184,4);
TASK_PP(16'hC185,4);
TASK_PP(16'hC186,4);
TASK_PP(16'hC187,4);
TASK_PP(16'hC188,4);
TASK_PP(16'hC189,4);
TASK_PP(16'hC18A,4);
TASK_PP(16'hC18B,4);
TASK_PP(16'hC18C,4);
TASK_PP(16'hC18D,4);
TASK_PP(16'hC18E,4);
TASK_PP(16'hC18F,4);
TASK_PP(16'hC190,4);
TASK_PP(16'hC191,4);
TASK_PP(16'hC192,4);
TASK_PP(16'hC193,4);
TASK_PP(16'hC194,4);
TASK_PP(16'hC195,4);
TASK_PP(16'hC196,4);
TASK_PP(16'hC197,4);
TASK_PP(16'hC198,4);
TASK_PP(16'hC199,4);
TASK_PP(16'hC19A,4);
TASK_PP(16'hC19B,4);
TASK_PP(16'hC19C,4);
TASK_PP(16'hC19D,4);
TASK_PP(16'hC19E,4);
TASK_PP(16'hC19F,4);
TASK_PP(16'hC1A0,4);
TASK_PP(16'hC1A1,4);
TASK_PP(16'hC1A2,4);
TASK_PP(16'hC1A3,4);
TASK_PP(16'hC1A4,4);
TASK_PP(16'hC1A5,4);
TASK_PP(16'hC1A6,4);
TASK_PP(16'hC1A7,4);
TASK_PP(16'hC1A8,4);
TASK_PP(16'hC1A9,4);
TASK_PP(16'hC1AA,4);
TASK_PP(16'hC1AB,4);
TASK_PP(16'hC1AC,4);
TASK_PP(16'hC1AD,4);
TASK_PP(16'hC1AE,4);
TASK_PP(16'hC1AF,4);
TASK_PP(16'hC1B0,4);
TASK_PP(16'hC1B1,4);
TASK_PP(16'hC1B2,4);
TASK_PP(16'hC1B3,4);
TASK_PP(16'hC1B4,4);
TASK_PP(16'hC1B5,4);
TASK_PP(16'hC1B6,4);
TASK_PP(16'hC1B7,4);
TASK_PP(16'hC1B8,4);
TASK_PP(16'hC1B9,4);
TASK_PP(16'hC1BA,4);
TASK_PP(16'hC1BB,4);
TASK_PP(16'hC1BC,4);
TASK_PP(16'hC1BD,4);
TASK_PP(16'hC1BE,4);
TASK_PP(16'hC1BF,4);
TASK_PP(16'hC1C0,4);
TASK_PP(16'hC1C1,4);
TASK_PP(16'hC1C2,4);
TASK_PP(16'hC1C3,4);
TASK_PP(16'hC1C4,4);
TASK_PP(16'hC1C5,4);
TASK_PP(16'hC1C6,4);
TASK_PP(16'hC1C7,4);
TASK_PP(16'hC1C8,4);
TASK_PP(16'hC1C9,4);
TASK_PP(16'hC1CA,4);
TASK_PP(16'hC1CB,4);
TASK_PP(16'hC1CC,4);
TASK_PP(16'hC1CD,4);
TASK_PP(16'hC1CE,4);
TASK_PP(16'hC1CF,4);
TASK_PP(16'hC1D0,4);
TASK_PP(16'hC1D1,4);
TASK_PP(16'hC1D2,4);
TASK_PP(16'hC1D3,4);
TASK_PP(16'hC1D4,4);
TASK_PP(16'hC1D5,4);
TASK_PP(16'hC1D6,4);
TASK_PP(16'hC1D7,4);
TASK_PP(16'hC1D8,4);
TASK_PP(16'hC1D9,4);
TASK_PP(16'hC1DA,4);
TASK_PP(16'hC1DB,4);
TASK_PP(16'hC1DC,4);
TASK_PP(16'hC1DD,4);
TASK_PP(16'hC1DE,4);
TASK_PP(16'hC1DF,4);
TASK_PP(16'hC1E0,4);
TASK_PP(16'hC1E1,4);
TASK_PP(16'hC1E2,4);
TASK_PP(16'hC1E3,4);
TASK_PP(16'hC1E4,4);
TASK_PP(16'hC1E5,4);
TASK_PP(16'hC1E6,4);
TASK_PP(16'hC1E7,4);
TASK_PP(16'hC1E8,4);
TASK_PP(16'hC1E9,4);
TASK_PP(16'hC1EA,4);
TASK_PP(16'hC1EB,4);
TASK_PP(16'hC1EC,4);
TASK_PP(16'hC1ED,4);
TASK_PP(16'hC1EE,4);
TASK_PP(16'hC1EF,4);
TASK_PP(16'hC1F0,4);
TASK_PP(16'hC1F1,4);
TASK_PP(16'hC1F2,4);
TASK_PP(16'hC1F3,4);
TASK_PP(16'hC1F4,4);
TASK_PP(16'hC1F5,4);
TASK_PP(16'hC1F6,4);
TASK_PP(16'hC1F7,4);
TASK_PP(16'hC1F8,4);
TASK_PP(16'hC1F9,4);
TASK_PP(16'hC1FA,4);
TASK_PP(16'hC1FB,4);
TASK_PP(16'hC1FC,4);
TASK_PP(16'hC1FD,4);
TASK_PP(16'hC1FE,4);
TASK_PP(16'hC1FF,4);
TASK_PP(16'hC200,4);
TASK_PP(16'hC201,4);
TASK_PP(16'hC202,4);
TASK_PP(16'hC203,4);
TASK_PP(16'hC204,4);
TASK_PP(16'hC205,4);
TASK_PP(16'hC206,4);
TASK_PP(16'hC207,4);
TASK_PP(16'hC208,4);
TASK_PP(16'hC209,4);
TASK_PP(16'hC20A,4);
TASK_PP(16'hC20B,4);
TASK_PP(16'hC20C,4);
TASK_PP(16'hC20D,4);
TASK_PP(16'hC20E,4);
TASK_PP(16'hC20F,4);
TASK_PP(16'hC210,4);
TASK_PP(16'hC211,4);
TASK_PP(16'hC212,4);
TASK_PP(16'hC213,4);
TASK_PP(16'hC214,4);
TASK_PP(16'hC215,4);
TASK_PP(16'hC216,4);
TASK_PP(16'hC217,4);
TASK_PP(16'hC218,4);
TASK_PP(16'hC219,4);
TASK_PP(16'hC21A,4);
TASK_PP(16'hC21B,4);
TASK_PP(16'hC21C,4);
TASK_PP(16'hC21D,4);
TASK_PP(16'hC21E,4);
TASK_PP(16'hC21F,4);
TASK_PP(16'hC220,4);
TASK_PP(16'hC221,4);
TASK_PP(16'hC222,4);
TASK_PP(16'hC223,4);
TASK_PP(16'hC224,4);
TASK_PP(16'hC225,4);
TASK_PP(16'hC226,4);
TASK_PP(16'hC227,4);
TASK_PP(16'hC228,4);
TASK_PP(16'hC229,4);
TASK_PP(16'hC22A,4);
TASK_PP(16'hC22B,4);
TASK_PP(16'hC22C,4);
TASK_PP(16'hC22D,4);
TASK_PP(16'hC22E,4);
TASK_PP(16'hC22F,4);
TASK_PP(16'hC230,4);
TASK_PP(16'hC231,4);
TASK_PP(16'hC232,4);
TASK_PP(16'hC233,4);
TASK_PP(16'hC234,4);
TASK_PP(16'hC235,4);
TASK_PP(16'hC236,4);
TASK_PP(16'hC237,4);
TASK_PP(16'hC238,4);
TASK_PP(16'hC239,4);
TASK_PP(16'hC23A,4);
TASK_PP(16'hC23B,4);
TASK_PP(16'hC23C,4);
TASK_PP(16'hC23D,4);
TASK_PP(16'hC23E,4);
TASK_PP(16'hC23F,4);
TASK_PP(16'hC240,4);
TASK_PP(16'hC241,4);
TASK_PP(16'hC242,4);
TASK_PP(16'hC243,4);
TASK_PP(16'hC244,4);
TASK_PP(16'hC245,4);
TASK_PP(16'hC246,4);
TASK_PP(16'hC247,4);
TASK_PP(16'hC248,4);
TASK_PP(16'hC249,4);
TASK_PP(16'hC24A,4);
TASK_PP(16'hC24B,4);
TASK_PP(16'hC24C,4);
TASK_PP(16'hC24D,4);
TASK_PP(16'hC24E,4);
TASK_PP(16'hC24F,4);
TASK_PP(16'hC250,4);
TASK_PP(16'hC251,4);
TASK_PP(16'hC252,4);
TASK_PP(16'hC253,4);
TASK_PP(16'hC254,4);
TASK_PP(16'hC255,4);
TASK_PP(16'hC256,4);
TASK_PP(16'hC257,4);
TASK_PP(16'hC258,4);
TASK_PP(16'hC259,4);
TASK_PP(16'hC25A,4);
TASK_PP(16'hC25B,4);
TASK_PP(16'hC25C,4);
TASK_PP(16'hC25D,4);
TASK_PP(16'hC25E,4);
TASK_PP(16'hC25F,4);
TASK_PP(16'hC260,4);
TASK_PP(16'hC261,4);
TASK_PP(16'hC262,4);
TASK_PP(16'hC263,4);
TASK_PP(16'hC264,4);
TASK_PP(16'hC265,4);
TASK_PP(16'hC266,4);
TASK_PP(16'hC267,4);
TASK_PP(16'hC268,4);
TASK_PP(16'hC269,4);
TASK_PP(16'hC26A,4);
TASK_PP(16'hC26B,4);
TASK_PP(16'hC26C,4);
TASK_PP(16'hC26D,4);
TASK_PP(16'hC26E,4);
TASK_PP(16'hC26F,4);
TASK_PP(16'hC270,4);
TASK_PP(16'hC271,4);
TASK_PP(16'hC272,4);
TASK_PP(16'hC273,4);
TASK_PP(16'hC274,4);
TASK_PP(16'hC275,4);
TASK_PP(16'hC276,4);
TASK_PP(16'hC277,4);
TASK_PP(16'hC278,4);
TASK_PP(16'hC279,4);
TASK_PP(16'hC27A,4);
TASK_PP(16'hC27B,4);
TASK_PP(16'hC27C,4);
TASK_PP(16'hC27D,4);
TASK_PP(16'hC27E,4);
TASK_PP(16'hC27F,4);
TASK_PP(16'hC280,4);
TASK_PP(16'hC281,4);
TASK_PP(16'hC282,4);
TASK_PP(16'hC283,4);
TASK_PP(16'hC284,4);
TASK_PP(16'hC285,4);
TASK_PP(16'hC286,4);
TASK_PP(16'hC287,4);
TASK_PP(16'hC288,4);
TASK_PP(16'hC289,4);
TASK_PP(16'hC28A,4);
TASK_PP(16'hC28B,4);
TASK_PP(16'hC28C,4);
TASK_PP(16'hC28D,4);
TASK_PP(16'hC28E,4);
TASK_PP(16'hC28F,4);
TASK_PP(16'hC290,4);
TASK_PP(16'hC291,4);
TASK_PP(16'hC292,4);
TASK_PP(16'hC293,4);
TASK_PP(16'hC294,4);
TASK_PP(16'hC295,4);
TASK_PP(16'hC296,4);
TASK_PP(16'hC297,4);
TASK_PP(16'hC298,4);
TASK_PP(16'hC299,4);
TASK_PP(16'hC29A,4);
TASK_PP(16'hC29B,4);
TASK_PP(16'hC29C,4);
TASK_PP(16'hC29D,4);
TASK_PP(16'hC29E,4);
TASK_PP(16'hC29F,4);
TASK_PP(16'hC2A0,4);
TASK_PP(16'hC2A1,4);
TASK_PP(16'hC2A2,4);
TASK_PP(16'hC2A3,4);
TASK_PP(16'hC2A4,4);
TASK_PP(16'hC2A5,4);
TASK_PP(16'hC2A6,4);
TASK_PP(16'hC2A7,4);
TASK_PP(16'hC2A8,4);
TASK_PP(16'hC2A9,4);
TASK_PP(16'hC2AA,4);
TASK_PP(16'hC2AB,4);
TASK_PP(16'hC2AC,4);
TASK_PP(16'hC2AD,4);
TASK_PP(16'hC2AE,4);
TASK_PP(16'hC2AF,4);
TASK_PP(16'hC2B0,4);
TASK_PP(16'hC2B1,4);
TASK_PP(16'hC2B2,4);
TASK_PP(16'hC2B3,4);
TASK_PP(16'hC2B4,4);
TASK_PP(16'hC2B5,4);
TASK_PP(16'hC2B6,4);
TASK_PP(16'hC2B7,4);
TASK_PP(16'hC2B8,4);
TASK_PP(16'hC2B9,4);
TASK_PP(16'hC2BA,4);
TASK_PP(16'hC2BB,4);
TASK_PP(16'hC2BC,4);
TASK_PP(16'hC2BD,4);
TASK_PP(16'hC2BE,4);
TASK_PP(16'hC2BF,4);
TASK_PP(16'hC2C0,4);
TASK_PP(16'hC2C1,4);
TASK_PP(16'hC2C2,4);
TASK_PP(16'hC2C3,4);
TASK_PP(16'hC2C4,4);
TASK_PP(16'hC2C5,4);
TASK_PP(16'hC2C6,4);
TASK_PP(16'hC2C7,4);
TASK_PP(16'hC2C8,4);
TASK_PP(16'hC2C9,4);
TASK_PP(16'hC2CA,4);
TASK_PP(16'hC2CB,4);
TASK_PP(16'hC2CC,4);
TASK_PP(16'hC2CD,4);
TASK_PP(16'hC2CE,4);
TASK_PP(16'hC2CF,4);
TASK_PP(16'hC2D0,4);
TASK_PP(16'hC2D1,4);
TASK_PP(16'hC2D2,4);
TASK_PP(16'hC2D3,4);
TASK_PP(16'hC2D4,4);
TASK_PP(16'hC2D5,4);
TASK_PP(16'hC2D6,4);
TASK_PP(16'hC2D7,4);
TASK_PP(16'hC2D8,4);
TASK_PP(16'hC2D9,4);
TASK_PP(16'hC2DA,4);
TASK_PP(16'hC2DB,4);
TASK_PP(16'hC2DC,4);
TASK_PP(16'hC2DD,4);
TASK_PP(16'hC2DE,4);
TASK_PP(16'hC2DF,4);
TASK_PP(16'hC2E0,4);
TASK_PP(16'hC2E1,4);
TASK_PP(16'hC2E2,4);
TASK_PP(16'hC2E3,4);
TASK_PP(16'hC2E4,4);
TASK_PP(16'hC2E5,4);
TASK_PP(16'hC2E6,4);
TASK_PP(16'hC2E7,4);
TASK_PP(16'hC2E8,4);
TASK_PP(16'hC2E9,4);
TASK_PP(16'hC2EA,4);
TASK_PP(16'hC2EB,4);
TASK_PP(16'hC2EC,4);
TASK_PP(16'hC2ED,4);
TASK_PP(16'hC2EE,4);
TASK_PP(16'hC2EF,4);
TASK_PP(16'hC2F0,4);
TASK_PP(16'hC2F1,4);
TASK_PP(16'hC2F2,4);
TASK_PP(16'hC2F3,4);
TASK_PP(16'hC2F4,4);
TASK_PP(16'hC2F5,4);
TASK_PP(16'hC2F6,4);
TASK_PP(16'hC2F7,4);
TASK_PP(16'hC2F8,4);
TASK_PP(16'hC2F9,4);
TASK_PP(16'hC2FA,4);
TASK_PP(16'hC2FB,4);
TASK_PP(16'hC2FC,4);
TASK_PP(16'hC2FD,4);
TASK_PP(16'hC2FE,4);
TASK_PP(16'hC2FF,4);
TASK_PP(16'hC300,4);
TASK_PP(16'hC301,4);
TASK_PP(16'hC302,4);
TASK_PP(16'hC303,4);
TASK_PP(16'hC304,4);
TASK_PP(16'hC305,4);
TASK_PP(16'hC306,4);
TASK_PP(16'hC307,4);
TASK_PP(16'hC308,4);
TASK_PP(16'hC309,4);
TASK_PP(16'hC30A,4);
TASK_PP(16'hC30B,4);
TASK_PP(16'hC30C,4);
TASK_PP(16'hC30D,4);
TASK_PP(16'hC30E,4);
TASK_PP(16'hC30F,4);
TASK_PP(16'hC310,4);
TASK_PP(16'hC311,4);
TASK_PP(16'hC312,4);
TASK_PP(16'hC313,4);
TASK_PP(16'hC314,4);
TASK_PP(16'hC315,4);
TASK_PP(16'hC316,4);
TASK_PP(16'hC317,4);
TASK_PP(16'hC318,4);
TASK_PP(16'hC319,4);
TASK_PP(16'hC31A,4);
TASK_PP(16'hC31B,4);
TASK_PP(16'hC31C,4);
TASK_PP(16'hC31D,4);
TASK_PP(16'hC31E,4);
TASK_PP(16'hC31F,4);
TASK_PP(16'hC320,4);
TASK_PP(16'hC321,4);
TASK_PP(16'hC322,4);
TASK_PP(16'hC323,4);
TASK_PP(16'hC324,4);
TASK_PP(16'hC325,4);
TASK_PP(16'hC326,4);
TASK_PP(16'hC327,4);
TASK_PP(16'hC328,4);
TASK_PP(16'hC329,4);
TASK_PP(16'hC32A,4);
TASK_PP(16'hC32B,4);
TASK_PP(16'hC32C,4);
TASK_PP(16'hC32D,4);
TASK_PP(16'hC32E,4);
TASK_PP(16'hC32F,4);
TASK_PP(16'hC330,4);
TASK_PP(16'hC331,4);
TASK_PP(16'hC332,4);
TASK_PP(16'hC333,4);
TASK_PP(16'hC334,4);
TASK_PP(16'hC335,4);
TASK_PP(16'hC336,4);
TASK_PP(16'hC337,4);
TASK_PP(16'hC338,4);
TASK_PP(16'hC339,4);
TASK_PP(16'hC33A,4);
TASK_PP(16'hC33B,4);
TASK_PP(16'hC33C,4);
TASK_PP(16'hC33D,4);
TASK_PP(16'hC33E,4);
TASK_PP(16'hC33F,4);
TASK_PP(16'hC340,4);
TASK_PP(16'hC341,4);
TASK_PP(16'hC342,4);
TASK_PP(16'hC343,4);
TASK_PP(16'hC344,4);
TASK_PP(16'hC345,4);
TASK_PP(16'hC346,4);
TASK_PP(16'hC347,4);
TASK_PP(16'hC348,4);
TASK_PP(16'hC349,4);
TASK_PP(16'hC34A,4);
TASK_PP(16'hC34B,4);
TASK_PP(16'hC34C,4);
TASK_PP(16'hC34D,4);
TASK_PP(16'hC34E,4);
TASK_PP(16'hC34F,4);
TASK_PP(16'hC350,4);
TASK_PP(16'hC351,4);
TASK_PP(16'hC352,4);
TASK_PP(16'hC353,4);
TASK_PP(16'hC354,4);
TASK_PP(16'hC355,4);
TASK_PP(16'hC356,4);
TASK_PP(16'hC357,4);
TASK_PP(16'hC358,4);
TASK_PP(16'hC359,4);
TASK_PP(16'hC35A,4);
TASK_PP(16'hC35B,4);
TASK_PP(16'hC35C,4);
TASK_PP(16'hC35D,4);
TASK_PP(16'hC35E,4);
TASK_PP(16'hC35F,4);
TASK_PP(16'hC360,4);
TASK_PP(16'hC361,4);
TASK_PP(16'hC362,4);
TASK_PP(16'hC363,4);
TASK_PP(16'hC364,4);
TASK_PP(16'hC365,4);
TASK_PP(16'hC366,4);
TASK_PP(16'hC367,4);
TASK_PP(16'hC368,4);
TASK_PP(16'hC369,4);
TASK_PP(16'hC36A,4);
TASK_PP(16'hC36B,4);
TASK_PP(16'hC36C,4);
TASK_PP(16'hC36D,4);
TASK_PP(16'hC36E,4);
TASK_PP(16'hC36F,4);
TASK_PP(16'hC370,4);
TASK_PP(16'hC371,4);
TASK_PP(16'hC372,4);
TASK_PP(16'hC373,4);
TASK_PP(16'hC374,4);
TASK_PP(16'hC375,4);
TASK_PP(16'hC376,4);
TASK_PP(16'hC377,4);
TASK_PP(16'hC378,4);
TASK_PP(16'hC379,4);
TASK_PP(16'hC37A,4);
TASK_PP(16'hC37B,4);
TASK_PP(16'hC37C,4);
TASK_PP(16'hC37D,4);
TASK_PP(16'hC37E,4);
TASK_PP(16'hC37F,4);
TASK_PP(16'hC380,4);
TASK_PP(16'hC381,4);
TASK_PP(16'hC382,4);
TASK_PP(16'hC383,4);
TASK_PP(16'hC384,4);
TASK_PP(16'hC385,4);
TASK_PP(16'hC386,4);
TASK_PP(16'hC387,4);
TASK_PP(16'hC388,4);
TASK_PP(16'hC389,4);
TASK_PP(16'hC38A,4);
TASK_PP(16'hC38B,4);
TASK_PP(16'hC38C,4);
TASK_PP(16'hC38D,4);
TASK_PP(16'hC38E,4);
TASK_PP(16'hC38F,4);
TASK_PP(16'hC390,4);
TASK_PP(16'hC391,4);
TASK_PP(16'hC392,4);
TASK_PP(16'hC393,4);
TASK_PP(16'hC394,4);
TASK_PP(16'hC395,4);
TASK_PP(16'hC396,4);
TASK_PP(16'hC397,4);
TASK_PP(16'hC398,4);
TASK_PP(16'hC399,4);
TASK_PP(16'hC39A,4);
TASK_PP(16'hC39B,4);
TASK_PP(16'hC39C,4);
TASK_PP(16'hC39D,4);
TASK_PP(16'hC39E,4);
TASK_PP(16'hC39F,4);
TASK_PP(16'hC3A0,4);
TASK_PP(16'hC3A1,4);
TASK_PP(16'hC3A2,4);
TASK_PP(16'hC3A3,4);
TASK_PP(16'hC3A4,4);
TASK_PP(16'hC3A5,4);
TASK_PP(16'hC3A6,4);
TASK_PP(16'hC3A7,4);
TASK_PP(16'hC3A8,4);
TASK_PP(16'hC3A9,4);
TASK_PP(16'hC3AA,4);
TASK_PP(16'hC3AB,4);
TASK_PP(16'hC3AC,4);
TASK_PP(16'hC3AD,4);
TASK_PP(16'hC3AE,4);
TASK_PP(16'hC3AF,4);
TASK_PP(16'hC3B0,4);
TASK_PP(16'hC3B1,4);
TASK_PP(16'hC3B2,4);
TASK_PP(16'hC3B3,4);
TASK_PP(16'hC3B4,4);
TASK_PP(16'hC3B5,4);
TASK_PP(16'hC3B6,4);
TASK_PP(16'hC3B7,4);
TASK_PP(16'hC3B8,4);
TASK_PP(16'hC3B9,4);
TASK_PP(16'hC3BA,4);
TASK_PP(16'hC3BB,4);
TASK_PP(16'hC3BC,4);
TASK_PP(16'hC3BD,4);
TASK_PP(16'hC3BE,4);
TASK_PP(16'hC3BF,4);
TASK_PP(16'hC3C0,4);
TASK_PP(16'hC3C1,4);
TASK_PP(16'hC3C2,4);
TASK_PP(16'hC3C3,4);
TASK_PP(16'hC3C4,4);
TASK_PP(16'hC3C5,4);
TASK_PP(16'hC3C6,4);
TASK_PP(16'hC3C7,4);
TASK_PP(16'hC3C8,4);
TASK_PP(16'hC3C9,4);
TASK_PP(16'hC3CA,4);
TASK_PP(16'hC3CB,4);
TASK_PP(16'hC3CC,4);
TASK_PP(16'hC3CD,4);
TASK_PP(16'hC3CE,4);
TASK_PP(16'hC3CF,4);
TASK_PP(16'hC3D0,4);
TASK_PP(16'hC3D1,4);
TASK_PP(16'hC3D2,4);
TASK_PP(16'hC3D3,4);
TASK_PP(16'hC3D4,4);
TASK_PP(16'hC3D5,4);
TASK_PP(16'hC3D6,4);
TASK_PP(16'hC3D7,4);
TASK_PP(16'hC3D8,4);
TASK_PP(16'hC3D9,4);
TASK_PP(16'hC3DA,4);
TASK_PP(16'hC3DB,4);
TASK_PP(16'hC3DC,4);
TASK_PP(16'hC3DD,4);
TASK_PP(16'hC3DE,4);
TASK_PP(16'hC3DF,4);
TASK_PP(16'hC3E0,4);
TASK_PP(16'hC3E1,4);
TASK_PP(16'hC3E2,4);
TASK_PP(16'hC3E3,4);
TASK_PP(16'hC3E4,4);
TASK_PP(16'hC3E5,4);
TASK_PP(16'hC3E6,4);
TASK_PP(16'hC3E7,4);
TASK_PP(16'hC3E8,4);
TASK_PP(16'hC3E9,4);
TASK_PP(16'hC3EA,4);
TASK_PP(16'hC3EB,4);
TASK_PP(16'hC3EC,4);
TASK_PP(16'hC3ED,4);
TASK_PP(16'hC3EE,4);
TASK_PP(16'hC3EF,4);
TASK_PP(16'hC3F0,4);
TASK_PP(16'hC3F1,4);
TASK_PP(16'hC3F2,4);
TASK_PP(16'hC3F3,4);
TASK_PP(16'hC3F4,4);
TASK_PP(16'hC3F5,4);
TASK_PP(16'hC3F6,4);
TASK_PP(16'hC3F7,4);
TASK_PP(16'hC3F8,4);
TASK_PP(16'hC3F9,4);
TASK_PP(16'hC3FA,4);
TASK_PP(16'hC3FB,4);
TASK_PP(16'hC3FC,4);
TASK_PP(16'hC3FD,4);
TASK_PP(16'hC3FE,4);
TASK_PP(16'hC3FF,4);
TASK_PP(16'hC400,4);
TASK_PP(16'hC401,4);
TASK_PP(16'hC402,4);
TASK_PP(16'hC403,4);
TASK_PP(16'hC404,4);
TASK_PP(16'hC405,4);
TASK_PP(16'hC406,4);
TASK_PP(16'hC407,4);
TASK_PP(16'hC408,4);
TASK_PP(16'hC409,4);
TASK_PP(16'hC40A,4);
TASK_PP(16'hC40B,4);
TASK_PP(16'hC40C,4);
TASK_PP(16'hC40D,4);
TASK_PP(16'hC40E,4);
TASK_PP(16'hC40F,4);
TASK_PP(16'hC410,4);
TASK_PP(16'hC411,4);
TASK_PP(16'hC412,4);
TASK_PP(16'hC413,4);
TASK_PP(16'hC414,4);
TASK_PP(16'hC415,4);
TASK_PP(16'hC416,4);
TASK_PP(16'hC417,4);
TASK_PP(16'hC418,4);
TASK_PP(16'hC419,4);
TASK_PP(16'hC41A,4);
TASK_PP(16'hC41B,4);
TASK_PP(16'hC41C,4);
TASK_PP(16'hC41D,4);
TASK_PP(16'hC41E,4);
TASK_PP(16'hC41F,4);
TASK_PP(16'hC420,4);
TASK_PP(16'hC421,4);
TASK_PP(16'hC422,4);
TASK_PP(16'hC423,4);
TASK_PP(16'hC424,4);
TASK_PP(16'hC425,4);
TASK_PP(16'hC426,4);
TASK_PP(16'hC427,4);
TASK_PP(16'hC428,4);
TASK_PP(16'hC429,4);
TASK_PP(16'hC42A,4);
TASK_PP(16'hC42B,4);
TASK_PP(16'hC42C,4);
TASK_PP(16'hC42D,4);
TASK_PP(16'hC42E,4);
TASK_PP(16'hC42F,4);
TASK_PP(16'hC430,4);
TASK_PP(16'hC431,4);
TASK_PP(16'hC432,4);
TASK_PP(16'hC433,4);
TASK_PP(16'hC434,4);
TASK_PP(16'hC435,4);
TASK_PP(16'hC436,4);
TASK_PP(16'hC437,4);
TASK_PP(16'hC438,4);
TASK_PP(16'hC439,4);
TASK_PP(16'hC43A,4);
TASK_PP(16'hC43B,4);
TASK_PP(16'hC43C,4);
TASK_PP(16'hC43D,4);
TASK_PP(16'hC43E,4);
TASK_PP(16'hC43F,4);
TASK_PP(16'hC440,4);
TASK_PP(16'hC441,4);
TASK_PP(16'hC442,4);
TASK_PP(16'hC443,4);
TASK_PP(16'hC444,4);
TASK_PP(16'hC445,4);
TASK_PP(16'hC446,4);
TASK_PP(16'hC447,4);
TASK_PP(16'hC448,4);
TASK_PP(16'hC449,4);
TASK_PP(16'hC44A,4);
TASK_PP(16'hC44B,4);
TASK_PP(16'hC44C,4);
TASK_PP(16'hC44D,4);
TASK_PP(16'hC44E,4);
TASK_PP(16'hC44F,4);
TASK_PP(16'hC450,4);
TASK_PP(16'hC451,4);
TASK_PP(16'hC452,4);
TASK_PP(16'hC453,4);
TASK_PP(16'hC454,4);
TASK_PP(16'hC455,4);
TASK_PP(16'hC456,4);
TASK_PP(16'hC457,4);
TASK_PP(16'hC458,4);
TASK_PP(16'hC459,4);
TASK_PP(16'hC45A,4);
TASK_PP(16'hC45B,4);
TASK_PP(16'hC45C,4);
TASK_PP(16'hC45D,4);
TASK_PP(16'hC45E,4);
TASK_PP(16'hC45F,4);
TASK_PP(16'hC460,4);
TASK_PP(16'hC461,4);
TASK_PP(16'hC462,4);
TASK_PP(16'hC463,4);
TASK_PP(16'hC464,4);
TASK_PP(16'hC465,4);
TASK_PP(16'hC466,4);
TASK_PP(16'hC467,4);
TASK_PP(16'hC468,4);
TASK_PP(16'hC469,4);
TASK_PP(16'hC46A,4);
TASK_PP(16'hC46B,4);
TASK_PP(16'hC46C,4);
TASK_PP(16'hC46D,4);
TASK_PP(16'hC46E,4);
TASK_PP(16'hC46F,4);
TASK_PP(16'hC470,4);
TASK_PP(16'hC471,4);
TASK_PP(16'hC472,4);
TASK_PP(16'hC473,4);
TASK_PP(16'hC474,4);
TASK_PP(16'hC475,4);
TASK_PP(16'hC476,4);
TASK_PP(16'hC477,4);
TASK_PP(16'hC478,4);
TASK_PP(16'hC479,4);
TASK_PP(16'hC47A,4);
TASK_PP(16'hC47B,4);
TASK_PP(16'hC47C,4);
TASK_PP(16'hC47D,4);
TASK_PP(16'hC47E,4);
TASK_PP(16'hC47F,4);
TASK_PP(16'hC480,4);
TASK_PP(16'hC481,4);
TASK_PP(16'hC482,4);
TASK_PP(16'hC483,4);
TASK_PP(16'hC484,4);
TASK_PP(16'hC485,4);
TASK_PP(16'hC486,4);
TASK_PP(16'hC487,4);
TASK_PP(16'hC488,4);
TASK_PP(16'hC489,4);
TASK_PP(16'hC48A,4);
TASK_PP(16'hC48B,4);
TASK_PP(16'hC48C,4);
TASK_PP(16'hC48D,4);
TASK_PP(16'hC48E,4);
TASK_PP(16'hC48F,4);
TASK_PP(16'hC490,4);
TASK_PP(16'hC491,4);
TASK_PP(16'hC492,4);
TASK_PP(16'hC493,4);
TASK_PP(16'hC494,4);
TASK_PP(16'hC495,4);
TASK_PP(16'hC496,4);
TASK_PP(16'hC497,4);
TASK_PP(16'hC498,4);
TASK_PP(16'hC499,4);
TASK_PP(16'hC49A,4);
TASK_PP(16'hC49B,4);
TASK_PP(16'hC49C,4);
TASK_PP(16'hC49D,4);
TASK_PP(16'hC49E,4);
TASK_PP(16'hC49F,4);
TASK_PP(16'hC4A0,4);
TASK_PP(16'hC4A1,4);
TASK_PP(16'hC4A2,4);
TASK_PP(16'hC4A3,4);
TASK_PP(16'hC4A4,4);
TASK_PP(16'hC4A5,4);
TASK_PP(16'hC4A6,4);
TASK_PP(16'hC4A7,4);
TASK_PP(16'hC4A8,4);
TASK_PP(16'hC4A9,4);
TASK_PP(16'hC4AA,4);
TASK_PP(16'hC4AB,4);
TASK_PP(16'hC4AC,4);
TASK_PP(16'hC4AD,4);
TASK_PP(16'hC4AE,4);
TASK_PP(16'hC4AF,4);
TASK_PP(16'hC4B0,4);
TASK_PP(16'hC4B1,4);
TASK_PP(16'hC4B2,4);
TASK_PP(16'hC4B3,4);
TASK_PP(16'hC4B4,4);
TASK_PP(16'hC4B5,4);
TASK_PP(16'hC4B6,4);
TASK_PP(16'hC4B7,4);
TASK_PP(16'hC4B8,4);
TASK_PP(16'hC4B9,4);
TASK_PP(16'hC4BA,4);
TASK_PP(16'hC4BB,4);
TASK_PP(16'hC4BC,4);
TASK_PP(16'hC4BD,4);
TASK_PP(16'hC4BE,4);
TASK_PP(16'hC4BF,4);
TASK_PP(16'hC4C0,4);
TASK_PP(16'hC4C1,4);
TASK_PP(16'hC4C2,4);
TASK_PP(16'hC4C3,4);
TASK_PP(16'hC4C4,4);
TASK_PP(16'hC4C5,4);
TASK_PP(16'hC4C6,4);
TASK_PP(16'hC4C7,4);
TASK_PP(16'hC4C8,4);
TASK_PP(16'hC4C9,4);
TASK_PP(16'hC4CA,4);
TASK_PP(16'hC4CB,4);
TASK_PP(16'hC4CC,4);
TASK_PP(16'hC4CD,4);
TASK_PP(16'hC4CE,4);
TASK_PP(16'hC4CF,4);
TASK_PP(16'hC4D0,4);
TASK_PP(16'hC4D1,4);
TASK_PP(16'hC4D2,4);
TASK_PP(16'hC4D3,4);
TASK_PP(16'hC4D4,4);
TASK_PP(16'hC4D5,4);
TASK_PP(16'hC4D6,4);
TASK_PP(16'hC4D7,4);
TASK_PP(16'hC4D8,4);
TASK_PP(16'hC4D9,4);
TASK_PP(16'hC4DA,4);
TASK_PP(16'hC4DB,4);
TASK_PP(16'hC4DC,4);
TASK_PP(16'hC4DD,4);
TASK_PP(16'hC4DE,4);
TASK_PP(16'hC4DF,4);
TASK_PP(16'hC4E0,4);
TASK_PP(16'hC4E1,4);
TASK_PP(16'hC4E2,4);
TASK_PP(16'hC4E3,4);
TASK_PP(16'hC4E4,4);
TASK_PP(16'hC4E5,4);
TASK_PP(16'hC4E6,4);
TASK_PP(16'hC4E7,4);
TASK_PP(16'hC4E8,4);
TASK_PP(16'hC4E9,4);
TASK_PP(16'hC4EA,4);
TASK_PP(16'hC4EB,4);
TASK_PP(16'hC4EC,4);
TASK_PP(16'hC4ED,4);
TASK_PP(16'hC4EE,4);
TASK_PP(16'hC4EF,4);
TASK_PP(16'hC4F0,4);
TASK_PP(16'hC4F1,4);
TASK_PP(16'hC4F2,4);
TASK_PP(16'hC4F3,4);
TASK_PP(16'hC4F4,4);
TASK_PP(16'hC4F5,4);
TASK_PP(16'hC4F6,4);
TASK_PP(16'hC4F7,4);
TASK_PP(16'hC4F8,4);
TASK_PP(16'hC4F9,4);
TASK_PP(16'hC4FA,4);
TASK_PP(16'hC4FB,4);
TASK_PP(16'hC4FC,4);
TASK_PP(16'hC4FD,4);
TASK_PP(16'hC4FE,4);
TASK_PP(16'hC4FF,4);
TASK_PP(16'hC500,4);
TASK_PP(16'hC501,4);
TASK_PP(16'hC502,4);
TASK_PP(16'hC503,4);
TASK_PP(16'hC504,4);
TASK_PP(16'hC505,4);
TASK_PP(16'hC506,4);
TASK_PP(16'hC507,4);
TASK_PP(16'hC508,4);
TASK_PP(16'hC509,4);
TASK_PP(16'hC50A,4);
TASK_PP(16'hC50B,4);
TASK_PP(16'hC50C,4);
TASK_PP(16'hC50D,4);
TASK_PP(16'hC50E,4);
TASK_PP(16'hC50F,4);
TASK_PP(16'hC510,4);
TASK_PP(16'hC511,4);
TASK_PP(16'hC512,4);
TASK_PP(16'hC513,4);
TASK_PP(16'hC514,4);
TASK_PP(16'hC515,4);
TASK_PP(16'hC516,4);
TASK_PP(16'hC517,4);
TASK_PP(16'hC518,4);
TASK_PP(16'hC519,4);
TASK_PP(16'hC51A,4);
TASK_PP(16'hC51B,4);
TASK_PP(16'hC51C,4);
TASK_PP(16'hC51D,4);
TASK_PP(16'hC51E,4);
TASK_PP(16'hC51F,4);
TASK_PP(16'hC520,4);
TASK_PP(16'hC521,4);
TASK_PP(16'hC522,4);
TASK_PP(16'hC523,4);
TASK_PP(16'hC524,4);
TASK_PP(16'hC525,4);
TASK_PP(16'hC526,4);
TASK_PP(16'hC527,4);
TASK_PP(16'hC528,4);
TASK_PP(16'hC529,4);
TASK_PP(16'hC52A,4);
TASK_PP(16'hC52B,4);
TASK_PP(16'hC52C,4);
TASK_PP(16'hC52D,4);
TASK_PP(16'hC52E,4);
TASK_PP(16'hC52F,4);
TASK_PP(16'hC530,4);
TASK_PP(16'hC531,4);
TASK_PP(16'hC532,4);
TASK_PP(16'hC533,4);
TASK_PP(16'hC534,4);
TASK_PP(16'hC535,4);
TASK_PP(16'hC536,4);
TASK_PP(16'hC537,4);
TASK_PP(16'hC538,4);
TASK_PP(16'hC539,4);
TASK_PP(16'hC53A,4);
TASK_PP(16'hC53B,4);
TASK_PP(16'hC53C,4);
TASK_PP(16'hC53D,4);
TASK_PP(16'hC53E,4);
TASK_PP(16'hC53F,4);
TASK_PP(16'hC540,4);
TASK_PP(16'hC541,4);
TASK_PP(16'hC542,4);
TASK_PP(16'hC543,4);
TASK_PP(16'hC544,4);
TASK_PP(16'hC545,4);
TASK_PP(16'hC546,4);
TASK_PP(16'hC547,4);
TASK_PP(16'hC548,4);
TASK_PP(16'hC549,4);
TASK_PP(16'hC54A,4);
TASK_PP(16'hC54B,4);
TASK_PP(16'hC54C,4);
TASK_PP(16'hC54D,4);
TASK_PP(16'hC54E,4);
TASK_PP(16'hC54F,4);
TASK_PP(16'hC550,4);
TASK_PP(16'hC551,4);
TASK_PP(16'hC552,4);
TASK_PP(16'hC553,4);
TASK_PP(16'hC554,4);
TASK_PP(16'hC555,4);
TASK_PP(16'hC556,4);
TASK_PP(16'hC557,4);
TASK_PP(16'hC558,4);
TASK_PP(16'hC559,4);
TASK_PP(16'hC55A,4);
TASK_PP(16'hC55B,4);
TASK_PP(16'hC55C,4);
TASK_PP(16'hC55D,4);
TASK_PP(16'hC55E,4);
TASK_PP(16'hC55F,4);
TASK_PP(16'hC560,4);
TASK_PP(16'hC561,4);
TASK_PP(16'hC562,4);
TASK_PP(16'hC563,4);
TASK_PP(16'hC564,4);
TASK_PP(16'hC565,4);
TASK_PP(16'hC566,4);
TASK_PP(16'hC567,4);
TASK_PP(16'hC568,4);
TASK_PP(16'hC569,4);
TASK_PP(16'hC56A,4);
TASK_PP(16'hC56B,4);
TASK_PP(16'hC56C,4);
TASK_PP(16'hC56D,4);
TASK_PP(16'hC56E,4);
TASK_PP(16'hC56F,4);
TASK_PP(16'hC570,4);
TASK_PP(16'hC571,4);
TASK_PP(16'hC572,4);
TASK_PP(16'hC573,4);
TASK_PP(16'hC574,4);
TASK_PP(16'hC575,4);
TASK_PP(16'hC576,4);
TASK_PP(16'hC577,4);
TASK_PP(16'hC578,4);
TASK_PP(16'hC579,4);
TASK_PP(16'hC57A,4);
TASK_PP(16'hC57B,4);
TASK_PP(16'hC57C,4);
TASK_PP(16'hC57D,4);
TASK_PP(16'hC57E,4);
TASK_PP(16'hC57F,4);
TASK_PP(16'hC580,4);
TASK_PP(16'hC581,4);
TASK_PP(16'hC582,4);
TASK_PP(16'hC583,4);
TASK_PP(16'hC584,4);
TASK_PP(16'hC585,4);
TASK_PP(16'hC586,4);
TASK_PP(16'hC587,4);
TASK_PP(16'hC588,4);
TASK_PP(16'hC589,4);
TASK_PP(16'hC58A,4);
TASK_PP(16'hC58B,4);
TASK_PP(16'hC58C,4);
TASK_PP(16'hC58D,4);
TASK_PP(16'hC58E,4);
TASK_PP(16'hC58F,4);
TASK_PP(16'hC590,4);
TASK_PP(16'hC591,4);
TASK_PP(16'hC592,4);
TASK_PP(16'hC593,4);
TASK_PP(16'hC594,4);
TASK_PP(16'hC595,4);
TASK_PP(16'hC596,4);
TASK_PP(16'hC597,4);
TASK_PP(16'hC598,4);
TASK_PP(16'hC599,4);
TASK_PP(16'hC59A,4);
TASK_PP(16'hC59B,4);
TASK_PP(16'hC59C,4);
TASK_PP(16'hC59D,4);
TASK_PP(16'hC59E,4);
TASK_PP(16'hC59F,4);
TASK_PP(16'hC5A0,4);
TASK_PP(16'hC5A1,4);
TASK_PP(16'hC5A2,4);
TASK_PP(16'hC5A3,4);
TASK_PP(16'hC5A4,4);
TASK_PP(16'hC5A5,4);
TASK_PP(16'hC5A6,4);
TASK_PP(16'hC5A7,4);
TASK_PP(16'hC5A8,4);
TASK_PP(16'hC5A9,4);
TASK_PP(16'hC5AA,4);
TASK_PP(16'hC5AB,4);
TASK_PP(16'hC5AC,4);
TASK_PP(16'hC5AD,4);
TASK_PP(16'hC5AE,4);
TASK_PP(16'hC5AF,4);
TASK_PP(16'hC5B0,4);
TASK_PP(16'hC5B1,4);
TASK_PP(16'hC5B2,4);
TASK_PP(16'hC5B3,4);
TASK_PP(16'hC5B4,4);
TASK_PP(16'hC5B5,4);
TASK_PP(16'hC5B6,4);
TASK_PP(16'hC5B7,4);
TASK_PP(16'hC5B8,4);
TASK_PP(16'hC5B9,4);
TASK_PP(16'hC5BA,4);
TASK_PP(16'hC5BB,4);
TASK_PP(16'hC5BC,4);
TASK_PP(16'hC5BD,4);
TASK_PP(16'hC5BE,4);
TASK_PP(16'hC5BF,4);
TASK_PP(16'hC5C0,4);
TASK_PP(16'hC5C1,4);
TASK_PP(16'hC5C2,4);
TASK_PP(16'hC5C3,4);
TASK_PP(16'hC5C4,4);
TASK_PP(16'hC5C5,4);
TASK_PP(16'hC5C6,4);
TASK_PP(16'hC5C7,4);
TASK_PP(16'hC5C8,4);
TASK_PP(16'hC5C9,4);
TASK_PP(16'hC5CA,4);
TASK_PP(16'hC5CB,4);
TASK_PP(16'hC5CC,4);
TASK_PP(16'hC5CD,4);
TASK_PP(16'hC5CE,4);
TASK_PP(16'hC5CF,4);
TASK_PP(16'hC5D0,4);
TASK_PP(16'hC5D1,4);
TASK_PP(16'hC5D2,4);
TASK_PP(16'hC5D3,4);
TASK_PP(16'hC5D4,4);
TASK_PP(16'hC5D5,4);
TASK_PP(16'hC5D6,4);
TASK_PP(16'hC5D7,4);
TASK_PP(16'hC5D8,4);
TASK_PP(16'hC5D9,4);
TASK_PP(16'hC5DA,4);
TASK_PP(16'hC5DB,4);
TASK_PP(16'hC5DC,4);
TASK_PP(16'hC5DD,4);
TASK_PP(16'hC5DE,4);
TASK_PP(16'hC5DF,4);
TASK_PP(16'hC5E0,4);
TASK_PP(16'hC5E1,4);
TASK_PP(16'hC5E2,4);
TASK_PP(16'hC5E3,4);
TASK_PP(16'hC5E4,4);
TASK_PP(16'hC5E5,4);
TASK_PP(16'hC5E6,4);
TASK_PP(16'hC5E7,4);
TASK_PP(16'hC5E8,4);
TASK_PP(16'hC5E9,4);
TASK_PP(16'hC5EA,4);
TASK_PP(16'hC5EB,4);
TASK_PP(16'hC5EC,4);
TASK_PP(16'hC5ED,4);
TASK_PP(16'hC5EE,4);
TASK_PP(16'hC5EF,4);
TASK_PP(16'hC5F0,4);
TASK_PP(16'hC5F1,4);
TASK_PP(16'hC5F2,4);
TASK_PP(16'hC5F3,4);
TASK_PP(16'hC5F4,4);
TASK_PP(16'hC5F5,4);
TASK_PP(16'hC5F6,4);
TASK_PP(16'hC5F7,4);
TASK_PP(16'hC5F8,4);
TASK_PP(16'hC5F9,4);
TASK_PP(16'hC5FA,4);
TASK_PP(16'hC5FB,4);
TASK_PP(16'hC5FC,4);
TASK_PP(16'hC5FD,4);
TASK_PP(16'hC5FE,4);
TASK_PP(16'hC5FF,4);
TASK_PP(16'hC600,4);
TASK_PP(16'hC601,4);
TASK_PP(16'hC602,4);
TASK_PP(16'hC603,4);
TASK_PP(16'hC604,4);
TASK_PP(16'hC605,4);
TASK_PP(16'hC606,4);
TASK_PP(16'hC607,4);
TASK_PP(16'hC608,4);
TASK_PP(16'hC609,4);
TASK_PP(16'hC60A,4);
TASK_PP(16'hC60B,4);
TASK_PP(16'hC60C,4);
TASK_PP(16'hC60D,4);
TASK_PP(16'hC60E,4);
TASK_PP(16'hC60F,4);
TASK_PP(16'hC610,4);
TASK_PP(16'hC611,4);
TASK_PP(16'hC612,4);
TASK_PP(16'hC613,4);
TASK_PP(16'hC614,4);
TASK_PP(16'hC615,4);
TASK_PP(16'hC616,4);
TASK_PP(16'hC617,4);
TASK_PP(16'hC618,4);
TASK_PP(16'hC619,4);
TASK_PP(16'hC61A,4);
TASK_PP(16'hC61B,4);
TASK_PP(16'hC61C,4);
TASK_PP(16'hC61D,4);
TASK_PP(16'hC61E,4);
TASK_PP(16'hC61F,4);
TASK_PP(16'hC620,4);
TASK_PP(16'hC621,4);
TASK_PP(16'hC622,4);
TASK_PP(16'hC623,4);
TASK_PP(16'hC624,4);
TASK_PP(16'hC625,4);
TASK_PP(16'hC626,4);
TASK_PP(16'hC627,4);
TASK_PP(16'hC628,4);
TASK_PP(16'hC629,4);
TASK_PP(16'hC62A,4);
TASK_PP(16'hC62B,4);
TASK_PP(16'hC62C,4);
TASK_PP(16'hC62D,4);
TASK_PP(16'hC62E,4);
TASK_PP(16'hC62F,4);
TASK_PP(16'hC630,4);
TASK_PP(16'hC631,4);
TASK_PP(16'hC632,4);
TASK_PP(16'hC633,4);
TASK_PP(16'hC634,4);
TASK_PP(16'hC635,4);
TASK_PP(16'hC636,4);
TASK_PP(16'hC637,4);
TASK_PP(16'hC638,4);
TASK_PP(16'hC639,4);
TASK_PP(16'hC63A,4);
TASK_PP(16'hC63B,4);
TASK_PP(16'hC63C,4);
TASK_PP(16'hC63D,4);
TASK_PP(16'hC63E,4);
TASK_PP(16'hC63F,4);
TASK_PP(16'hC640,4);
TASK_PP(16'hC641,4);
TASK_PP(16'hC642,4);
TASK_PP(16'hC643,4);
TASK_PP(16'hC644,4);
TASK_PP(16'hC645,4);
TASK_PP(16'hC646,4);
TASK_PP(16'hC647,4);
TASK_PP(16'hC648,4);
TASK_PP(16'hC649,4);
TASK_PP(16'hC64A,4);
TASK_PP(16'hC64B,4);
TASK_PP(16'hC64C,4);
TASK_PP(16'hC64D,4);
TASK_PP(16'hC64E,4);
TASK_PP(16'hC64F,4);
TASK_PP(16'hC650,4);
TASK_PP(16'hC651,4);
TASK_PP(16'hC652,4);
TASK_PP(16'hC653,4);
TASK_PP(16'hC654,4);
TASK_PP(16'hC655,4);
TASK_PP(16'hC656,4);
TASK_PP(16'hC657,4);
TASK_PP(16'hC658,4);
TASK_PP(16'hC659,4);
TASK_PP(16'hC65A,4);
TASK_PP(16'hC65B,4);
TASK_PP(16'hC65C,4);
TASK_PP(16'hC65D,4);
TASK_PP(16'hC65E,4);
TASK_PP(16'hC65F,4);
TASK_PP(16'hC660,4);
TASK_PP(16'hC661,4);
TASK_PP(16'hC662,4);
TASK_PP(16'hC663,4);
TASK_PP(16'hC664,4);
TASK_PP(16'hC665,4);
TASK_PP(16'hC666,4);
TASK_PP(16'hC667,4);
TASK_PP(16'hC668,4);
TASK_PP(16'hC669,4);
TASK_PP(16'hC66A,4);
TASK_PP(16'hC66B,4);
TASK_PP(16'hC66C,4);
TASK_PP(16'hC66D,4);
TASK_PP(16'hC66E,4);
TASK_PP(16'hC66F,4);
TASK_PP(16'hC670,4);
TASK_PP(16'hC671,4);
TASK_PP(16'hC672,4);
TASK_PP(16'hC673,4);
TASK_PP(16'hC674,4);
TASK_PP(16'hC675,4);
TASK_PP(16'hC676,4);
TASK_PP(16'hC677,4);
TASK_PP(16'hC678,4);
TASK_PP(16'hC679,4);
TASK_PP(16'hC67A,4);
TASK_PP(16'hC67B,4);
TASK_PP(16'hC67C,4);
TASK_PP(16'hC67D,4);
TASK_PP(16'hC67E,4);
TASK_PP(16'hC67F,4);
TASK_PP(16'hC680,4);
TASK_PP(16'hC681,4);
TASK_PP(16'hC682,4);
TASK_PP(16'hC683,4);
TASK_PP(16'hC684,4);
TASK_PP(16'hC685,4);
TASK_PP(16'hC686,4);
TASK_PP(16'hC687,4);
TASK_PP(16'hC688,4);
TASK_PP(16'hC689,4);
TASK_PP(16'hC68A,4);
TASK_PP(16'hC68B,4);
TASK_PP(16'hC68C,4);
TASK_PP(16'hC68D,4);
TASK_PP(16'hC68E,4);
TASK_PP(16'hC68F,4);
TASK_PP(16'hC690,4);
TASK_PP(16'hC691,4);
TASK_PP(16'hC692,4);
TASK_PP(16'hC693,4);
TASK_PP(16'hC694,4);
TASK_PP(16'hC695,4);
TASK_PP(16'hC696,4);
TASK_PP(16'hC697,4);
TASK_PP(16'hC698,4);
TASK_PP(16'hC699,4);
TASK_PP(16'hC69A,4);
TASK_PP(16'hC69B,4);
TASK_PP(16'hC69C,4);
TASK_PP(16'hC69D,4);
TASK_PP(16'hC69E,4);
TASK_PP(16'hC69F,4);
TASK_PP(16'hC6A0,4);
TASK_PP(16'hC6A1,4);
TASK_PP(16'hC6A2,4);
TASK_PP(16'hC6A3,4);
TASK_PP(16'hC6A4,4);
TASK_PP(16'hC6A5,4);
TASK_PP(16'hC6A6,4);
TASK_PP(16'hC6A7,4);
TASK_PP(16'hC6A8,4);
TASK_PP(16'hC6A9,4);
TASK_PP(16'hC6AA,4);
TASK_PP(16'hC6AB,4);
TASK_PP(16'hC6AC,4);
TASK_PP(16'hC6AD,4);
TASK_PP(16'hC6AE,4);
TASK_PP(16'hC6AF,4);
TASK_PP(16'hC6B0,4);
TASK_PP(16'hC6B1,4);
TASK_PP(16'hC6B2,4);
TASK_PP(16'hC6B3,4);
TASK_PP(16'hC6B4,4);
TASK_PP(16'hC6B5,4);
TASK_PP(16'hC6B6,4);
TASK_PP(16'hC6B7,4);
TASK_PP(16'hC6B8,4);
TASK_PP(16'hC6B9,4);
TASK_PP(16'hC6BA,4);
TASK_PP(16'hC6BB,4);
TASK_PP(16'hC6BC,4);
TASK_PP(16'hC6BD,4);
TASK_PP(16'hC6BE,4);
TASK_PP(16'hC6BF,4);
TASK_PP(16'hC6C0,4);
TASK_PP(16'hC6C1,4);
TASK_PP(16'hC6C2,4);
TASK_PP(16'hC6C3,4);
TASK_PP(16'hC6C4,4);
TASK_PP(16'hC6C5,4);
TASK_PP(16'hC6C6,4);
TASK_PP(16'hC6C7,4);
TASK_PP(16'hC6C8,4);
TASK_PP(16'hC6C9,4);
TASK_PP(16'hC6CA,4);
TASK_PP(16'hC6CB,4);
TASK_PP(16'hC6CC,4);
TASK_PP(16'hC6CD,4);
TASK_PP(16'hC6CE,4);
TASK_PP(16'hC6CF,4);
TASK_PP(16'hC6D0,4);
TASK_PP(16'hC6D1,4);
TASK_PP(16'hC6D2,4);
TASK_PP(16'hC6D3,4);
TASK_PP(16'hC6D4,4);
TASK_PP(16'hC6D5,4);
TASK_PP(16'hC6D6,4);
TASK_PP(16'hC6D7,4);
TASK_PP(16'hC6D8,4);
TASK_PP(16'hC6D9,4);
TASK_PP(16'hC6DA,4);
TASK_PP(16'hC6DB,4);
TASK_PP(16'hC6DC,4);
TASK_PP(16'hC6DD,4);
TASK_PP(16'hC6DE,4);
TASK_PP(16'hC6DF,4);
TASK_PP(16'hC6E0,4);
TASK_PP(16'hC6E1,4);
TASK_PP(16'hC6E2,4);
TASK_PP(16'hC6E3,4);
TASK_PP(16'hC6E4,4);
TASK_PP(16'hC6E5,4);
TASK_PP(16'hC6E6,4);
TASK_PP(16'hC6E7,4);
TASK_PP(16'hC6E8,4);
TASK_PP(16'hC6E9,4);
TASK_PP(16'hC6EA,4);
TASK_PP(16'hC6EB,4);
TASK_PP(16'hC6EC,4);
TASK_PP(16'hC6ED,4);
TASK_PP(16'hC6EE,4);
TASK_PP(16'hC6EF,4);
TASK_PP(16'hC6F0,4);
TASK_PP(16'hC6F1,4);
TASK_PP(16'hC6F2,4);
TASK_PP(16'hC6F3,4);
TASK_PP(16'hC6F4,4);
TASK_PP(16'hC6F5,4);
TASK_PP(16'hC6F6,4);
TASK_PP(16'hC6F7,4);
TASK_PP(16'hC6F8,4);
TASK_PP(16'hC6F9,4);
TASK_PP(16'hC6FA,4);
TASK_PP(16'hC6FB,4);
TASK_PP(16'hC6FC,4);
TASK_PP(16'hC6FD,4);
TASK_PP(16'hC6FE,4);
TASK_PP(16'hC6FF,4);
TASK_PP(16'hC700,4);
TASK_PP(16'hC701,4);
TASK_PP(16'hC702,4);
TASK_PP(16'hC703,4);
TASK_PP(16'hC704,4);
TASK_PP(16'hC705,4);
TASK_PP(16'hC706,4);
TASK_PP(16'hC707,4);
TASK_PP(16'hC708,4);
TASK_PP(16'hC709,4);
TASK_PP(16'hC70A,4);
TASK_PP(16'hC70B,4);
TASK_PP(16'hC70C,4);
TASK_PP(16'hC70D,4);
TASK_PP(16'hC70E,4);
TASK_PP(16'hC70F,4);
TASK_PP(16'hC710,4);
TASK_PP(16'hC711,4);
TASK_PP(16'hC712,4);
TASK_PP(16'hC713,4);
TASK_PP(16'hC714,4);
TASK_PP(16'hC715,4);
TASK_PP(16'hC716,4);
TASK_PP(16'hC717,4);
TASK_PP(16'hC718,4);
TASK_PP(16'hC719,4);
TASK_PP(16'hC71A,4);
TASK_PP(16'hC71B,4);
TASK_PP(16'hC71C,4);
TASK_PP(16'hC71D,4);
TASK_PP(16'hC71E,4);
TASK_PP(16'hC71F,4);
TASK_PP(16'hC720,4);
TASK_PP(16'hC721,4);
TASK_PP(16'hC722,4);
TASK_PP(16'hC723,4);
TASK_PP(16'hC724,4);
TASK_PP(16'hC725,4);
TASK_PP(16'hC726,4);
TASK_PP(16'hC727,4);
TASK_PP(16'hC728,4);
TASK_PP(16'hC729,4);
TASK_PP(16'hC72A,4);
TASK_PP(16'hC72B,4);
TASK_PP(16'hC72C,4);
TASK_PP(16'hC72D,4);
TASK_PP(16'hC72E,4);
TASK_PP(16'hC72F,4);
TASK_PP(16'hC730,4);
TASK_PP(16'hC731,4);
TASK_PP(16'hC732,4);
TASK_PP(16'hC733,4);
TASK_PP(16'hC734,4);
TASK_PP(16'hC735,4);
TASK_PP(16'hC736,4);
TASK_PP(16'hC737,4);
TASK_PP(16'hC738,4);
TASK_PP(16'hC739,4);
TASK_PP(16'hC73A,4);
TASK_PP(16'hC73B,4);
TASK_PP(16'hC73C,4);
TASK_PP(16'hC73D,4);
TASK_PP(16'hC73E,4);
TASK_PP(16'hC73F,4);
TASK_PP(16'hC740,4);
TASK_PP(16'hC741,4);
TASK_PP(16'hC742,4);
TASK_PP(16'hC743,4);
TASK_PP(16'hC744,4);
TASK_PP(16'hC745,4);
TASK_PP(16'hC746,4);
TASK_PP(16'hC747,4);
TASK_PP(16'hC748,4);
TASK_PP(16'hC749,4);
TASK_PP(16'hC74A,4);
TASK_PP(16'hC74B,4);
TASK_PP(16'hC74C,4);
TASK_PP(16'hC74D,4);
TASK_PP(16'hC74E,4);
TASK_PP(16'hC74F,4);
TASK_PP(16'hC750,4);
TASK_PP(16'hC751,4);
TASK_PP(16'hC752,4);
TASK_PP(16'hC753,4);
TASK_PP(16'hC754,4);
TASK_PP(16'hC755,4);
TASK_PP(16'hC756,4);
TASK_PP(16'hC757,4);
TASK_PP(16'hC758,4);
TASK_PP(16'hC759,4);
TASK_PP(16'hC75A,4);
TASK_PP(16'hC75B,4);
TASK_PP(16'hC75C,4);
TASK_PP(16'hC75D,4);
TASK_PP(16'hC75E,4);
TASK_PP(16'hC75F,4);
TASK_PP(16'hC760,4);
TASK_PP(16'hC761,4);
TASK_PP(16'hC762,4);
TASK_PP(16'hC763,4);
TASK_PP(16'hC764,4);
TASK_PP(16'hC765,4);
TASK_PP(16'hC766,4);
TASK_PP(16'hC767,4);
TASK_PP(16'hC768,4);
TASK_PP(16'hC769,4);
TASK_PP(16'hC76A,4);
TASK_PP(16'hC76B,4);
TASK_PP(16'hC76C,4);
TASK_PP(16'hC76D,4);
TASK_PP(16'hC76E,4);
TASK_PP(16'hC76F,4);
TASK_PP(16'hC770,4);
TASK_PP(16'hC771,4);
TASK_PP(16'hC772,4);
TASK_PP(16'hC773,4);
TASK_PP(16'hC774,4);
TASK_PP(16'hC775,4);
TASK_PP(16'hC776,4);
TASK_PP(16'hC777,4);
TASK_PP(16'hC778,4);
TASK_PP(16'hC779,4);
TASK_PP(16'hC77A,4);
TASK_PP(16'hC77B,4);
TASK_PP(16'hC77C,4);
TASK_PP(16'hC77D,4);
TASK_PP(16'hC77E,4);
TASK_PP(16'hC77F,4);
TASK_PP(16'hC780,4);
TASK_PP(16'hC781,4);
TASK_PP(16'hC782,4);
TASK_PP(16'hC783,4);
TASK_PP(16'hC784,4);
TASK_PP(16'hC785,4);
TASK_PP(16'hC786,4);
TASK_PP(16'hC787,4);
TASK_PP(16'hC788,4);
TASK_PP(16'hC789,4);
TASK_PP(16'hC78A,4);
TASK_PP(16'hC78B,4);
TASK_PP(16'hC78C,4);
TASK_PP(16'hC78D,4);
TASK_PP(16'hC78E,4);
TASK_PP(16'hC78F,4);
TASK_PP(16'hC790,4);
TASK_PP(16'hC791,4);
TASK_PP(16'hC792,4);
TASK_PP(16'hC793,4);
TASK_PP(16'hC794,4);
TASK_PP(16'hC795,4);
TASK_PP(16'hC796,4);
TASK_PP(16'hC797,4);
TASK_PP(16'hC798,4);
TASK_PP(16'hC799,4);
TASK_PP(16'hC79A,4);
TASK_PP(16'hC79B,4);
TASK_PP(16'hC79C,4);
TASK_PP(16'hC79D,4);
TASK_PP(16'hC79E,4);
TASK_PP(16'hC79F,4);
TASK_PP(16'hC7A0,4);
TASK_PP(16'hC7A1,4);
TASK_PP(16'hC7A2,4);
TASK_PP(16'hC7A3,4);
TASK_PP(16'hC7A4,4);
TASK_PP(16'hC7A5,4);
TASK_PP(16'hC7A6,4);
TASK_PP(16'hC7A7,4);
TASK_PP(16'hC7A8,4);
TASK_PP(16'hC7A9,4);
TASK_PP(16'hC7AA,4);
TASK_PP(16'hC7AB,4);
TASK_PP(16'hC7AC,4);
TASK_PP(16'hC7AD,4);
TASK_PP(16'hC7AE,4);
TASK_PP(16'hC7AF,4);
TASK_PP(16'hC7B0,4);
TASK_PP(16'hC7B1,4);
TASK_PP(16'hC7B2,4);
TASK_PP(16'hC7B3,4);
TASK_PP(16'hC7B4,4);
TASK_PP(16'hC7B5,4);
TASK_PP(16'hC7B6,4);
TASK_PP(16'hC7B7,4);
TASK_PP(16'hC7B8,4);
TASK_PP(16'hC7B9,4);
TASK_PP(16'hC7BA,4);
TASK_PP(16'hC7BB,4);
TASK_PP(16'hC7BC,4);
TASK_PP(16'hC7BD,4);
TASK_PP(16'hC7BE,4);
TASK_PP(16'hC7BF,4);
TASK_PP(16'hC7C0,4);
TASK_PP(16'hC7C1,4);
TASK_PP(16'hC7C2,4);
TASK_PP(16'hC7C3,4);
TASK_PP(16'hC7C4,4);
TASK_PP(16'hC7C5,4);
TASK_PP(16'hC7C6,4);
TASK_PP(16'hC7C7,4);
TASK_PP(16'hC7C8,4);
TASK_PP(16'hC7C9,4);
TASK_PP(16'hC7CA,4);
TASK_PP(16'hC7CB,4);
TASK_PP(16'hC7CC,4);
TASK_PP(16'hC7CD,4);
TASK_PP(16'hC7CE,4);
TASK_PP(16'hC7CF,4);
TASK_PP(16'hC7D0,4);
TASK_PP(16'hC7D1,4);
TASK_PP(16'hC7D2,4);
TASK_PP(16'hC7D3,4);
TASK_PP(16'hC7D4,4);
TASK_PP(16'hC7D5,4);
TASK_PP(16'hC7D6,4);
TASK_PP(16'hC7D7,4);
TASK_PP(16'hC7D8,4);
TASK_PP(16'hC7D9,4);
TASK_PP(16'hC7DA,4);
TASK_PP(16'hC7DB,4);
TASK_PP(16'hC7DC,4);
TASK_PP(16'hC7DD,4);
TASK_PP(16'hC7DE,4);
TASK_PP(16'hC7DF,4);
TASK_PP(16'hC7E0,4);
TASK_PP(16'hC7E1,4);
TASK_PP(16'hC7E2,4);
TASK_PP(16'hC7E3,4);
TASK_PP(16'hC7E4,4);
TASK_PP(16'hC7E5,4);
TASK_PP(16'hC7E6,4);
TASK_PP(16'hC7E7,4);
TASK_PP(16'hC7E8,4);
TASK_PP(16'hC7E9,4);
TASK_PP(16'hC7EA,4);
TASK_PP(16'hC7EB,4);
TASK_PP(16'hC7EC,4);
TASK_PP(16'hC7ED,4);
TASK_PP(16'hC7EE,4);
TASK_PP(16'hC7EF,4);
TASK_PP(16'hC7F0,4);
TASK_PP(16'hC7F1,4);
TASK_PP(16'hC7F2,4);
TASK_PP(16'hC7F3,4);
TASK_PP(16'hC7F4,4);
TASK_PP(16'hC7F5,4);
TASK_PP(16'hC7F6,4);
TASK_PP(16'hC7F7,4);
TASK_PP(16'hC7F8,4);
TASK_PP(16'hC7F9,4);
TASK_PP(16'hC7FA,4);
TASK_PP(16'hC7FB,4);
TASK_PP(16'hC7FC,4);
TASK_PP(16'hC7FD,4);
TASK_PP(16'hC7FE,4);
TASK_PP(16'hC7FF,4);
TASK_PP(16'hC800,4);
TASK_PP(16'hC801,4);
TASK_PP(16'hC802,4);
TASK_PP(16'hC803,4);
TASK_PP(16'hC804,4);
TASK_PP(16'hC805,4);
TASK_PP(16'hC806,4);
TASK_PP(16'hC807,4);
TASK_PP(16'hC808,4);
TASK_PP(16'hC809,4);
TASK_PP(16'hC80A,4);
TASK_PP(16'hC80B,4);
TASK_PP(16'hC80C,4);
TASK_PP(16'hC80D,4);
TASK_PP(16'hC80E,4);
TASK_PP(16'hC80F,4);
TASK_PP(16'hC810,4);
TASK_PP(16'hC811,4);
TASK_PP(16'hC812,4);
TASK_PP(16'hC813,4);
TASK_PP(16'hC814,4);
TASK_PP(16'hC815,4);
TASK_PP(16'hC816,4);
TASK_PP(16'hC817,4);
TASK_PP(16'hC818,4);
TASK_PP(16'hC819,4);
TASK_PP(16'hC81A,4);
TASK_PP(16'hC81B,4);
TASK_PP(16'hC81C,4);
TASK_PP(16'hC81D,4);
TASK_PP(16'hC81E,4);
TASK_PP(16'hC81F,4);
TASK_PP(16'hC820,4);
TASK_PP(16'hC821,4);
TASK_PP(16'hC822,4);
TASK_PP(16'hC823,4);
TASK_PP(16'hC824,4);
TASK_PP(16'hC825,4);
TASK_PP(16'hC826,4);
TASK_PP(16'hC827,4);
TASK_PP(16'hC828,4);
TASK_PP(16'hC829,4);
TASK_PP(16'hC82A,4);
TASK_PP(16'hC82B,4);
TASK_PP(16'hC82C,4);
TASK_PP(16'hC82D,4);
TASK_PP(16'hC82E,4);
TASK_PP(16'hC82F,4);
TASK_PP(16'hC830,4);
TASK_PP(16'hC831,4);
TASK_PP(16'hC832,4);
TASK_PP(16'hC833,4);
TASK_PP(16'hC834,4);
TASK_PP(16'hC835,4);
TASK_PP(16'hC836,4);
TASK_PP(16'hC837,4);
TASK_PP(16'hC838,4);
TASK_PP(16'hC839,4);
TASK_PP(16'hC83A,4);
TASK_PP(16'hC83B,4);
TASK_PP(16'hC83C,4);
TASK_PP(16'hC83D,4);
TASK_PP(16'hC83E,4);
TASK_PP(16'hC83F,4);
TASK_PP(16'hC840,4);
TASK_PP(16'hC841,4);
TASK_PP(16'hC842,4);
TASK_PP(16'hC843,4);
TASK_PP(16'hC844,4);
TASK_PP(16'hC845,4);
TASK_PP(16'hC846,4);
TASK_PP(16'hC847,4);
TASK_PP(16'hC848,4);
TASK_PP(16'hC849,4);
TASK_PP(16'hC84A,4);
TASK_PP(16'hC84B,4);
TASK_PP(16'hC84C,4);
TASK_PP(16'hC84D,4);
TASK_PP(16'hC84E,4);
TASK_PP(16'hC84F,4);
TASK_PP(16'hC850,4);
TASK_PP(16'hC851,4);
TASK_PP(16'hC852,4);
TASK_PP(16'hC853,4);
TASK_PP(16'hC854,4);
TASK_PP(16'hC855,4);
TASK_PP(16'hC856,4);
TASK_PP(16'hC857,4);
TASK_PP(16'hC858,4);
TASK_PP(16'hC859,4);
TASK_PP(16'hC85A,4);
TASK_PP(16'hC85B,4);
TASK_PP(16'hC85C,4);
TASK_PP(16'hC85D,4);
TASK_PP(16'hC85E,4);
TASK_PP(16'hC85F,4);
TASK_PP(16'hC860,4);
TASK_PP(16'hC861,4);
TASK_PP(16'hC862,4);
TASK_PP(16'hC863,4);
TASK_PP(16'hC864,4);
TASK_PP(16'hC865,4);
TASK_PP(16'hC866,4);
TASK_PP(16'hC867,4);
TASK_PP(16'hC868,4);
TASK_PP(16'hC869,4);
TASK_PP(16'hC86A,4);
TASK_PP(16'hC86B,4);
TASK_PP(16'hC86C,4);
TASK_PP(16'hC86D,4);
TASK_PP(16'hC86E,4);
TASK_PP(16'hC86F,4);
TASK_PP(16'hC870,4);
TASK_PP(16'hC871,4);
TASK_PP(16'hC872,4);
TASK_PP(16'hC873,4);
TASK_PP(16'hC874,4);
TASK_PP(16'hC875,4);
TASK_PP(16'hC876,4);
TASK_PP(16'hC877,4);
TASK_PP(16'hC878,4);
TASK_PP(16'hC879,4);
TASK_PP(16'hC87A,4);
TASK_PP(16'hC87B,4);
TASK_PP(16'hC87C,4);
TASK_PP(16'hC87D,4);
TASK_PP(16'hC87E,4);
TASK_PP(16'hC87F,4);
TASK_PP(16'hC880,4);
TASK_PP(16'hC881,4);
TASK_PP(16'hC882,4);
TASK_PP(16'hC883,4);
TASK_PP(16'hC884,4);
TASK_PP(16'hC885,4);
TASK_PP(16'hC886,4);
TASK_PP(16'hC887,4);
TASK_PP(16'hC888,4);
TASK_PP(16'hC889,4);
TASK_PP(16'hC88A,4);
TASK_PP(16'hC88B,4);
TASK_PP(16'hC88C,4);
TASK_PP(16'hC88D,4);
TASK_PP(16'hC88E,4);
TASK_PP(16'hC88F,4);
TASK_PP(16'hC890,4);
TASK_PP(16'hC891,4);
TASK_PP(16'hC892,4);
TASK_PP(16'hC893,4);
TASK_PP(16'hC894,4);
TASK_PP(16'hC895,4);
TASK_PP(16'hC896,4);
TASK_PP(16'hC897,4);
TASK_PP(16'hC898,4);
TASK_PP(16'hC899,4);
TASK_PP(16'hC89A,4);
TASK_PP(16'hC89B,4);
TASK_PP(16'hC89C,4);
TASK_PP(16'hC89D,4);
TASK_PP(16'hC89E,4);
TASK_PP(16'hC89F,4);
TASK_PP(16'hC8A0,4);
TASK_PP(16'hC8A1,4);
TASK_PP(16'hC8A2,4);
TASK_PP(16'hC8A3,4);
TASK_PP(16'hC8A4,4);
TASK_PP(16'hC8A5,4);
TASK_PP(16'hC8A6,4);
TASK_PP(16'hC8A7,4);
TASK_PP(16'hC8A8,4);
TASK_PP(16'hC8A9,4);
TASK_PP(16'hC8AA,4);
TASK_PP(16'hC8AB,4);
TASK_PP(16'hC8AC,4);
TASK_PP(16'hC8AD,4);
TASK_PP(16'hC8AE,4);
TASK_PP(16'hC8AF,4);
TASK_PP(16'hC8B0,4);
TASK_PP(16'hC8B1,4);
TASK_PP(16'hC8B2,4);
TASK_PP(16'hC8B3,4);
TASK_PP(16'hC8B4,4);
TASK_PP(16'hC8B5,4);
TASK_PP(16'hC8B6,4);
TASK_PP(16'hC8B7,4);
TASK_PP(16'hC8B8,4);
TASK_PP(16'hC8B9,4);
TASK_PP(16'hC8BA,4);
TASK_PP(16'hC8BB,4);
TASK_PP(16'hC8BC,4);
TASK_PP(16'hC8BD,4);
TASK_PP(16'hC8BE,4);
TASK_PP(16'hC8BF,4);
TASK_PP(16'hC8C0,4);
TASK_PP(16'hC8C1,4);
TASK_PP(16'hC8C2,4);
TASK_PP(16'hC8C3,4);
TASK_PP(16'hC8C4,4);
TASK_PP(16'hC8C5,4);
TASK_PP(16'hC8C6,4);
TASK_PP(16'hC8C7,4);
TASK_PP(16'hC8C8,4);
TASK_PP(16'hC8C9,4);
TASK_PP(16'hC8CA,4);
TASK_PP(16'hC8CB,4);
TASK_PP(16'hC8CC,4);
TASK_PP(16'hC8CD,4);
TASK_PP(16'hC8CE,4);
TASK_PP(16'hC8CF,4);
TASK_PP(16'hC8D0,4);
TASK_PP(16'hC8D1,4);
TASK_PP(16'hC8D2,4);
TASK_PP(16'hC8D3,4);
TASK_PP(16'hC8D4,4);
TASK_PP(16'hC8D5,4);
TASK_PP(16'hC8D6,4);
TASK_PP(16'hC8D7,4);
TASK_PP(16'hC8D8,4);
TASK_PP(16'hC8D9,4);
TASK_PP(16'hC8DA,4);
TASK_PP(16'hC8DB,4);
TASK_PP(16'hC8DC,4);
TASK_PP(16'hC8DD,4);
TASK_PP(16'hC8DE,4);
TASK_PP(16'hC8DF,4);
TASK_PP(16'hC8E0,4);
TASK_PP(16'hC8E1,4);
TASK_PP(16'hC8E2,4);
TASK_PP(16'hC8E3,4);
TASK_PP(16'hC8E4,4);
TASK_PP(16'hC8E5,4);
TASK_PP(16'hC8E6,4);
TASK_PP(16'hC8E7,4);
TASK_PP(16'hC8E8,4);
TASK_PP(16'hC8E9,4);
TASK_PP(16'hC8EA,4);
TASK_PP(16'hC8EB,4);
TASK_PP(16'hC8EC,4);
TASK_PP(16'hC8ED,4);
TASK_PP(16'hC8EE,4);
TASK_PP(16'hC8EF,4);
TASK_PP(16'hC8F0,4);
TASK_PP(16'hC8F1,4);
TASK_PP(16'hC8F2,4);
TASK_PP(16'hC8F3,4);
TASK_PP(16'hC8F4,4);
TASK_PP(16'hC8F5,4);
TASK_PP(16'hC8F6,4);
TASK_PP(16'hC8F7,4);
TASK_PP(16'hC8F8,4);
TASK_PP(16'hC8F9,4);
TASK_PP(16'hC8FA,4);
TASK_PP(16'hC8FB,4);
TASK_PP(16'hC8FC,4);
TASK_PP(16'hC8FD,4);
TASK_PP(16'hC8FE,4);
TASK_PP(16'hC8FF,4);
TASK_PP(16'hC900,4);
TASK_PP(16'hC901,4);
TASK_PP(16'hC902,4);
TASK_PP(16'hC903,4);
TASK_PP(16'hC904,4);
TASK_PP(16'hC905,4);
TASK_PP(16'hC906,4);
TASK_PP(16'hC907,4);
TASK_PP(16'hC908,4);
TASK_PP(16'hC909,4);
TASK_PP(16'hC90A,4);
TASK_PP(16'hC90B,4);
TASK_PP(16'hC90C,4);
TASK_PP(16'hC90D,4);
TASK_PP(16'hC90E,4);
TASK_PP(16'hC90F,4);
TASK_PP(16'hC910,4);
TASK_PP(16'hC911,4);
TASK_PP(16'hC912,4);
TASK_PP(16'hC913,4);
TASK_PP(16'hC914,4);
TASK_PP(16'hC915,4);
TASK_PP(16'hC916,4);
TASK_PP(16'hC917,4);
TASK_PP(16'hC918,4);
TASK_PP(16'hC919,4);
TASK_PP(16'hC91A,4);
TASK_PP(16'hC91B,4);
TASK_PP(16'hC91C,4);
TASK_PP(16'hC91D,4);
TASK_PP(16'hC91E,4);
TASK_PP(16'hC91F,4);
TASK_PP(16'hC920,4);
TASK_PP(16'hC921,4);
TASK_PP(16'hC922,4);
TASK_PP(16'hC923,4);
TASK_PP(16'hC924,4);
TASK_PP(16'hC925,4);
TASK_PP(16'hC926,4);
TASK_PP(16'hC927,4);
TASK_PP(16'hC928,4);
TASK_PP(16'hC929,4);
TASK_PP(16'hC92A,4);
TASK_PP(16'hC92B,4);
TASK_PP(16'hC92C,4);
TASK_PP(16'hC92D,4);
TASK_PP(16'hC92E,4);
TASK_PP(16'hC92F,4);
TASK_PP(16'hC930,4);
TASK_PP(16'hC931,4);
TASK_PP(16'hC932,4);
TASK_PP(16'hC933,4);
TASK_PP(16'hC934,4);
TASK_PP(16'hC935,4);
TASK_PP(16'hC936,4);
TASK_PP(16'hC937,4);
TASK_PP(16'hC938,4);
TASK_PP(16'hC939,4);
TASK_PP(16'hC93A,4);
TASK_PP(16'hC93B,4);
TASK_PP(16'hC93C,4);
TASK_PP(16'hC93D,4);
TASK_PP(16'hC93E,4);
TASK_PP(16'hC93F,4);
TASK_PP(16'hC940,4);
TASK_PP(16'hC941,4);
TASK_PP(16'hC942,4);
TASK_PP(16'hC943,4);
TASK_PP(16'hC944,4);
TASK_PP(16'hC945,4);
TASK_PP(16'hC946,4);
TASK_PP(16'hC947,4);
TASK_PP(16'hC948,4);
TASK_PP(16'hC949,4);
TASK_PP(16'hC94A,4);
TASK_PP(16'hC94B,4);
TASK_PP(16'hC94C,4);
TASK_PP(16'hC94D,4);
TASK_PP(16'hC94E,4);
TASK_PP(16'hC94F,4);
TASK_PP(16'hC950,4);
TASK_PP(16'hC951,4);
TASK_PP(16'hC952,4);
TASK_PP(16'hC953,4);
TASK_PP(16'hC954,4);
TASK_PP(16'hC955,4);
TASK_PP(16'hC956,4);
TASK_PP(16'hC957,4);
TASK_PP(16'hC958,4);
TASK_PP(16'hC959,4);
TASK_PP(16'hC95A,4);
TASK_PP(16'hC95B,4);
TASK_PP(16'hC95C,4);
TASK_PP(16'hC95D,4);
TASK_PP(16'hC95E,4);
TASK_PP(16'hC95F,4);
TASK_PP(16'hC960,4);
TASK_PP(16'hC961,4);
TASK_PP(16'hC962,4);
TASK_PP(16'hC963,4);
TASK_PP(16'hC964,4);
TASK_PP(16'hC965,4);
TASK_PP(16'hC966,4);
TASK_PP(16'hC967,4);
TASK_PP(16'hC968,4);
TASK_PP(16'hC969,4);
TASK_PP(16'hC96A,4);
TASK_PP(16'hC96B,4);
TASK_PP(16'hC96C,4);
TASK_PP(16'hC96D,4);
TASK_PP(16'hC96E,4);
TASK_PP(16'hC96F,4);
TASK_PP(16'hC970,4);
TASK_PP(16'hC971,4);
TASK_PP(16'hC972,4);
TASK_PP(16'hC973,4);
TASK_PP(16'hC974,4);
TASK_PP(16'hC975,4);
TASK_PP(16'hC976,4);
TASK_PP(16'hC977,4);
TASK_PP(16'hC978,4);
TASK_PP(16'hC979,4);
TASK_PP(16'hC97A,4);
TASK_PP(16'hC97B,4);
TASK_PP(16'hC97C,4);
TASK_PP(16'hC97D,4);
TASK_PP(16'hC97E,4);
TASK_PP(16'hC97F,4);
TASK_PP(16'hC980,4);
TASK_PP(16'hC981,4);
TASK_PP(16'hC982,4);
TASK_PP(16'hC983,4);
TASK_PP(16'hC984,4);
TASK_PP(16'hC985,4);
TASK_PP(16'hC986,4);
TASK_PP(16'hC987,4);
TASK_PP(16'hC988,4);
TASK_PP(16'hC989,4);
TASK_PP(16'hC98A,4);
TASK_PP(16'hC98B,4);
TASK_PP(16'hC98C,4);
TASK_PP(16'hC98D,4);
TASK_PP(16'hC98E,4);
TASK_PP(16'hC98F,4);
TASK_PP(16'hC990,4);
TASK_PP(16'hC991,4);
TASK_PP(16'hC992,4);
TASK_PP(16'hC993,4);
TASK_PP(16'hC994,4);
TASK_PP(16'hC995,4);
TASK_PP(16'hC996,4);
TASK_PP(16'hC997,4);
TASK_PP(16'hC998,4);
TASK_PP(16'hC999,4);
TASK_PP(16'hC99A,4);
TASK_PP(16'hC99B,4);
TASK_PP(16'hC99C,4);
TASK_PP(16'hC99D,4);
TASK_PP(16'hC99E,4);
TASK_PP(16'hC99F,4);
TASK_PP(16'hC9A0,4);
TASK_PP(16'hC9A1,4);
TASK_PP(16'hC9A2,4);
TASK_PP(16'hC9A3,4);
TASK_PP(16'hC9A4,4);
TASK_PP(16'hC9A5,4);
TASK_PP(16'hC9A6,4);
TASK_PP(16'hC9A7,4);
TASK_PP(16'hC9A8,4);
TASK_PP(16'hC9A9,4);
TASK_PP(16'hC9AA,4);
TASK_PP(16'hC9AB,4);
TASK_PP(16'hC9AC,4);
TASK_PP(16'hC9AD,4);
TASK_PP(16'hC9AE,4);
TASK_PP(16'hC9AF,4);
TASK_PP(16'hC9B0,4);
TASK_PP(16'hC9B1,4);
TASK_PP(16'hC9B2,4);
TASK_PP(16'hC9B3,4);
TASK_PP(16'hC9B4,4);
TASK_PP(16'hC9B5,4);
TASK_PP(16'hC9B6,4);
TASK_PP(16'hC9B7,4);
TASK_PP(16'hC9B8,4);
TASK_PP(16'hC9B9,4);
TASK_PP(16'hC9BA,4);
TASK_PP(16'hC9BB,4);
TASK_PP(16'hC9BC,4);
TASK_PP(16'hC9BD,4);
TASK_PP(16'hC9BE,4);
TASK_PP(16'hC9BF,4);
TASK_PP(16'hC9C0,4);
TASK_PP(16'hC9C1,4);
TASK_PP(16'hC9C2,4);
TASK_PP(16'hC9C3,4);
TASK_PP(16'hC9C4,4);
TASK_PP(16'hC9C5,4);
TASK_PP(16'hC9C6,4);
TASK_PP(16'hC9C7,4);
TASK_PP(16'hC9C8,4);
TASK_PP(16'hC9C9,4);
TASK_PP(16'hC9CA,4);
TASK_PP(16'hC9CB,4);
TASK_PP(16'hC9CC,4);
TASK_PP(16'hC9CD,4);
TASK_PP(16'hC9CE,4);
TASK_PP(16'hC9CF,4);
TASK_PP(16'hC9D0,4);
TASK_PP(16'hC9D1,4);
TASK_PP(16'hC9D2,4);
TASK_PP(16'hC9D3,4);
TASK_PP(16'hC9D4,4);
TASK_PP(16'hC9D5,4);
TASK_PP(16'hC9D6,4);
TASK_PP(16'hC9D7,4);
TASK_PP(16'hC9D8,4);
TASK_PP(16'hC9D9,4);
TASK_PP(16'hC9DA,4);
TASK_PP(16'hC9DB,4);
TASK_PP(16'hC9DC,4);
TASK_PP(16'hC9DD,4);
TASK_PP(16'hC9DE,4);
TASK_PP(16'hC9DF,4);
TASK_PP(16'hC9E0,4);
TASK_PP(16'hC9E1,4);
TASK_PP(16'hC9E2,4);
TASK_PP(16'hC9E3,4);
TASK_PP(16'hC9E4,4);
TASK_PP(16'hC9E5,4);
TASK_PP(16'hC9E6,4);
TASK_PP(16'hC9E7,4);
TASK_PP(16'hC9E8,4);
TASK_PP(16'hC9E9,4);
TASK_PP(16'hC9EA,4);
TASK_PP(16'hC9EB,4);
TASK_PP(16'hC9EC,4);
TASK_PP(16'hC9ED,4);
TASK_PP(16'hC9EE,4);
TASK_PP(16'hC9EF,4);
TASK_PP(16'hC9F0,4);
TASK_PP(16'hC9F1,4);
TASK_PP(16'hC9F2,4);
TASK_PP(16'hC9F3,4);
TASK_PP(16'hC9F4,4);
TASK_PP(16'hC9F5,4);
TASK_PP(16'hC9F6,4);
TASK_PP(16'hC9F7,4);
TASK_PP(16'hC9F8,4);
TASK_PP(16'hC9F9,4);
TASK_PP(16'hC9FA,4);
TASK_PP(16'hC9FB,4);
TASK_PP(16'hC9FC,4);
TASK_PP(16'hC9FD,4);
TASK_PP(16'hC9FE,4);
TASK_PP(16'hC9FF,4);
TASK_PP(16'hCA00,4);
TASK_PP(16'hCA01,4);
TASK_PP(16'hCA02,4);
TASK_PP(16'hCA03,4);
TASK_PP(16'hCA04,4);
TASK_PP(16'hCA05,4);
TASK_PP(16'hCA06,4);
TASK_PP(16'hCA07,4);
TASK_PP(16'hCA08,4);
TASK_PP(16'hCA09,4);
TASK_PP(16'hCA0A,4);
TASK_PP(16'hCA0B,4);
TASK_PP(16'hCA0C,4);
TASK_PP(16'hCA0D,4);
TASK_PP(16'hCA0E,4);
TASK_PP(16'hCA0F,4);
TASK_PP(16'hCA10,4);
TASK_PP(16'hCA11,4);
TASK_PP(16'hCA12,4);
TASK_PP(16'hCA13,4);
TASK_PP(16'hCA14,4);
TASK_PP(16'hCA15,4);
TASK_PP(16'hCA16,4);
TASK_PP(16'hCA17,4);
TASK_PP(16'hCA18,4);
TASK_PP(16'hCA19,4);
TASK_PP(16'hCA1A,4);
TASK_PP(16'hCA1B,4);
TASK_PP(16'hCA1C,4);
TASK_PP(16'hCA1D,4);
TASK_PP(16'hCA1E,4);
TASK_PP(16'hCA1F,4);
TASK_PP(16'hCA20,4);
TASK_PP(16'hCA21,4);
TASK_PP(16'hCA22,4);
TASK_PP(16'hCA23,4);
TASK_PP(16'hCA24,4);
TASK_PP(16'hCA25,4);
TASK_PP(16'hCA26,4);
TASK_PP(16'hCA27,4);
TASK_PP(16'hCA28,4);
TASK_PP(16'hCA29,4);
TASK_PP(16'hCA2A,4);
TASK_PP(16'hCA2B,4);
TASK_PP(16'hCA2C,4);
TASK_PP(16'hCA2D,4);
TASK_PP(16'hCA2E,4);
TASK_PP(16'hCA2F,4);
TASK_PP(16'hCA30,4);
TASK_PP(16'hCA31,4);
TASK_PP(16'hCA32,4);
TASK_PP(16'hCA33,4);
TASK_PP(16'hCA34,4);
TASK_PP(16'hCA35,4);
TASK_PP(16'hCA36,4);
TASK_PP(16'hCA37,4);
TASK_PP(16'hCA38,4);
TASK_PP(16'hCA39,4);
TASK_PP(16'hCA3A,4);
TASK_PP(16'hCA3B,4);
TASK_PP(16'hCA3C,4);
TASK_PP(16'hCA3D,4);
TASK_PP(16'hCA3E,4);
TASK_PP(16'hCA3F,4);
TASK_PP(16'hCA40,4);
TASK_PP(16'hCA41,4);
TASK_PP(16'hCA42,4);
TASK_PP(16'hCA43,4);
TASK_PP(16'hCA44,4);
TASK_PP(16'hCA45,4);
TASK_PP(16'hCA46,4);
TASK_PP(16'hCA47,4);
TASK_PP(16'hCA48,4);
TASK_PP(16'hCA49,4);
TASK_PP(16'hCA4A,4);
TASK_PP(16'hCA4B,4);
TASK_PP(16'hCA4C,4);
TASK_PP(16'hCA4D,4);
TASK_PP(16'hCA4E,4);
TASK_PP(16'hCA4F,4);
TASK_PP(16'hCA50,4);
TASK_PP(16'hCA51,4);
TASK_PP(16'hCA52,4);
TASK_PP(16'hCA53,4);
TASK_PP(16'hCA54,4);
TASK_PP(16'hCA55,4);
TASK_PP(16'hCA56,4);
TASK_PP(16'hCA57,4);
TASK_PP(16'hCA58,4);
TASK_PP(16'hCA59,4);
TASK_PP(16'hCA5A,4);
TASK_PP(16'hCA5B,4);
TASK_PP(16'hCA5C,4);
TASK_PP(16'hCA5D,4);
TASK_PP(16'hCA5E,4);
TASK_PP(16'hCA5F,4);
TASK_PP(16'hCA60,4);
TASK_PP(16'hCA61,4);
TASK_PP(16'hCA62,4);
TASK_PP(16'hCA63,4);
TASK_PP(16'hCA64,4);
TASK_PP(16'hCA65,4);
TASK_PP(16'hCA66,4);
TASK_PP(16'hCA67,4);
TASK_PP(16'hCA68,4);
TASK_PP(16'hCA69,4);
TASK_PP(16'hCA6A,4);
TASK_PP(16'hCA6B,4);
TASK_PP(16'hCA6C,4);
TASK_PP(16'hCA6D,4);
TASK_PP(16'hCA6E,4);
TASK_PP(16'hCA6F,4);
TASK_PP(16'hCA70,4);
TASK_PP(16'hCA71,4);
TASK_PP(16'hCA72,4);
TASK_PP(16'hCA73,4);
TASK_PP(16'hCA74,4);
TASK_PP(16'hCA75,4);
TASK_PP(16'hCA76,4);
TASK_PP(16'hCA77,4);
TASK_PP(16'hCA78,4);
TASK_PP(16'hCA79,4);
TASK_PP(16'hCA7A,4);
TASK_PP(16'hCA7B,4);
TASK_PP(16'hCA7C,4);
TASK_PP(16'hCA7D,4);
TASK_PP(16'hCA7E,4);
TASK_PP(16'hCA7F,4);
TASK_PP(16'hCA80,4);
TASK_PP(16'hCA81,4);
TASK_PP(16'hCA82,4);
TASK_PP(16'hCA83,4);
TASK_PP(16'hCA84,4);
TASK_PP(16'hCA85,4);
TASK_PP(16'hCA86,4);
TASK_PP(16'hCA87,4);
TASK_PP(16'hCA88,4);
TASK_PP(16'hCA89,4);
TASK_PP(16'hCA8A,4);
TASK_PP(16'hCA8B,4);
TASK_PP(16'hCA8C,4);
TASK_PP(16'hCA8D,4);
TASK_PP(16'hCA8E,4);
TASK_PP(16'hCA8F,4);
TASK_PP(16'hCA90,4);
TASK_PP(16'hCA91,4);
TASK_PP(16'hCA92,4);
TASK_PP(16'hCA93,4);
TASK_PP(16'hCA94,4);
TASK_PP(16'hCA95,4);
TASK_PP(16'hCA96,4);
TASK_PP(16'hCA97,4);
TASK_PP(16'hCA98,4);
TASK_PP(16'hCA99,4);
TASK_PP(16'hCA9A,4);
TASK_PP(16'hCA9B,4);
TASK_PP(16'hCA9C,4);
TASK_PP(16'hCA9D,4);
TASK_PP(16'hCA9E,4);
TASK_PP(16'hCA9F,4);
TASK_PP(16'hCAA0,4);
TASK_PP(16'hCAA1,4);
TASK_PP(16'hCAA2,4);
TASK_PP(16'hCAA3,4);
TASK_PP(16'hCAA4,4);
TASK_PP(16'hCAA5,4);
TASK_PP(16'hCAA6,4);
TASK_PP(16'hCAA7,4);
TASK_PP(16'hCAA8,4);
TASK_PP(16'hCAA9,4);
TASK_PP(16'hCAAA,4);
TASK_PP(16'hCAAB,4);
TASK_PP(16'hCAAC,4);
TASK_PP(16'hCAAD,4);
TASK_PP(16'hCAAE,4);
TASK_PP(16'hCAAF,4);
TASK_PP(16'hCAB0,4);
TASK_PP(16'hCAB1,4);
TASK_PP(16'hCAB2,4);
TASK_PP(16'hCAB3,4);
TASK_PP(16'hCAB4,4);
TASK_PP(16'hCAB5,4);
TASK_PP(16'hCAB6,4);
TASK_PP(16'hCAB7,4);
TASK_PP(16'hCAB8,4);
TASK_PP(16'hCAB9,4);
TASK_PP(16'hCABA,4);
TASK_PP(16'hCABB,4);
TASK_PP(16'hCABC,4);
TASK_PP(16'hCABD,4);
TASK_PP(16'hCABE,4);
TASK_PP(16'hCABF,4);
TASK_PP(16'hCAC0,4);
TASK_PP(16'hCAC1,4);
TASK_PP(16'hCAC2,4);
TASK_PP(16'hCAC3,4);
TASK_PP(16'hCAC4,4);
TASK_PP(16'hCAC5,4);
TASK_PP(16'hCAC6,4);
TASK_PP(16'hCAC7,4);
TASK_PP(16'hCAC8,4);
TASK_PP(16'hCAC9,4);
TASK_PP(16'hCACA,4);
TASK_PP(16'hCACB,4);
TASK_PP(16'hCACC,4);
TASK_PP(16'hCACD,4);
TASK_PP(16'hCACE,4);
TASK_PP(16'hCACF,4);
TASK_PP(16'hCAD0,4);
TASK_PP(16'hCAD1,4);
TASK_PP(16'hCAD2,4);
TASK_PP(16'hCAD3,4);
TASK_PP(16'hCAD4,4);
TASK_PP(16'hCAD5,4);
TASK_PP(16'hCAD6,4);
TASK_PP(16'hCAD7,4);
TASK_PP(16'hCAD8,4);
TASK_PP(16'hCAD9,4);
TASK_PP(16'hCADA,4);
TASK_PP(16'hCADB,4);
TASK_PP(16'hCADC,4);
TASK_PP(16'hCADD,4);
TASK_PP(16'hCADE,4);
TASK_PP(16'hCADF,4);
TASK_PP(16'hCAE0,4);
TASK_PP(16'hCAE1,4);
TASK_PP(16'hCAE2,4);
TASK_PP(16'hCAE3,4);
TASK_PP(16'hCAE4,4);
TASK_PP(16'hCAE5,4);
TASK_PP(16'hCAE6,4);
TASK_PP(16'hCAE7,4);
TASK_PP(16'hCAE8,4);
TASK_PP(16'hCAE9,4);
TASK_PP(16'hCAEA,4);
TASK_PP(16'hCAEB,4);
TASK_PP(16'hCAEC,4);
TASK_PP(16'hCAED,4);
TASK_PP(16'hCAEE,4);
TASK_PP(16'hCAEF,4);
TASK_PP(16'hCAF0,4);
TASK_PP(16'hCAF1,4);
TASK_PP(16'hCAF2,4);
TASK_PP(16'hCAF3,4);
TASK_PP(16'hCAF4,4);
TASK_PP(16'hCAF5,4);
TASK_PP(16'hCAF6,4);
TASK_PP(16'hCAF7,4);
TASK_PP(16'hCAF8,4);
TASK_PP(16'hCAF9,4);
TASK_PP(16'hCAFA,4);
TASK_PP(16'hCAFB,4);
TASK_PP(16'hCAFC,4);
TASK_PP(16'hCAFD,4);
TASK_PP(16'hCAFE,4);
TASK_PP(16'hCAFF,4);
TASK_PP(16'hCB00,4);
TASK_PP(16'hCB01,4);
TASK_PP(16'hCB02,4);
TASK_PP(16'hCB03,4);
TASK_PP(16'hCB04,4);
TASK_PP(16'hCB05,4);
TASK_PP(16'hCB06,4);
TASK_PP(16'hCB07,4);
TASK_PP(16'hCB08,4);
TASK_PP(16'hCB09,4);
TASK_PP(16'hCB0A,4);
TASK_PP(16'hCB0B,4);
TASK_PP(16'hCB0C,4);
TASK_PP(16'hCB0D,4);
TASK_PP(16'hCB0E,4);
TASK_PP(16'hCB0F,4);
TASK_PP(16'hCB10,4);
TASK_PP(16'hCB11,4);
TASK_PP(16'hCB12,4);
TASK_PP(16'hCB13,4);
TASK_PP(16'hCB14,4);
TASK_PP(16'hCB15,4);
TASK_PP(16'hCB16,4);
TASK_PP(16'hCB17,4);
TASK_PP(16'hCB18,4);
TASK_PP(16'hCB19,4);
TASK_PP(16'hCB1A,4);
TASK_PP(16'hCB1B,4);
TASK_PP(16'hCB1C,4);
TASK_PP(16'hCB1D,4);
TASK_PP(16'hCB1E,4);
TASK_PP(16'hCB1F,4);
TASK_PP(16'hCB20,4);
TASK_PP(16'hCB21,4);
TASK_PP(16'hCB22,4);
TASK_PP(16'hCB23,4);
TASK_PP(16'hCB24,4);
TASK_PP(16'hCB25,4);
TASK_PP(16'hCB26,4);
TASK_PP(16'hCB27,4);
TASK_PP(16'hCB28,4);
TASK_PP(16'hCB29,4);
TASK_PP(16'hCB2A,4);
TASK_PP(16'hCB2B,4);
TASK_PP(16'hCB2C,4);
TASK_PP(16'hCB2D,4);
TASK_PP(16'hCB2E,4);
TASK_PP(16'hCB2F,4);
TASK_PP(16'hCB30,4);
TASK_PP(16'hCB31,4);
TASK_PP(16'hCB32,4);
TASK_PP(16'hCB33,4);
TASK_PP(16'hCB34,4);
TASK_PP(16'hCB35,4);
TASK_PP(16'hCB36,4);
TASK_PP(16'hCB37,4);
TASK_PP(16'hCB38,4);
TASK_PP(16'hCB39,4);
TASK_PP(16'hCB3A,4);
TASK_PP(16'hCB3B,4);
TASK_PP(16'hCB3C,4);
TASK_PP(16'hCB3D,4);
TASK_PP(16'hCB3E,4);
TASK_PP(16'hCB3F,4);
TASK_PP(16'hCB40,4);
TASK_PP(16'hCB41,4);
TASK_PP(16'hCB42,4);
TASK_PP(16'hCB43,4);
TASK_PP(16'hCB44,4);
TASK_PP(16'hCB45,4);
TASK_PP(16'hCB46,4);
TASK_PP(16'hCB47,4);
TASK_PP(16'hCB48,4);
TASK_PP(16'hCB49,4);
TASK_PP(16'hCB4A,4);
TASK_PP(16'hCB4B,4);
TASK_PP(16'hCB4C,4);
TASK_PP(16'hCB4D,4);
TASK_PP(16'hCB4E,4);
TASK_PP(16'hCB4F,4);
TASK_PP(16'hCB50,4);
TASK_PP(16'hCB51,4);
TASK_PP(16'hCB52,4);
TASK_PP(16'hCB53,4);
TASK_PP(16'hCB54,4);
TASK_PP(16'hCB55,4);
TASK_PP(16'hCB56,4);
TASK_PP(16'hCB57,4);
TASK_PP(16'hCB58,4);
TASK_PP(16'hCB59,4);
TASK_PP(16'hCB5A,4);
TASK_PP(16'hCB5B,4);
TASK_PP(16'hCB5C,4);
TASK_PP(16'hCB5D,4);
TASK_PP(16'hCB5E,4);
TASK_PP(16'hCB5F,4);
TASK_PP(16'hCB60,4);
TASK_PP(16'hCB61,4);
TASK_PP(16'hCB62,4);
TASK_PP(16'hCB63,4);
TASK_PP(16'hCB64,4);
TASK_PP(16'hCB65,4);
TASK_PP(16'hCB66,4);
TASK_PP(16'hCB67,4);
TASK_PP(16'hCB68,4);
TASK_PP(16'hCB69,4);
TASK_PP(16'hCB6A,4);
TASK_PP(16'hCB6B,4);
TASK_PP(16'hCB6C,4);
TASK_PP(16'hCB6D,4);
TASK_PP(16'hCB6E,4);
TASK_PP(16'hCB6F,4);
TASK_PP(16'hCB70,4);
TASK_PP(16'hCB71,4);
TASK_PP(16'hCB72,4);
TASK_PP(16'hCB73,4);
TASK_PP(16'hCB74,4);
TASK_PP(16'hCB75,4);
TASK_PP(16'hCB76,4);
TASK_PP(16'hCB77,4);
TASK_PP(16'hCB78,4);
TASK_PP(16'hCB79,4);
TASK_PP(16'hCB7A,4);
TASK_PP(16'hCB7B,4);
TASK_PP(16'hCB7C,4);
TASK_PP(16'hCB7D,4);
TASK_PP(16'hCB7E,4);
TASK_PP(16'hCB7F,4);
TASK_PP(16'hCB80,4);
TASK_PP(16'hCB81,4);
TASK_PP(16'hCB82,4);
TASK_PP(16'hCB83,4);
TASK_PP(16'hCB84,4);
TASK_PP(16'hCB85,4);
TASK_PP(16'hCB86,4);
TASK_PP(16'hCB87,4);
TASK_PP(16'hCB88,4);
TASK_PP(16'hCB89,4);
TASK_PP(16'hCB8A,4);
TASK_PP(16'hCB8B,4);
TASK_PP(16'hCB8C,4);
TASK_PP(16'hCB8D,4);
TASK_PP(16'hCB8E,4);
TASK_PP(16'hCB8F,4);
TASK_PP(16'hCB90,4);
TASK_PP(16'hCB91,4);
TASK_PP(16'hCB92,4);
TASK_PP(16'hCB93,4);
TASK_PP(16'hCB94,4);
TASK_PP(16'hCB95,4);
TASK_PP(16'hCB96,4);
TASK_PP(16'hCB97,4);
TASK_PP(16'hCB98,4);
TASK_PP(16'hCB99,4);
TASK_PP(16'hCB9A,4);
TASK_PP(16'hCB9B,4);
TASK_PP(16'hCB9C,4);
TASK_PP(16'hCB9D,4);
TASK_PP(16'hCB9E,4);
TASK_PP(16'hCB9F,4);
TASK_PP(16'hCBA0,4);
TASK_PP(16'hCBA1,4);
TASK_PP(16'hCBA2,4);
TASK_PP(16'hCBA3,4);
TASK_PP(16'hCBA4,4);
TASK_PP(16'hCBA5,4);
TASK_PP(16'hCBA6,4);
TASK_PP(16'hCBA7,4);
TASK_PP(16'hCBA8,4);
TASK_PP(16'hCBA9,4);
TASK_PP(16'hCBAA,4);
TASK_PP(16'hCBAB,4);
TASK_PP(16'hCBAC,4);
TASK_PP(16'hCBAD,4);
TASK_PP(16'hCBAE,4);
TASK_PP(16'hCBAF,4);
TASK_PP(16'hCBB0,4);
TASK_PP(16'hCBB1,4);
TASK_PP(16'hCBB2,4);
TASK_PP(16'hCBB3,4);
TASK_PP(16'hCBB4,4);
TASK_PP(16'hCBB5,4);
TASK_PP(16'hCBB6,4);
TASK_PP(16'hCBB7,4);
TASK_PP(16'hCBB8,4);
TASK_PP(16'hCBB9,4);
TASK_PP(16'hCBBA,4);
TASK_PP(16'hCBBB,4);
TASK_PP(16'hCBBC,4);
TASK_PP(16'hCBBD,4);
TASK_PP(16'hCBBE,4);
TASK_PP(16'hCBBF,4);
TASK_PP(16'hCBC0,4);
TASK_PP(16'hCBC1,4);
TASK_PP(16'hCBC2,4);
TASK_PP(16'hCBC3,4);
TASK_PP(16'hCBC4,4);
TASK_PP(16'hCBC5,4);
TASK_PP(16'hCBC6,4);
TASK_PP(16'hCBC7,4);
TASK_PP(16'hCBC8,4);
TASK_PP(16'hCBC9,4);
TASK_PP(16'hCBCA,4);
TASK_PP(16'hCBCB,4);
TASK_PP(16'hCBCC,4);
TASK_PP(16'hCBCD,4);
TASK_PP(16'hCBCE,4);
TASK_PP(16'hCBCF,4);
TASK_PP(16'hCBD0,4);
TASK_PP(16'hCBD1,4);
TASK_PP(16'hCBD2,4);
TASK_PP(16'hCBD3,4);
TASK_PP(16'hCBD4,4);
TASK_PP(16'hCBD5,4);
TASK_PP(16'hCBD6,4);
TASK_PP(16'hCBD7,4);
TASK_PP(16'hCBD8,4);
TASK_PP(16'hCBD9,4);
TASK_PP(16'hCBDA,4);
TASK_PP(16'hCBDB,4);
TASK_PP(16'hCBDC,4);
TASK_PP(16'hCBDD,4);
TASK_PP(16'hCBDE,4);
TASK_PP(16'hCBDF,4);
TASK_PP(16'hCBE0,4);
TASK_PP(16'hCBE1,4);
TASK_PP(16'hCBE2,4);
TASK_PP(16'hCBE3,4);
TASK_PP(16'hCBE4,4);
TASK_PP(16'hCBE5,4);
TASK_PP(16'hCBE6,4);
TASK_PP(16'hCBE7,4);
TASK_PP(16'hCBE8,4);
TASK_PP(16'hCBE9,4);
TASK_PP(16'hCBEA,4);
TASK_PP(16'hCBEB,4);
TASK_PP(16'hCBEC,4);
TASK_PP(16'hCBED,4);
TASK_PP(16'hCBEE,4);
TASK_PP(16'hCBEF,4);
TASK_PP(16'hCBF0,4);
TASK_PP(16'hCBF1,4);
TASK_PP(16'hCBF2,4);
TASK_PP(16'hCBF3,4);
TASK_PP(16'hCBF4,4);
TASK_PP(16'hCBF5,4);
TASK_PP(16'hCBF6,4);
TASK_PP(16'hCBF7,4);
TASK_PP(16'hCBF8,4);
TASK_PP(16'hCBF9,4);
TASK_PP(16'hCBFA,4);
TASK_PP(16'hCBFB,4);
TASK_PP(16'hCBFC,4);
TASK_PP(16'hCBFD,4);
TASK_PP(16'hCBFE,4);
TASK_PP(16'hCBFF,4);
TASK_PP(16'hCC00,4);
TASK_PP(16'hCC01,4);
TASK_PP(16'hCC02,4);
TASK_PP(16'hCC03,4);
TASK_PP(16'hCC04,4);
TASK_PP(16'hCC05,4);
TASK_PP(16'hCC06,4);
TASK_PP(16'hCC07,4);
TASK_PP(16'hCC08,4);
TASK_PP(16'hCC09,4);
TASK_PP(16'hCC0A,4);
TASK_PP(16'hCC0B,4);
TASK_PP(16'hCC0C,4);
TASK_PP(16'hCC0D,4);
TASK_PP(16'hCC0E,4);
TASK_PP(16'hCC0F,4);
TASK_PP(16'hCC10,4);
TASK_PP(16'hCC11,4);
TASK_PP(16'hCC12,4);
TASK_PP(16'hCC13,4);
TASK_PP(16'hCC14,4);
TASK_PP(16'hCC15,4);
TASK_PP(16'hCC16,4);
TASK_PP(16'hCC17,4);
TASK_PP(16'hCC18,4);
TASK_PP(16'hCC19,4);
TASK_PP(16'hCC1A,4);
TASK_PP(16'hCC1B,4);
TASK_PP(16'hCC1C,4);
TASK_PP(16'hCC1D,4);
TASK_PP(16'hCC1E,4);
TASK_PP(16'hCC1F,4);
TASK_PP(16'hCC20,4);
TASK_PP(16'hCC21,4);
TASK_PP(16'hCC22,4);
TASK_PP(16'hCC23,4);
TASK_PP(16'hCC24,4);
TASK_PP(16'hCC25,4);
TASK_PP(16'hCC26,4);
TASK_PP(16'hCC27,4);
TASK_PP(16'hCC28,4);
TASK_PP(16'hCC29,4);
TASK_PP(16'hCC2A,4);
TASK_PP(16'hCC2B,4);
TASK_PP(16'hCC2C,4);
TASK_PP(16'hCC2D,4);
TASK_PP(16'hCC2E,4);
TASK_PP(16'hCC2F,4);
TASK_PP(16'hCC30,4);
TASK_PP(16'hCC31,4);
TASK_PP(16'hCC32,4);
TASK_PP(16'hCC33,4);
TASK_PP(16'hCC34,4);
TASK_PP(16'hCC35,4);
TASK_PP(16'hCC36,4);
TASK_PP(16'hCC37,4);
TASK_PP(16'hCC38,4);
TASK_PP(16'hCC39,4);
TASK_PP(16'hCC3A,4);
TASK_PP(16'hCC3B,4);
TASK_PP(16'hCC3C,4);
TASK_PP(16'hCC3D,4);
TASK_PP(16'hCC3E,4);
TASK_PP(16'hCC3F,4);
TASK_PP(16'hCC40,4);
TASK_PP(16'hCC41,4);
TASK_PP(16'hCC42,4);
TASK_PP(16'hCC43,4);
TASK_PP(16'hCC44,4);
TASK_PP(16'hCC45,4);
TASK_PP(16'hCC46,4);
TASK_PP(16'hCC47,4);
TASK_PP(16'hCC48,4);
TASK_PP(16'hCC49,4);
TASK_PP(16'hCC4A,4);
TASK_PP(16'hCC4B,4);
TASK_PP(16'hCC4C,4);
TASK_PP(16'hCC4D,4);
TASK_PP(16'hCC4E,4);
TASK_PP(16'hCC4F,4);
TASK_PP(16'hCC50,4);
TASK_PP(16'hCC51,4);
TASK_PP(16'hCC52,4);
TASK_PP(16'hCC53,4);
TASK_PP(16'hCC54,4);
TASK_PP(16'hCC55,4);
TASK_PP(16'hCC56,4);
TASK_PP(16'hCC57,4);
TASK_PP(16'hCC58,4);
TASK_PP(16'hCC59,4);
TASK_PP(16'hCC5A,4);
TASK_PP(16'hCC5B,4);
TASK_PP(16'hCC5C,4);
TASK_PP(16'hCC5D,4);
TASK_PP(16'hCC5E,4);
TASK_PP(16'hCC5F,4);
TASK_PP(16'hCC60,4);
TASK_PP(16'hCC61,4);
TASK_PP(16'hCC62,4);
TASK_PP(16'hCC63,4);
TASK_PP(16'hCC64,4);
TASK_PP(16'hCC65,4);
TASK_PP(16'hCC66,4);
TASK_PP(16'hCC67,4);
TASK_PP(16'hCC68,4);
TASK_PP(16'hCC69,4);
TASK_PP(16'hCC6A,4);
TASK_PP(16'hCC6B,4);
TASK_PP(16'hCC6C,4);
TASK_PP(16'hCC6D,4);
TASK_PP(16'hCC6E,4);
TASK_PP(16'hCC6F,4);
TASK_PP(16'hCC70,4);
TASK_PP(16'hCC71,4);
TASK_PP(16'hCC72,4);
TASK_PP(16'hCC73,4);
TASK_PP(16'hCC74,4);
TASK_PP(16'hCC75,4);
TASK_PP(16'hCC76,4);
TASK_PP(16'hCC77,4);
TASK_PP(16'hCC78,4);
TASK_PP(16'hCC79,4);
TASK_PP(16'hCC7A,4);
TASK_PP(16'hCC7B,4);
TASK_PP(16'hCC7C,4);
TASK_PP(16'hCC7D,4);
TASK_PP(16'hCC7E,4);
TASK_PP(16'hCC7F,4);
TASK_PP(16'hCC80,4);
TASK_PP(16'hCC81,4);
TASK_PP(16'hCC82,4);
TASK_PP(16'hCC83,4);
TASK_PP(16'hCC84,4);
TASK_PP(16'hCC85,4);
TASK_PP(16'hCC86,4);
TASK_PP(16'hCC87,4);
TASK_PP(16'hCC88,4);
TASK_PP(16'hCC89,4);
TASK_PP(16'hCC8A,4);
TASK_PP(16'hCC8B,4);
TASK_PP(16'hCC8C,4);
TASK_PP(16'hCC8D,4);
TASK_PP(16'hCC8E,4);
TASK_PP(16'hCC8F,4);
TASK_PP(16'hCC90,4);
TASK_PP(16'hCC91,4);
TASK_PP(16'hCC92,4);
TASK_PP(16'hCC93,4);
TASK_PP(16'hCC94,4);
TASK_PP(16'hCC95,4);
TASK_PP(16'hCC96,4);
TASK_PP(16'hCC97,4);
TASK_PP(16'hCC98,4);
TASK_PP(16'hCC99,4);
TASK_PP(16'hCC9A,4);
TASK_PP(16'hCC9B,4);
TASK_PP(16'hCC9C,4);
TASK_PP(16'hCC9D,4);
TASK_PP(16'hCC9E,4);
TASK_PP(16'hCC9F,4);
TASK_PP(16'hCCA0,4);
TASK_PP(16'hCCA1,4);
TASK_PP(16'hCCA2,4);
TASK_PP(16'hCCA3,4);
TASK_PP(16'hCCA4,4);
TASK_PP(16'hCCA5,4);
TASK_PP(16'hCCA6,4);
TASK_PP(16'hCCA7,4);
TASK_PP(16'hCCA8,4);
TASK_PP(16'hCCA9,4);
TASK_PP(16'hCCAA,4);
TASK_PP(16'hCCAB,4);
TASK_PP(16'hCCAC,4);
TASK_PP(16'hCCAD,4);
TASK_PP(16'hCCAE,4);
TASK_PP(16'hCCAF,4);
TASK_PP(16'hCCB0,4);
TASK_PP(16'hCCB1,4);
TASK_PP(16'hCCB2,4);
TASK_PP(16'hCCB3,4);
TASK_PP(16'hCCB4,4);
TASK_PP(16'hCCB5,4);
TASK_PP(16'hCCB6,4);
TASK_PP(16'hCCB7,4);
TASK_PP(16'hCCB8,4);
TASK_PP(16'hCCB9,4);
TASK_PP(16'hCCBA,4);
TASK_PP(16'hCCBB,4);
TASK_PP(16'hCCBC,4);
TASK_PP(16'hCCBD,4);
TASK_PP(16'hCCBE,4);
TASK_PP(16'hCCBF,4);
TASK_PP(16'hCCC0,4);
TASK_PP(16'hCCC1,4);
TASK_PP(16'hCCC2,4);
TASK_PP(16'hCCC3,4);
TASK_PP(16'hCCC4,4);
TASK_PP(16'hCCC5,4);
TASK_PP(16'hCCC6,4);
TASK_PP(16'hCCC7,4);
TASK_PP(16'hCCC8,4);
TASK_PP(16'hCCC9,4);
TASK_PP(16'hCCCA,4);
TASK_PP(16'hCCCB,4);
TASK_PP(16'hCCCC,4);
TASK_PP(16'hCCCD,4);
TASK_PP(16'hCCCE,4);
TASK_PP(16'hCCCF,4);
TASK_PP(16'hCCD0,4);
TASK_PP(16'hCCD1,4);
TASK_PP(16'hCCD2,4);
TASK_PP(16'hCCD3,4);
TASK_PP(16'hCCD4,4);
TASK_PP(16'hCCD5,4);
TASK_PP(16'hCCD6,4);
TASK_PP(16'hCCD7,4);
TASK_PP(16'hCCD8,4);
TASK_PP(16'hCCD9,4);
TASK_PP(16'hCCDA,4);
TASK_PP(16'hCCDB,4);
TASK_PP(16'hCCDC,4);
TASK_PP(16'hCCDD,4);
TASK_PP(16'hCCDE,4);
TASK_PP(16'hCCDF,4);
TASK_PP(16'hCCE0,4);
TASK_PP(16'hCCE1,4);
TASK_PP(16'hCCE2,4);
TASK_PP(16'hCCE3,4);
TASK_PP(16'hCCE4,4);
TASK_PP(16'hCCE5,4);
TASK_PP(16'hCCE6,4);
TASK_PP(16'hCCE7,4);
TASK_PP(16'hCCE8,4);
TASK_PP(16'hCCE9,4);
TASK_PP(16'hCCEA,4);
TASK_PP(16'hCCEB,4);
TASK_PP(16'hCCEC,4);
TASK_PP(16'hCCED,4);
TASK_PP(16'hCCEE,4);
TASK_PP(16'hCCEF,4);
TASK_PP(16'hCCF0,4);
TASK_PP(16'hCCF1,4);
TASK_PP(16'hCCF2,4);
TASK_PP(16'hCCF3,4);
TASK_PP(16'hCCF4,4);
TASK_PP(16'hCCF5,4);
TASK_PP(16'hCCF6,4);
TASK_PP(16'hCCF7,4);
TASK_PP(16'hCCF8,4);
TASK_PP(16'hCCF9,4);
TASK_PP(16'hCCFA,4);
TASK_PP(16'hCCFB,4);
TASK_PP(16'hCCFC,4);
TASK_PP(16'hCCFD,4);
TASK_PP(16'hCCFE,4);
TASK_PP(16'hCCFF,4);
TASK_PP(16'hCD00,4);
TASK_PP(16'hCD01,4);
TASK_PP(16'hCD02,4);
TASK_PP(16'hCD03,4);
TASK_PP(16'hCD04,4);
TASK_PP(16'hCD05,4);
TASK_PP(16'hCD06,4);
TASK_PP(16'hCD07,4);
TASK_PP(16'hCD08,4);
TASK_PP(16'hCD09,4);
TASK_PP(16'hCD0A,4);
TASK_PP(16'hCD0B,4);
TASK_PP(16'hCD0C,4);
TASK_PP(16'hCD0D,4);
TASK_PP(16'hCD0E,4);
TASK_PP(16'hCD0F,4);
TASK_PP(16'hCD10,4);
TASK_PP(16'hCD11,4);
TASK_PP(16'hCD12,4);
TASK_PP(16'hCD13,4);
TASK_PP(16'hCD14,4);
TASK_PP(16'hCD15,4);
TASK_PP(16'hCD16,4);
TASK_PP(16'hCD17,4);
TASK_PP(16'hCD18,4);
TASK_PP(16'hCD19,4);
TASK_PP(16'hCD1A,4);
TASK_PP(16'hCD1B,4);
TASK_PP(16'hCD1C,4);
TASK_PP(16'hCD1D,4);
TASK_PP(16'hCD1E,4);
TASK_PP(16'hCD1F,4);
TASK_PP(16'hCD20,4);
TASK_PP(16'hCD21,4);
TASK_PP(16'hCD22,4);
TASK_PP(16'hCD23,4);
TASK_PP(16'hCD24,4);
TASK_PP(16'hCD25,4);
TASK_PP(16'hCD26,4);
TASK_PP(16'hCD27,4);
TASK_PP(16'hCD28,4);
TASK_PP(16'hCD29,4);
TASK_PP(16'hCD2A,4);
TASK_PP(16'hCD2B,4);
TASK_PP(16'hCD2C,4);
TASK_PP(16'hCD2D,4);
TASK_PP(16'hCD2E,4);
TASK_PP(16'hCD2F,4);
TASK_PP(16'hCD30,4);
TASK_PP(16'hCD31,4);
TASK_PP(16'hCD32,4);
TASK_PP(16'hCD33,4);
TASK_PP(16'hCD34,4);
TASK_PP(16'hCD35,4);
TASK_PP(16'hCD36,4);
TASK_PP(16'hCD37,4);
TASK_PP(16'hCD38,4);
TASK_PP(16'hCD39,4);
TASK_PP(16'hCD3A,4);
TASK_PP(16'hCD3B,4);
TASK_PP(16'hCD3C,4);
TASK_PP(16'hCD3D,4);
TASK_PP(16'hCD3E,4);
TASK_PP(16'hCD3F,4);
TASK_PP(16'hCD40,4);
TASK_PP(16'hCD41,4);
TASK_PP(16'hCD42,4);
TASK_PP(16'hCD43,4);
TASK_PP(16'hCD44,4);
TASK_PP(16'hCD45,4);
TASK_PP(16'hCD46,4);
TASK_PP(16'hCD47,4);
TASK_PP(16'hCD48,4);
TASK_PP(16'hCD49,4);
TASK_PP(16'hCD4A,4);
TASK_PP(16'hCD4B,4);
TASK_PP(16'hCD4C,4);
TASK_PP(16'hCD4D,4);
TASK_PP(16'hCD4E,4);
TASK_PP(16'hCD4F,4);
TASK_PP(16'hCD50,4);
TASK_PP(16'hCD51,4);
TASK_PP(16'hCD52,4);
TASK_PP(16'hCD53,4);
TASK_PP(16'hCD54,4);
TASK_PP(16'hCD55,4);
TASK_PP(16'hCD56,4);
TASK_PP(16'hCD57,4);
TASK_PP(16'hCD58,4);
TASK_PP(16'hCD59,4);
TASK_PP(16'hCD5A,4);
TASK_PP(16'hCD5B,4);
TASK_PP(16'hCD5C,4);
TASK_PP(16'hCD5D,4);
TASK_PP(16'hCD5E,4);
TASK_PP(16'hCD5F,4);
TASK_PP(16'hCD60,4);
TASK_PP(16'hCD61,4);
TASK_PP(16'hCD62,4);
TASK_PP(16'hCD63,4);
TASK_PP(16'hCD64,4);
TASK_PP(16'hCD65,4);
TASK_PP(16'hCD66,4);
TASK_PP(16'hCD67,4);
TASK_PP(16'hCD68,4);
TASK_PP(16'hCD69,4);
TASK_PP(16'hCD6A,4);
TASK_PP(16'hCD6B,4);
TASK_PP(16'hCD6C,4);
TASK_PP(16'hCD6D,4);
TASK_PP(16'hCD6E,4);
TASK_PP(16'hCD6F,4);
TASK_PP(16'hCD70,4);
TASK_PP(16'hCD71,4);
TASK_PP(16'hCD72,4);
TASK_PP(16'hCD73,4);
TASK_PP(16'hCD74,4);
TASK_PP(16'hCD75,4);
TASK_PP(16'hCD76,4);
TASK_PP(16'hCD77,4);
TASK_PP(16'hCD78,4);
TASK_PP(16'hCD79,4);
TASK_PP(16'hCD7A,4);
TASK_PP(16'hCD7B,4);
TASK_PP(16'hCD7C,4);
TASK_PP(16'hCD7D,4);
TASK_PP(16'hCD7E,4);
TASK_PP(16'hCD7F,4);
TASK_PP(16'hCD80,4);
TASK_PP(16'hCD81,4);
TASK_PP(16'hCD82,4);
TASK_PP(16'hCD83,4);
TASK_PP(16'hCD84,4);
TASK_PP(16'hCD85,4);
TASK_PP(16'hCD86,4);
TASK_PP(16'hCD87,4);
TASK_PP(16'hCD88,4);
TASK_PP(16'hCD89,4);
TASK_PP(16'hCD8A,4);
TASK_PP(16'hCD8B,4);
TASK_PP(16'hCD8C,4);
TASK_PP(16'hCD8D,4);
TASK_PP(16'hCD8E,4);
TASK_PP(16'hCD8F,4);
TASK_PP(16'hCD90,4);
TASK_PP(16'hCD91,4);
TASK_PP(16'hCD92,4);
TASK_PP(16'hCD93,4);
TASK_PP(16'hCD94,4);
TASK_PP(16'hCD95,4);
TASK_PP(16'hCD96,4);
TASK_PP(16'hCD97,4);
TASK_PP(16'hCD98,4);
TASK_PP(16'hCD99,4);
TASK_PP(16'hCD9A,4);
TASK_PP(16'hCD9B,4);
TASK_PP(16'hCD9C,4);
TASK_PP(16'hCD9D,4);
TASK_PP(16'hCD9E,4);
TASK_PP(16'hCD9F,4);
TASK_PP(16'hCDA0,4);
TASK_PP(16'hCDA1,4);
TASK_PP(16'hCDA2,4);
TASK_PP(16'hCDA3,4);
TASK_PP(16'hCDA4,4);
TASK_PP(16'hCDA5,4);
TASK_PP(16'hCDA6,4);
TASK_PP(16'hCDA7,4);
TASK_PP(16'hCDA8,4);
TASK_PP(16'hCDA9,4);
TASK_PP(16'hCDAA,4);
TASK_PP(16'hCDAB,4);
TASK_PP(16'hCDAC,4);
TASK_PP(16'hCDAD,4);
TASK_PP(16'hCDAE,4);
TASK_PP(16'hCDAF,4);
TASK_PP(16'hCDB0,4);
TASK_PP(16'hCDB1,4);
TASK_PP(16'hCDB2,4);
TASK_PP(16'hCDB3,4);
TASK_PP(16'hCDB4,4);
TASK_PP(16'hCDB5,4);
TASK_PP(16'hCDB6,4);
TASK_PP(16'hCDB7,4);
TASK_PP(16'hCDB8,4);
TASK_PP(16'hCDB9,4);
TASK_PP(16'hCDBA,4);
TASK_PP(16'hCDBB,4);
TASK_PP(16'hCDBC,4);
TASK_PP(16'hCDBD,4);
TASK_PP(16'hCDBE,4);
TASK_PP(16'hCDBF,4);
TASK_PP(16'hCDC0,4);
TASK_PP(16'hCDC1,4);
TASK_PP(16'hCDC2,4);
TASK_PP(16'hCDC3,4);
TASK_PP(16'hCDC4,4);
TASK_PP(16'hCDC5,4);
TASK_PP(16'hCDC6,4);
TASK_PP(16'hCDC7,4);
TASK_PP(16'hCDC8,4);
TASK_PP(16'hCDC9,4);
TASK_PP(16'hCDCA,4);
TASK_PP(16'hCDCB,4);
TASK_PP(16'hCDCC,4);
TASK_PP(16'hCDCD,4);
TASK_PP(16'hCDCE,4);
TASK_PP(16'hCDCF,4);
TASK_PP(16'hCDD0,4);
TASK_PP(16'hCDD1,4);
TASK_PP(16'hCDD2,4);
TASK_PP(16'hCDD3,4);
TASK_PP(16'hCDD4,4);
TASK_PP(16'hCDD5,4);
TASK_PP(16'hCDD6,4);
TASK_PP(16'hCDD7,4);
TASK_PP(16'hCDD8,4);
TASK_PP(16'hCDD9,4);
TASK_PP(16'hCDDA,4);
TASK_PP(16'hCDDB,4);
TASK_PP(16'hCDDC,4);
TASK_PP(16'hCDDD,4);
TASK_PP(16'hCDDE,4);
TASK_PP(16'hCDDF,4);
TASK_PP(16'hCDE0,4);
TASK_PP(16'hCDE1,4);
TASK_PP(16'hCDE2,4);
TASK_PP(16'hCDE3,4);
TASK_PP(16'hCDE4,4);
TASK_PP(16'hCDE5,4);
TASK_PP(16'hCDE6,4);
TASK_PP(16'hCDE7,4);
TASK_PP(16'hCDE8,4);
TASK_PP(16'hCDE9,4);
TASK_PP(16'hCDEA,4);
TASK_PP(16'hCDEB,4);
TASK_PP(16'hCDEC,4);
TASK_PP(16'hCDED,4);
TASK_PP(16'hCDEE,4);
TASK_PP(16'hCDEF,4);
TASK_PP(16'hCDF0,4);
TASK_PP(16'hCDF1,4);
TASK_PP(16'hCDF2,4);
TASK_PP(16'hCDF3,4);
TASK_PP(16'hCDF4,4);
TASK_PP(16'hCDF5,4);
TASK_PP(16'hCDF6,4);
TASK_PP(16'hCDF7,4);
TASK_PP(16'hCDF8,4);
TASK_PP(16'hCDF9,4);
TASK_PP(16'hCDFA,4);
TASK_PP(16'hCDFB,4);
TASK_PP(16'hCDFC,4);
TASK_PP(16'hCDFD,4);
TASK_PP(16'hCDFE,4);
TASK_PP(16'hCDFF,4);
TASK_PP(16'hCE00,4);
TASK_PP(16'hCE01,4);
TASK_PP(16'hCE02,4);
TASK_PP(16'hCE03,4);
TASK_PP(16'hCE04,4);
TASK_PP(16'hCE05,4);
TASK_PP(16'hCE06,4);
TASK_PP(16'hCE07,4);
TASK_PP(16'hCE08,4);
TASK_PP(16'hCE09,4);
TASK_PP(16'hCE0A,4);
TASK_PP(16'hCE0B,4);
TASK_PP(16'hCE0C,4);
TASK_PP(16'hCE0D,4);
TASK_PP(16'hCE0E,4);
TASK_PP(16'hCE0F,4);
TASK_PP(16'hCE10,4);
TASK_PP(16'hCE11,4);
TASK_PP(16'hCE12,4);
TASK_PP(16'hCE13,4);
TASK_PP(16'hCE14,4);
TASK_PP(16'hCE15,4);
TASK_PP(16'hCE16,4);
TASK_PP(16'hCE17,4);
TASK_PP(16'hCE18,4);
TASK_PP(16'hCE19,4);
TASK_PP(16'hCE1A,4);
TASK_PP(16'hCE1B,4);
TASK_PP(16'hCE1C,4);
TASK_PP(16'hCE1D,4);
TASK_PP(16'hCE1E,4);
TASK_PP(16'hCE1F,4);
TASK_PP(16'hCE20,4);
TASK_PP(16'hCE21,4);
TASK_PP(16'hCE22,4);
TASK_PP(16'hCE23,4);
TASK_PP(16'hCE24,4);
TASK_PP(16'hCE25,4);
TASK_PP(16'hCE26,4);
TASK_PP(16'hCE27,4);
TASK_PP(16'hCE28,4);
TASK_PP(16'hCE29,4);
TASK_PP(16'hCE2A,4);
TASK_PP(16'hCE2B,4);
TASK_PP(16'hCE2C,4);
TASK_PP(16'hCE2D,4);
TASK_PP(16'hCE2E,4);
TASK_PP(16'hCE2F,4);
TASK_PP(16'hCE30,4);
TASK_PP(16'hCE31,4);
TASK_PP(16'hCE32,4);
TASK_PP(16'hCE33,4);
TASK_PP(16'hCE34,4);
TASK_PP(16'hCE35,4);
TASK_PP(16'hCE36,4);
TASK_PP(16'hCE37,4);
TASK_PP(16'hCE38,4);
TASK_PP(16'hCE39,4);
TASK_PP(16'hCE3A,4);
TASK_PP(16'hCE3B,4);
TASK_PP(16'hCE3C,4);
TASK_PP(16'hCE3D,4);
TASK_PP(16'hCE3E,4);
TASK_PP(16'hCE3F,4);
TASK_PP(16'hCE40,4);
TASK_PP(16'hCE41,4);
TASK_PP(16'hCE42,4);
TASK_PP(16'hCE43,4);
TASK_PP(16'hCE44,4);
TASK_PP(16'hCE45,4);
TASK_PP(16'hCE46,4);
TASK_PP(16'hCE47,4);
TASK_PP(16'hCE48,4);
TASK_PP(16'hCE49,4);
TASK_PP(16'hCE4A,4);
TASK_PP(16'hCE4B,4);
TASK_PP(16'hCE4C,4);
TASK_PP(16'hCE4D,4);
TASK_PP(16'hCE4E,4);
TASK_PP(16'hCE4F,4);
TASK_PP(16'hCE50,4);
TASK_PP(16'hCE51,4);
TASK_PP(16'hCE52,4);
TASK_PP(16'hCE53,4);
TASK_PP(16'hCE54,4);
TASK_PP(16'hCE55,4);
TASK_PP(16'hCE56,4);
TASK_PP(16'hCE57,4);
TASK_PP(16'hCE58,4);
TASK_PP(16'hCE59,4);
TASK_PP(16'hCE5A,4);
TASK_PP(16'hCE5B,4);
TASK_PP(16'hCE5C,4);
TASK_PP(16'hCE5D,4);
TASK_PP(16'hCE5E,4);
TASK_PP(16'hCE5F,4);
TASK_PP(16'hCE60,4);
TASK_PP(16'hCE61,4);
TASK_PP(16'hCE62,4);
TASK_PP(16'hCE63,4);
TASK_PP(16'hCE64,4);
TASK_PP(16'hCE65,4);
TASK_PP(16'hCE66,4);
TASK_PP(16'hCE67,4);
TASK_PP(16'hCE68,4);
TASK_PP(16'hCE69,4);
TASK_PP(16'hCE6A,4);
TASK_PP(16'hCE6B,4);
TASK_PP(16'hCE6C,4);
TASK_PP(16'hCE6D,4);
TASK_PP(16'hCE6E,4);
TASK_PP(16'hCE6F,4);
TASK_PP(16'hCE70,4);
TASK_PP(16'hCE71,4);
TASK_PP(16'hCE72,4);
TASK_PP(16'hCE73,4);
TASK_PP(16'hCE74,4);
TASK_PP(16'hCE75,4);
TASK_PP(16'hCE76,4);
TASK_PP(16'hCE77,4);
TASK_PP(16'hCE78,4);
TASK_PP(16'hCE79,4);
TASK_PP(16'hCE7A,4);
TASK_PP(16'hCE7B,4);
TASK_PP(16'hCE7C,4);
TASK_PP(16'hCE7D,4);
TASK_PP(16'hCE7E,4);
TASK_PP(16'hCE7F,4);
TASK_PP(16'hCE80,4);
TASK_PP(16'hCE81,4);
TASK_PP(16'hCE82,4);
TASK_PP(16'hCE83,4);
TASK_PP(16'hCE84,4);
TASK_PP(16'hCE85,4);
TASK_PP(16'hCE86,4);
TASK_PP(16'hCE87,4);
TASK_PP(16'hCE88,4);
TASK_PP(16'hCE89,4);
TASK_PP(16'hCE8A,4);
TASK_PP(16'hCE8B,4);
TASK_PP(16'hCE8C,4);
TASK_PP(16'hCE8D,4);
TASK_PP(16'hCE8E,4);
TASK_PP(16'hCE8F,4);
TASK_PP(16'hCE90,4);
TASK_PP(16'hCE91,4);
TASK_PP(16'hCE92,4);
TASK_PP(16'hCE93,4);
TASK_PP(16'hCE94,4);
TASK_PP(16'hCE95,4);
TASK_PP(16'hCE96,4);
TASK_PP(16'hCE97,4);
TASK_PP(16'hCE98,4);
TASK_PP(16'hCE99,4);
TASK_PP(16'hCE9A,4);
TASK_PP(16'hCE9B,4);
TASK_PP(16'hCE9C,4);
TASK_PP(16'hCE9D,4);
TASK_PP(16'hCE9E,4);
TASK_PP(16'hCE9F,4);
TASK_PP(16'hCEA0,4);
TASK_PP(16'hCEA1,4);
TASK_PP(16'hCEA2,4);
TASK_PP(16'hCEA3,4);
TASK_PP(16'hCEA4,4);
TASK_PP(16'hCEA5,4);
TASK_PP(16'hCEA6,4);
TASK_PP(16'hCEA7,4);
TASK_PP(16'hCEA8,4);
TASK_PP(16'hCEA9,4);
TASK_PP(16'hCEAA,4);
TASK_PP(16'hCEAB,4);
TASK_PP(16'hCEAC,4);
TASK_PP(16'hCEAD,4);
TASK_PP(16'hCEAE,4);
TASK_PP(16'hCEAF,4);
TASK_PP(16'hCEB0,4);
TASK_PP(16'hCEB1,4);
TASK_PP(16'hCEB2,4);
TASK_PP(16'hCEB3,4);
TASK_PP(16'hCEB4,4);
TASK_PP(16'hCEB5,4);
TASK_PP(16'hCEB6,4);
TASK_PP(16'hCEB7,4);
TASK_PP(16'hCEB8,4);
TASK_PP(16'hCEB9,4);
TASK_PP(16'hCEBA,4);
TASK_PP(16'hCEBB,4);
TASK_PP(16'hCEBC,4);
TASK_PP(16'hCEBD,4);
TASK_PP(16'hCEBE,4);
TASK_PP(16'hCEBF,4);
TASK_PP(16'hCEC0,4);
TASK_PP(16'hCEC1,4);
TASK_PP(16'hCEC2,4);
TASK_PP(16'hCEC3,4);
TASK_PP(16'hCEC4,4);
TASK_PP(16'hCEC5,4);
TASK_PP(16'hCEC6,4);
TASK_PP(16'hCEC7,4);
TASK_PP(16'hCEC8,4);
TASK_PP(16'hCEC9,4);
TASK_PP(16'hCECA,4);
TASK_PP(16'hCECB,4);
TASK_PP(16'hCECC,4);
TASK_PP(16'hCECD,4);
TASK_PP(16'hCECE,4);
TASK_PP(16'hCECF,4);
TASK_PP(16'hCED0,4);
TASK_PP(16'hCED1,4);
TASK_PP(16'hCED2,4);
TASK_PP(16'hCED3,4);
TASK_PP(16'hCED4,4);
TASK_PP(16'hCED5,4);
TASK_PP(16'hCED6,4);
TASK_PP(16'hCED7,4);
TASK_PP(16'hCED8,4);
TASK_PP(16'hCED9,4);
TASK_PP(16'hCEDA,4);
TASK_PP(16'hCEDB,4);
TASK_PP(16'hCEDC,4);
TASK_PP(16'hCEDD,4);
TASK_PP(16'hCEDE,4);
TASK_PP(16'hCEDF,4);
TASK_PP(16'hCEE0,4);
TASK_PP(16'hCEE1,4);
TASK_PP(16'hCEE2,4);
TASK_PP(16'hCEE3,4);
TASK_PP(16'hCEE4,4);
TASK_PP(16'hCEE5,4);
TASK_PP(16'hCEE6,4);
TASK_PP(16'hCEE7,4);
TASK_PP(16'hCEE8,4);
TASK_PP(16'hCEE9,4);
TASK_PP(16'hCEEA,4);
TASK_PP(16'hCEEB,4);
TASK_PP(16'hCEEC,4);
TASK_PP(16'hCEED,4);
TASK_PP(16'hCEEE,4);
TASK_PP(16'hCEEF,4);
TASK_PP(16'hCEF0,4);
TASK_PP(16'hCEF1,4);
TASK_PP(16'hCEF2,4);
TASK_PP(16'hCEF3,4);
TASK_PP(16'hCEF4,4);
TASK_PP(16'hCEF5,4);
TASK_PP(16'hCEF6,4);
TASK_PP(16'hCEF7,4);
TASK_PP(16'hCEF8,4);
TASK_PP(16'hCEF9,4);
TASK_PP(16'hCEFA,4);
TASK_PP(16'hCEFB,4);
TASK_PP(16'hCEFC,4);
TASK_PP(16'hCEFD,4);
TASK_PP(16'hCEFE,4);
TASK_PP(16'hCEFF,4);
TASK_PP(16'hCF00,4);
TASK_PP(16'hCF01,4);
TASK_PP(16'hCF02,4);
TASK_PP(16'hCF03,4);
TASK_PP(16'hCF04,4);
TASK_PP(16'hCF05,4);
TASK_PP(16'hCF06,4);
TASK_PP(16'hCF07,4);
TASK_PP(16'hCF08,4);
TASK_PP(16'hCF09,4);
TASK_PP(16'hCF0A,4);
TASK_PP(16'hCF0B,4);
TASK_PP(16'hCF0C,4);
TASK_PP(16'hCF0D,4);
TASK_PP(16'hCF0E,4);
TASK_PP(16'hCF0F,4);
TASK_PP(16'hCF10,4);
TASK_PP(16'hCF11,4);
TASK_PP(16'hCF12,4);
TASK_PP(16'hCF13,4);
TASK_PP(16'hCF14,4);
TASK_PP(16'hCF15,4);
TASK_PP(16'hCF16,4);
TASK_PP(16'hCF17,4);
TASK_PP(16'hCF18,4);
TASK_PP(16'hCF19,4);
TASK_PP(16'hCF1A,4);
TASK_PP(16'hCF1B,4);
TASK_PP(16'hCF1C,4);
TASK_PP(16'hCF1D,4);
TASK_PP(16'hCF1E,4);
TASK_PP(16'hCF1F,4);
TASK_PP(16'hCF20,4);
TASK_PP(16'hCF21,4);
TASK_PP(16'hCF22,4);
TASK_PP(16'hCF23,4);
TASK_PP(16'hCF24,4);
TASK_PP(16'hCF25,4);
TASK_PP(16'hCF26,4);
TASK_PP(16'hCF27,4);
TASK_PP(16'hCF28,4);
TASK_PP(16'hCF29,4);
TASK_PP(16'hCF2A,4);
TASK_PP(16'hCF2B,4);
TASK_PP(16'hCF2C,4);
TASK_PP(16'hCF2D,4);
TASK_PP(16'hCF2E,4);
TASK_PP(16'hCF2F,4);
TASK_PP(16'hCF30,4);
TASK_PP(16'hCF31,4);
TASK_PP(16'hCF32,4);
TASK_PP(16'hCF33,4);
TASK_PP(16'hCF34,4);
TASK_PP(16'hCF35,4);
TASK_PP(16'hCF36,4);
TASK_PP(16'hCF37,4);
TASK_PP(16'hCF38,4);
TASK_PP(16'hCF39,4);
TASK_PP(16'hCF3A,4);
TASK_PP(16'hCF3B,4);
TASK_PP(16'hCF3C,4);
TASK_PP(16'hCF3D,4);
TASK_PP(16'hCF3E,4);
TASK_PP(16'hCF3F,4);
TASK_PP(16'hCF40,4);
TASK_PP(16'hCF41,4);
TASK_PP(16'hCF42,4);
TASK_PP(16'hCF43,4);
TASK_PP(16'hCF44,4);
TASK_PP(16'hCF45,4);
TASK_PP(16'hCF46,4);
TASK_PP(16'hCF47,4);
TASK_PP(16'hCF48,4);
TASK_PP(16'hCF49,4);
TASK_PP(16'hCF4A,4);
TASK_PP(16'hCF4B,4);
TASK_PP(16'hCF4C,4);
TASK_PP(16'hCF4D,4);
TASK_PP(16'hCF4E,4);
TASK_PP(16'hCF4F,4);
TASK_PP(16'hCF50,4);
TASK_PP(16'hCF51,4);
TASK_PP(16'hCF52,4);
TASK_PP(16'hCF53,4);
TASK_PP(16'hCF54,4);
TASK_PP(16'hCF55,4);
TASK_PP(16'hCF56,4);
TASK_PP(16'hCF57,4);
TASK_PP(16'hCF58,4);
TASK_PP(16'hCF59,4);
TASK_PP(16'hCF5A,4);
TASK_PP(16'hCF5B,4);
TASK_PP(16'hCF5C,4);
TASK_PP(16'hCF5D,4);
TASK_PP(16'hCF5E,4);
TASK_PP(16'hCF5F,4);
TASK_PP(16'hCF60,4);
TASK_PP(16'hCF61,4);
TASK_PP(16'hCF62,4);
TASK_PP(16'hCF63,4);
TASK_PP(16'hCF64,4);
TASK_PP(16'hCF65,4);
TASK_PP(16'hCF66,4);
TASK_PP(16'hCF67,4);
TASK_PP(16'hCF68,4);
TASK_PP(16'hCF69,4);
TASK_PP(16'hCF6A,4);
TASK_PP(16'hCF6B,4);
TASK_PP(16'hCF6C,4);
TASK_PP(16'hCF6D,4);
TASK_PP(16'hCF6E,4);
TASK_PP(16'hCF6F,4);
TASK_PP(16'hCF70,4);
TASK_PP(16'hCF71,4);
TASK_PP(16'hCF72,4);
TASK_PP(16'hCF73,4);
TASK_PP(16'hCF74,4);
TASK_PP(16'hCF75,4);
TASK_PP(16'hCF76,4);
TASK_PP(16'hCF77,4);
TASK_PP(16'hCF78,4);
TASK_PP(16'hCF79,4);
TASK_PP(16'hCF7A,4);
TASK_PP(16'hCF7B,4);
TASK_PP(16'hCF7C,4);
TASK_PP(16'hCF7D,4);
TASK_PP(16'hCF7E,4);
TASK_PP(16'hCF7F,4);
TASK_PP(16'hCF80,4);
TASK_PP(16'hCF81,4);
TASK_PP(16'hCF82,4);
TASK_PP(16'hCF83,4);
TASK_PP(16'hCF84,4);
TASK_PP(16'hCF85,4);
TASK_PP(16'hCF86,4);
TASK_PP(16'hCF87,4);
TASK_PP(16'hCF88,4);
TASK_PP(16'hCF89,4);
TASK_PP(16'hCF8A,4);
TASK_PP(16'hCF8B,4);
TASK_PP(16'hCF8C,4);
TASK_PP(16'hCF8D,4);
TASK_PP(16'hCF8E,4);
TASK_PP(16'hCF8F,4);
TASK_PP(16'hCF90,4);
TASK_PP(16'hCF91,4);
TASK_PP(16'hCF92,4);
TASK_PP(16'hCF93,4);
TASK_PP(16'hCF94,4);
TASK_PP(16'hCF95,4);
TASK_PP(16'hCF96,4);
TASK_PP(16'hCF97,4);
TASK_PP(16'hCF98,4);
TASK_PP(16'hCF99,4);
TASK_PP(16'hCF9A,4);
TASK_PP(16'hCF9B,4);
TASK_PP(16'hCF9C,4);
TASK_PP(16'hCF9D,4);
TASK_PP(16'hCF9E,4);
TASK_PP(16'hCF9F,4);
TASK_PP(16'hCFA0,4);
TASK_PP(16'hCFA1,4);
TASK_PP(16'hCFA2,4);
TASK_PP(16'hCFA3,4);
TASK_PP(16'hCFA4,4);
TASK_PP(16'hCFA5,4);
TASK_PP(16'hCFA6,4);
TASK_PP(16'hCFA7,4);
TASK_PP(16'hCFA8,4);
TASK_PP(16'hCFA9,4);
TASK_PP(16'hCFAA,4);
TASK_PP(16'hCFAB,4);
TASK_PP(16'hCFAC,4);
TASK_PP(16'hCFAD,4);
TASK_PP(16'hCFAE,4);
TASK_PP(16'hCFAF,4);
TASK_PP(16'hCFB0,4);
TASK_PP(16'hCFB1,4);
TASK_PP(16'hCFB2,4);
TASK_PP(16'hCFB3,4);
TASK_PP(16'hCFB4,4);
TASK_PP(16'hCFB5,4);
TASK_PP(16'hCFB6,4);
TASK_PP(16'hCFB7,4);
TASK_PP(16'hCFB8,4);
TASK_PP(16'hCFB9,4);
TASK_PP(16'hCFBA,4);
TASK_PP(16'hCFBB,4);
TASK_PP(16'hCFBC,4);
TASK_PP(16'hCFBD,4);
TASK_PP(16'hCFBE,4);
TASK_PP(16'hCFBF,4);
TASK_PP(16'hCFC0,4);
TASK_PP(16'hCFC1,4);
TASK_PP(16'hCFC2,4);
TASK_PP(16'hCFC3,4);
TASK_PP(16'hCFC4,4);
TASK_PP(16'hCFC5,4);
TASK_PP(16'hCFC6,4);
TASK_PP(16'hCFC7,4);
TASK_PP(16'hCFC8,4);
TASK_PP(16'hCFC9,4);
TASK_PP(16'hCFCA,4);
TASK_PP(16'hCFCB,4);
TASK_PP(16'hCFCC,4);
TASK_PP(16'hCFCD,4);
TASK_PP(16'hCFCE,4);
TASK_PP(16'hCFCF,4);
TASK_PP(16'hCFD0,4);
TASK_PP(16'hCFD1,4);
TASK_PP(16'hCFD2,4);
TASK_PP(16'hCFD3,4);
TASK_PP(16'hCFD4,4);
TASK_PP(16'hCFD5,4);
TASK_PP(16'hCFD6,4);
TASK_PP(16'hCFD7,4);
TASK_PP(16'hCFD8,4);
TASK_PP(16'hCFD9,4);
TASK_PP(16'hCFDA,4);
TASK_PP(16'hCFDB,4);
TASK_PP(16'hCFDC,4);
TASK_PP(16'hCFDD,4);
TASK_PP(16'hCFDE,4);
TASK_PP(16'hCFDF,4);
TASK_PP(16'hCFE0,4);
TASK_PP(16'hCFE1,4);
TASK_PP(16'hCFE2,4);
TASK_PP(16'hCFE3,4);
TASK_PP(16'hCFE4,4);
TASK_PP(16'hCFE5,4);
TASK_PP(16'hCFE6,4);
TASK_PP(16'hCFE7,4);
TASK_PP(16'hCFE8,4);
TASK_PP(16'hCFE9,4);
TASK_PP(16'hCFEA,4);
TASK_PP(16'hCFEB,4);
TASK_PP(16'hCFEC,4);
TASK_PP(16'hCFED,4);
TASK_PP(16'hCFEE,4);
TASK_PP(16'hCFEF,4);
TASK_PP(16'hCFF0,4);
TASK_PP(16'hCFF1,4);
TASK_PP(16'hCFF2,4);
TASK_PP(16'hCFF3,4);
TASK_PP(16'hCFF4,4);
TASK_PP(16'hCFF5,4);
TASK_PP(16'hCFF6,4);
TASK_PP(16'hCFF7,4);
TASK_PP(16'hCFF8,4);
TASK_PP(16'hCFF9,4);
TASK_PP(16'hCFFA,4);
TASK_PP(16'hCFFB,4);
TASK_PP(16'hCFFC,4);
TASK_PP(16'hCFFD,4);
TASK_PP(16'hCFFE,4);
TASK_PP(16'hCFFF,4);
TASK_PP(16'hD000,4);
TASK_PP(16'hD001,4);
TASK_PP(16'hD002,4);
TASK_PP(16'hD003,4);
TASK_PP(16'hD004,4);
TASK_PP(16'hD005,4);
TASK_PP(16'hD006,4);
TASK_PP(16'hD007,4);
TASK_PP(16'hD008,4);
TASK_PP(16'hD009,4);
TASK_PP(16'hD00A,4);
TASK_PP(16'hD00B,4);
TASK_PP(16'hD00C,4);
TASK_PP(16'hD00D,4);
TASK_PP(16'hD00E,4);
TASK_PP(16'hD00F,4);
TASK_PP(16'hD010,4);
TASK_PP(16'hD011,4);
TASK_PP(16'hD012,4);
TASK_PP(16'hD013,4);
TASK_PP(16'hD014,4);
TASK_PP(16'hD015,4);
TASK_PP(16'hD016,4);
TASK_PP(16'hD017,4);
TASK_PP(16'hD018,4);
TASK_PP(16'hD019,4);
TASK_PP(16'hD01A,4);
TASK_PP(16'hD01B,4);
TASK_PP(16'hD01C,4);
TASK_PP(16'hD01D,4);
TASK_PP(16'hD01E,4);
TASK_PP(16'hD01F,4);
TASK_PP(16'hD020,4);
TASK_PP(16'hD021,4);
TASK_PP(16'hD022,4);
TASK_PP(16'hD023,4);
TASK_PP(16'hD024,4);
TASK_PP(16'hD025,4);
TASK_PP(16'hD026,4);
TASK_PP(16'hD027,4);
TASK_PP(16'hD028,4);
TASK_PP(16'hD029,4);
TASK_PP(16'hD02A,4);
TASK_PP(16'hD02B,4);
TASK_PP(16'hD02C,4);
TASK_PP(16'hD02D,4);
TASK_PP(16'hD02E,4);
TASK_PP(16'hD02F,4);
TASK_PP(16'hD030,4);
TASK_PP(16'hD031,4);
TASK_PP(16'hD032,4);
TASK_PP(16'hD033,4);
TASK_PP(16'hD034,4);
TASK_PP(16'hD035,4);
TASK_PP(16'hD036,4);
TASK_PP(16'hD037,4);
TASK_PP(16'hD038,4);
TASK_PP(16'hD039,4);
TASK_PP(16'hD03A,4);
TASK_PP(16'hD03B,4);
TASK_PP(16'hD03C,4);
TASK_PP(16'hD03D,4);
TASK_PP(16'hD03E,4);
TASK_PP(16'hD03F,4);
TASK_PP(16'hD040,4);
TASK_PP(16'hD041,4);
TASK_PP(16'hD042,4);
TASK_PP(16'hD043,4);
TASK_PP(16'hD044,4);
TASK_PP(16'hD045,4);
TASK_PP(16'hD046,4);
TASK_PP(16'hD047,4);
TASK_PP(16'hD048,4);
TASK_PP(16'hD049,4);
TASK_PP(16'hD04A,4);
TASK_PP(16'hD04B,4);
TASK_PP(16'hD04C,4);
TASK_PP(16'hD04D,4);
TASK_PP(16'hD04E,4);
TASK_PP(16'hD04F,4);
TASK_PP(16'hD050,4);
TASK_PP(16'hD051,4);
TASK_PP(16'hD052,4);
TASK_PP(16'hD053,4);
TASK_PP(16'hD054,4);
TASK_PP(16'hD055,4);
TASK_PP(16'hD056,4);
TASK_PP(16'hD057,4);
TASK_PP(16'hD058,4);
TASK_PP(16'hD059,4);
TASK_PP(16'hD05A,4);
TASK_PP(16'hD05B,4);
TASK_PP(16'hD05C,4);
TASK_PP(16'hD05D,4);
TASK_PP(16'hD05E,4);
TASK_PP(16'hD05F,4);
TASK_PP(16'hD060,4);
TASK_PP(16'hD061,4);
TASK_PP(16'hD062,4);
TASK_PP(16'hD063,4);
TASK_PP(16'hD064,4);
TASK_PP(16'hD065,4);
TASK_PP(16'hD066,4);
TASK_PP(16'hD067,4);
TASK_PP(16'hD068,4);
TASK_PP(16'hD069,4);
TASK_PP(16'hD06A,4);
TASK_PP(16'hD06B,4);
TASK_PP(16'hD06C,4);
TASK_PP(16'hD06D,4);
TASK_PP(16'hD06E,4);
TASK_PP(16'hD06F,4);
TASK_PP(16'hD070,4);
TASK_PP(16'hD071,4);
TASK_PP(16'hD072,4);
TASK_PP(16'hD073,4);
TASK_PP(16'hD074,4);
TASK_PP(16'hD075,4);
TASK_PP(16'hD076,4);
TASK_PP(16'hD077,4);
TASK_PP(16'hD078,4);
TASK_PP(16'hD079,4);
TASK_PP(16'hD07A,4);
TASK_PP(16'hD07B,4);
TASK_PP(16'hD07C,4);
TASK_PP(16'hD07D,4);
TASK_PP(16'hD07E,4);
TASK_PP(16'hD07F,4);
TASK_PP(16'hD080,4);
TASK_PP(16'hD081,4);
TASK_PP(16'hD082,4);
TASK_PP(16'hD083,4);
TASK_PP(16'hD084,4);
TASK_PP(16'hD085,4);
TASK_PP(16'hD086,4);
TASK_PP(16'hD087,4);
TASK_PP(16'hD088,4);
TASK_PP(16'hD089,4);
TASK_PP(16'hD08A,4);
TASK_PP(16'hD08B,4);
TASK_PP(16'hD08C,4);
TASK_PP(16'hD08D,4);
TASK_PP(16'hD08E,4);
TASK_PP(16'hD08F,4);
TASK_PP(16'hD090,4);
TASK_PP(16'hD091,4);
TASK_PP(16'hD092,4);
TASK_PP(16'hD093,4);
TASK_PP(16'hD094,4);
TASK_PP(16'hD095,4);
TASK_PP(16'hD096,4);
TASK_PP(16'hD097,4);
TASK_PP(16'hD098,4);
TASK_PP(16'hD099,4);
TASK_PP(16'hD09A,4);
TASK_PP(16'hD09B,4);
TASK_PP(16'hD09C,4);
TASK_PP(16'hD09D,4);
TASK_PP(16'hD09E,4);
TASK_PP(16'hD09F,4);
TASK_PP(16'hD0A0,4);
TASK_PP(16'hD0A1,4);
TASK_PP(16'hD0A2,4);
TASK_PP(16'hD0A3,4);
TASK_PP(16'hD0A4,4);
TASK_PP(16'hD0A5,4);
TASK_PP(16'hD0A6,4);
TASK_PP(16'hD0A7,4);
TASK_PP(16'hD0A8,4);
TASK_PP(16'hD0A9,4);
TASK_PP(16'hD0AA,4);
TASK_PP(16'hD0AB,4);
TASK_PP(16'hD0AC,4);
TASK_PP(16'hD0AD,4);
TASK_PP(16'hD0AE,4);
TASK_PP(16'hD0AF,4);
TASK_PP(16'hD0B0,4);
TASK_PP(16'hD0B1,4);
TASK_PP(16'hD0B2,4);
TASK_PP(16'hD0B3,4);
TASK_PP(16'hD0B4,4);
TASK_PP(16'hD0B5,4);
TASK_PP(16'hD0B6,4);
TASK_PP(16'hD0B7,4);
TASK_PP(16'hD0B8,4);
TASK_PP(16'hD0B9,4);
TASK_PP(16'hD0BA,4);
TASK_PP(16'hD0BB,4);
TASK_PP(16'hD0BC,4);
TASK_PP(16'hD0BD,4);
TASK_PP(16'hD0BE,4);
TASK_PP(16'hD0BF,4);
TASK_PP(16'hD0C0,4);
TASK_PP(16'hD0C1,4);
TASK_PP(16'hD0C2,4);
TASK_PP(16'hD0C3,4);
TASK_PP(16'hD0C4,4);
TASK_PP(16'hD0C5,4);
TASK_PP(16'hD0C6,4);
TASK_PP(16'hD0C7,4);
TASK_PP(16'hD0C8,4);
TASK_PP(16'hD0C9,4);
TASK_PP(16'hD0CA,4);
TASK_PP(16'hD0CB,4);
TASK_PP(16'hD0CC,4);
TASK_PP(16'hD0CD,4);
TASK_PP(16'hD0CE,4);
TASK_PP(16'hD0CF,4);
TASK_PP(16'hD0D0,4);
TASK_PP(16'hD0D1,4);
TASK_PP(16'hD0D2,4);
TASK_PP(16'hD0D3,4);
TASK_PP(16'hD0D4,4);
TASK_PP(16'hD0D5,4);
TASK_PP(16'hD0D6,4);
TASK_PP(16'hD0D7,4);
TASK_PP(16'hD0D8,4);
TASK_PP(16'hD0D9,4);
TASK_PP(16'hD0DA,4);
TASK_PP(16'hD0DB,4);
TASK_PP(16'hD0DC,4);
TASK_PP(16'hD0DD,4);
TASK_PP(16'hD0DE,4);
TASK_PP(16'hD0DF,4);
TASK_PP(16'hD0E0,4);
TASK_PP(16'hD0E1,4);
TASK_PP(16'hD0E2,4);
TASK_PP(16'hD0E3,4);
TASK_PP(16'hD0E4,4);
TASK_PP(16'hD0E5,4);
TASK_PP(16'hD0E6,4);
TASK_PP(16'hD0E7,4);
TASK_PP(16'hD0E8,4);
TASK_PP(16'hD0E9,4);
TASK_PP(16'hD0EA,4);
TASK_PP(16'hD0EB,4);
TASK_PP(16'hD0EC,4);
TASK_PP(16'hD0ED,4);
TASK_PP(16'hD0EE,4);
TASK_PP(16'hD0EF,4);
TASK_PP(16'hD0F0,4);
TASK_PP(16'hD0F1,4);
TASK_PP(16'hD0F2,4);
TASK_PP(16'hD0F3,4);
TASK_PP(16'hD0F4,4);
TASK_PP(16'hD0F5,4);
TASK_PP(16'hD0F6,4);
TASK_PP(16'hD0F7,4);
TASK_PP(16'hD0F8,4);
TASK_PP(16'hD0F9,4);
TASK_PP(16'hD0FA,4);
TASK_PP(16'hD0FB,4);
TASK_PP(16'hD0FC,4);
TASK_PP(16'hD0FD,4);
TASK_PP(16'hD0FE,4);
TASK_PP(16'hD0FF,4);
TASK_PP(16'hD100,4);
TASK_PP(16'hD101,4);
TASK_PP(16'hD102,4);
TASK_PP(16'hD103,4);
TASK_PP(16'hD104,4);
TASK_PP(16'hD105,4);
TASK_PP(16'hD106,4);
TASK_PP(16'hD107,4);
TASK_PP(16'hD108,4);
TASK_PP(16'hD109,4);
TASK_PP(16'hD10A,4);
TASK_PP(16'hD10B,4);
TASK_PP(16'hD10C,4);
TASK_PP(16'hD10D,4);
TASK_PP(16'hD10E,4);
TASK_PP(16'hD10F,4);
TASK_PP(16'hD110,4);
TASK_PP(16'hD111,4);
TASK_PP(16'hD112,4);
TASK_PP(16'hD113,4);
TASK_PP(16'hD114,4);
TASK_PP(16'hD115,4);
TASK_PP(16'hD116,4);
TASK_PP(16'hD117,4);
TASK_PP(16'hD118,4);
TASK_PP(16'hD119,4);
TASK_PP(16'hD11A,4);
TASK_PP(16'hD11B,4);
TASK_PP(16'hD11C,4);
TASK_PP(16'hD11D,4);
TASK_PP(16'hD11E,4);
TASK_PP(16'hD11F,4);
TASK_PP(16'hD120,4);
TASK_PP(16'hD121,4);
TASK_PP(16'hD122,4);
TASK_PP(16'hD123,4);
TASK_PP(16'hD124,4);
TASK_PP(16'hD125,4);
TASK_PP(16'hD126,4);
TASK_PP(16'hD127,4);
TASK_PP(16'hD128,4);
TASK_PP(16'hD129,4);
TASK_PP(16'hD12A,4);
TASK_PP(16'hD12B,4);
TASK_PP(16'hD12C,4);
TASK_PP(16'hD12D,4);
TASK_PP(16'hD12E,4);
TASK_PP(16'hD12F,4);
TASK_PP(16'hD130,4);
TASK_PP(16'hD131,4);
TASK_PP(16'hD132,4);
TASK_PP(16'hD133,4);
TASK_PP(16'hD134,4);
TASK_PP(16'hD135,4);
TASK_PP(16'hD136,4);
TASK_PP(16'hD137,4);
TASK_PP(16'hD138,4);
TASK_PP(16'hD139,4);
TASK_PP(16'hD13A,4);
TASK_PP(16'hD13B,4);
TASK_PP(16'hD13C,4);
TASK_PP(16'hD13D,4);
TASK_PP(16'hD13E,4);
TASK_PP(16'hD13F,4);
TASK_PP(16'hD140,4);
TASK_PP(16'hD141,4);
TASK_PP(16'hD142,4);
TASK_PP(16'hD143,4);
TASK_PP(16'hD144,4);
TASK_PP(16'hD145,4);
TASK_PP(16'hD146,4);
TASK_PP(16'hD147,4);
TASK_PP(16'hD148,4);
TASK_PP(16'hD149,4);
TASK_PP(16'hD14A,4);
TASK_PP(16'hD14B,4);
TASK_PP(16'hD14C,4);
TASK_PP(16'hD14D,4);
TASK_PP(16'hD14E,4);
TASK_PP(16'hD14F,4);
TASK_PP(16'hD150,4);
TASK_PP(16'hD151,4);
TASK_PP(16'hD152,4);
TASK_PP(16'hD153,4);
TASK_PP(16'hD154,4);
TASK_PP(16'hD155,4);
TASK_PP(16'hD156,4);
TASK_PP(16'hD157,4);
TASK_PP(16'hD158,4);
TASK_PP(16'hD159,4);
TASK_PP(16'hD15A,4);
TASK_PP(16'hD15B,4);
TASK_PP(16'hD15C,4);
TASK_PP(16'hD15D,4);
TASK_PP(16'hD15E,4);
TASK_PP(16'hD15F,4);
TASK_PP(16'hD160,4);
TASK_PP(16'hD161,4);
TASK_PP(16'hD162,4);
TASK_PP(16'hD163,4);
TASK_PP(16'hD164,4);
TASK_PP(16'hD165,4);
TASK_PP(16'hD166,4);
TASK_PP(16'hD167,4);
TASK_PP(16'hD168,4);
TASK_PP(16'hD169,4);
TASK_PP(16'hD16A,4);
TASK_PP(16'hD16B,4);
TASK_PP(16'hD16C,4);
TASK_PP(16'hD16D,4);
TASK_PP(16'hD16E,4);
TASK_PP(16'hD16F,4);
TASK_PP(16'hD170,4);
TASK_PP(16'hD171,4);
TASK_PP(16'hD172,4);
TASK_PP(16'hD173,4);
TASK_PP(16'hD174,4);
TASK_PP(16'hD175,4);
TASK_PP(16'hD176,4);
TASK_PP(16'hD177,4);
TASK_PP(16'hD178,4);
TASK_PP(16'hD179,4);
TASK_PP(16'hD17A,4);
TASK_PP(16'hD17B,4);
TASK_PP(16'hD17C,4);
TASK_PP(16'hD17D,4);
TASK_PP(16'hD17E,4);
TASK_PP(16'hD17F,4);
TASK_PP(16'hD180,4);
TASK_PP(16'hD181,4);
TASK_PP(16'hD182,4);
TASK_PP(16'hD183,4);
TASK_PP(16'hD184,4);
TASK_PP(16'hD185,4);
TASK_PP(16'hD186,4);
TASK_PP(16'hD187,4);
TASK_PP(16'hD188,4);
TASK_PP(16'hD189,4);
TASK_PP(16'hD18A,4);
TASK_PP(16'hD18B,4);
TASK_PP(16'hD18C,4);
TASK_PP(16'hD18D,4);
TASK_PP(16'hD18E,4);
TASK_PP(16'hD18F,4);
TASK_PP(16'hD190,4);
TASK_PP(16'hD191,4);
TASK_PP(16'hD192,4);
TASK_PP(16'hD193,4);
TASK_PP(16'hD194,4);
TASK_PP(16'hD195,4);
TASK_PP(16'hD196,4);
TASK_PP(16'hD197,4);
TASK_PP(16'hD198,4);
TASK_PP(16'hD199,4);
TASK_PP(16'hD19A,4);
TASK_PP(16'hD19B,4);
TASK_PP(16'hD19C,4);
TASK_PP(16'hD19D,4);
TASK_PP(16'hD19E,4);
TASK_PP(16'hD19F,4);
TASK_PP(16'hD1A0,4);
TASK_PP(16'hD1A1,4);
TASK_PP(16'hD1A2,4);
TASK_PP(16'hD1A3,4);
TASK_PP(16'hD1A4,4);
TASK_PP(16'hD1A5,4);
TASK_PP(16'hD1A6,4);
TASK_PP(16'hD1A7,4);
TASK_PP(16'hD1A8,4);
TASK_PP(16'hD1A9,4);
TASK_PP(16'hD1AA,4);
TASK_PP(16'hD1AB,4);
TASK_PP(16'hD1AC,4);
TASK_PP(16'hD1AD,4);
TASK_PP(16'hD1AE,4);
TASK_PP(16'hD1AF,4);
TASK_PP(16'hD1B0,4);
TASK_PP(16'hD1B1,4);
TASK_PP(16'hD1B2,4);
TASK_PP(16'hD1B3,4);
TASK_PP(16'hD1B4,4);
TASK_PP(16'hD1B5,4);
TASK_PP(16'hD1B6,4);
TASK_PP(16'hD1B7,4);
TASK_PP(16'hD1B8,4);
TASK_PP(16'hD1B9,4);
TASK_PP(16'hD1BA,4);
TASK_PP(16'hD1BB,4);
TASK_PP(16'hD1BC,4);
TASK_PP(16'hD1BD,4);
TASK_PP(16'hD1BE,4);
TASK_PP(16'hD1BF,4);
TASK_PP(16'hD1C0,4);
TASK_PP(16'hD1C1,4);
TASK_PP(16'hD1C2,4);
TASK_PP(16'hD1C3,4);
TASK_PP(16'hD1C4,4);
TASK_PP(16'hD1C5,4);
TASK_PP(16'hD1C6,4);
TASK_PP(16'hD1C7,4);
TASK_PP(16'hD1C8,4);
TASK_PP(16'hD1C9,4);
TASK_PP(16'hD1CA,4);
TASK_PP(16'hD1CB,4);
TASK_PP(16'hD1CC,4);
TASK_PP(16'hD1CD,4);
TASK_PP(16'hD1CE,4);
TASK_PP(16'hD1CF,4);
TASK_PP(16'hD1D0,4);
TASK_PP(16'hD1D1,4);
TASK_PP(16'hD1D2,4);
TASK_PP(16'hD1D3,4);
TASK_PP(16'hD1D4,4);
TASK_PP(16'hD1D5,4);
TASK_PP(16'hD1D6,4);
TASK_PP(16'hD1D7,4);
TASK_PP(16'hD1D8,4);
TASK_PP(16'hD1D9,4);
TASK_PP(16'hD1DA,4);
TASK_PP(16'hD1DB,4);
TASK_PP(16'hD1DC,4);
TASK_PP(16'hD1DD,4);
TASK_PP(16'hD1DE,4);
TASK_PP(16'hD1DF,4);
TASK_PP(16'hD1E0,4);
TASK_PP(16'hD1E1,4);
TASK_PP(16'hD1E2,4);
TASK_PP(16'hD1E3,4);
TASK_PP(16'hD1E4,4);
TASK_PP(16'hD1E5,4);
TASK_PP(16'hD1E6,4);
TASK_PP(16'hD1E7,4);
TASK_PP(16'hD1E8,4);
TASK_PP(16'hD1E9,4);
TASK_PP(16'hD1EA,4);
TASK_PP(16'hD1EB,4);
TASK_PP(16'hD1EC,4);
TASK_PP(16'hD1ED,4);
TASK_PP(16'hD1EE,4);
TASK_PP(16'hD1EF,4);
TASK_PP(16'hD1F0,4);
TASK_PP(16'hD1F1,4);
TASK_PP(16'hD1F2,4);
TASK_PP(16'hD1F3,4);
TASK_PP(16'hD1F4,4);
TASK_PP(16'hD1F5,4);
TASK_PP(16'hD1F6,4);
TASK_PP(16'hD1F7,4);
TASK_PP(16'hD1F8,4);
TASK_PP(16'hD1F9,4);
TASK_PP(16'hD1FA,4);
TASK_PP(16'hD1FB,4);
TASK_PP(16'hD1FC,4);
TASK_PP(16'hD1FD,4);
TASK_PP(16'hD1FE,4);
TASK_PP(16'hD1FF,4);
TASK_PP(16'hD200,4);
TASK_PP(16'hD201,4);
TASK_PP(16'hD202,4);
TASK_PP(16'hD203,4);
TASK_PP(16'hD204,4);
TASK_PP(16'hD205,4);
TASK_PP(16'hD206,4);
TASK_PP(16'hD207,4);
TASK_PP(16'hD208,4);
TASK_PP(16'hD209,4);
TASK_PP(16'hD20A,4);
TASK_PP(16'hD20B,4);
TASK_PP(16'hD20C,4);
TASK_PP(16'hD20D,4);
TASK_PP(16'hD20E,4);
TASK_PP(16'hD20F,4);
TASK_PP(16'hD210,4);
TASK_PP(16'hD211,4);
TASK_PP(16'hD212,4);
TASK_PP(16'hD213,4);
TASK_PP(16'hD214,4);
TASK_PP(16'hD215,4);
TASK_PP(16'hD216,4);
TASK_PP(16'hD217,4);
TASK_PP(16'hD218,4);
TASK_PP(16'hD219,4);
TASK_PP(16'hD21A,4);
TASK_PP(16'hD21B,4);
TASK_PP(16'hD21C,4);
TASK_PP(16'hD21D,4);
TASK_PP(16'hD21E,4);
TASK_PP(16'hD21F,4);
TASK_PP(16'hD220,4);
TASK_PP(16'hD221,4);
TASK_PP(16'hD222,4);
TASK_PP(16'hD223,4);
TASK_PP(16'hD224,4);
TASK_PP(16'hD225,4);
TASK_PP(16'hD226,4);
TASK_PP(16'hD227,4);
TASK_PP(16'hD228,4);
TASK_PP(16'hD229,4);
TASK_PP(16'hD22A,4);
TASK_PP(16'hD22B,4);
TASK_PP(16'hD22C,4);
TASK_PP(16'hD22D,4);
TASK_PP(16'hD22E,4);
TASK_PP(16'hD22F,4);
TASK_PP(16'hD230,4);
TASK_PP(16'hD231,4);
TASK_PP(16'hD232,4);
TASK_PP(16'hD233,4);
TASK_PP(16'hD234,4);
TASK_PP(16'hD235,4);
TASK_PP(16'hD236,4);
TASK_PP(16'hD237,4);
TASK_PP(16'hD238,4);
TASK_PP(16'hD239,4);
TASK_PP(16'hD23A,4);
TASK_PP(16'hD23B,4);
TASK_PP(16'hD23C,4);
TASK_PP(16'hD23D,4);
TASK_PP(16'hD23E,4);
TASK_PP(16'hD23F,4);
TASK_PP(16'hD240,4);
TASK_PP(16'hD241,4);
TASK_PP(16'hD242,4);
TASK_PP(16'hD243,4);
TASK_PP(16'hD244,4);
TASK_PP(16'hD245,4);
TASK_PP(16'hD246,4);
TASK_PP(16'hD247,4);
TASK_PP(16'hD248,4);
TASK_PP(16'hD249,4);
TASK_PP(16'hD24A,4);
TASK_PP(16'hD24B,4);
TASK_PP(16'hD24C,4);
TASK_PP(16'hD24D,4);
TASK_PP(16'hD24E,4);
TASK_PP(16'hD24F,4);
TASK_PP(16'hD250,4);
TASK_PP(16'hD251,4);
TASK_PP(16'hD252,4);
TASK_PP(16'hD253,4);
TASK_PP(16'hD254,4);
TASK_PP(16'hD255,4);
TASK_PP(16'hD256,4);
TASK_PP(16'hD257,4);
TASK_PP(16'hD258,4);
TASK_PP(16'hD259,4);
TASK_PP(16'hD25A,4);
TASK_PP(16'hD25B,4);
TASK_PP(16'hD25C,4);
TASK_PP(16'hD25D,4);
TASK_PP(16'hD25E,4);
TASK_PP(16'hD25F,4);
TASK_PP(16'hD260,4);
TASK_PP(16'hD261,4);
TASK_PP(16'hD262,4);
TASK_PP(16'hD263,4);
TASK_PP(16'hD264,4);
TASK_PP(16'hD265,4);
TASK_PP(16'hD266,4);
TASK_PP(16'hD267,4);
TASK_PP(16'hD268,4);
TASK_PP(16'hD269,4);
TASK_PP(16'hD26A,4);
TASK_PP(16'hD26B,4);
TASK_PP(16'hD26C,4);
TASK_PP(16'hD26D,4);
TASK_PP(16'hD26E,4);
TASK_PP(16'hD26F,4);
TASK_PP(16'hD270,4);
TASK_PP(16'hD271,4);
TASK_PP(16'hD272,4);
TASK_PP(16'hD273,4);
TASK_PP(16'hD274,4);
TASK_PP(16'hD275,4);
TASK_PP(16'hD276,4);
TASK_PP(16'hD277,4);
TASK_PP(16'hD278,4);
TASK_PP(16'hD279,4);
TASK_PP(16'hD27A,4);
TASK_PP(16'hD27B,4);
TASK_PP(16'hD27C,4);
TASK_PP(16'hD27D,4);
TASK_PP(16'hD27E,4);
TASK_PP(16'hD27F,4);
TASK_PP(16'hD280,4);
TASK_PP(16'hD281,4);
TASK_PP(16'hD282,4);
TASK_PP(16'hD283,4);
TASK_PP(16'hD284,4);
TASK_PP(16'hD285,4);
TASK_PP(16'hD286,4);
TASK_PP(16'hD287,4);
TASK_PP(16'hD288,4);
TASK_PP(16'hD289,4);
TASK_PP(16'hD28A,4);
TASK_PP(16'hD28B,4);
TASK_PP(16'hD28C,4);
TASK_PP(16'hD28D,4);
TASK_PP(16'hD28E,4);
TASK_PP(16'hD28F,4);
TASK_PP(16'hD290,4);
TASK_PP(16'hD291,4);
TASK_PP(16'hD292,4);
TASK_PP(16'hD293,4);
TASK_PP(16'hD294,4);
TASK_PP(16'hD295,4);
TASK_PP(16'hD296,4);
TASK_PP(16'hD297,4);
TASK_PP(16'hD298,4);
TASK_PP(16'hD299,4);
TASK_PP(16'hD29A,4);
TASK_PP(16'hD29B,4);
TASK_PP(16'hD29C,4);
TASK_PP(16'hD29D,4);
TASK_PP(16'hD29E,4);
TASK_PP(16'hD29F,4);
TASK_PP(16'hD2A0,4);
TASK_PP(16'hD2A1,4);
TASK_PP(16'hD2A2,4);
TASK_PP(16'hD2A3,4);
TASK_PP(16'hD2A4,4);
TASK_PP(16'hD2A5,4);
TASK_PP(16'hD2A6,4);
TASK_PP(16'hD2A7,4);
TASK_PP(16'hD2A8,4);
TASK_PP(16'hD2A9,4);
TASK_PP(16'hD2AA,4);
TASK_PP(16'hD2AB,4);
TASK_PP(16'hD2AC,4);
TASK_PP(16'hD2AD,4);
TASK_PP(16'hD2AE,4);
TASK_PP(16'hD2AF,4);
TASK_PP(16'hD2B0,4);
TASK_PP(16'hD2B1,4);
TASK_PP(16'hD2B2,4);
TASK_PP(16'hD2B3,4);
TASK_PP(16'hD2B4,4);
TASK_PP(16'hD2B5,4);
TASK_PP(16'hD2B6,4);
TASK_PP(16'hD2B7,4);
TASK_PP(16'hD2B8,4);
TASK_PP(16'hD2B9,4);
TASK_PP(16'hD2BA,4);
TASK_PP(16'hD2BB,4);
TASK_PP(16'hD2BC,4);
TASK_PP(16'hD2BD,4);
TASK_PP(16'hD2BE,4);
TASK_PP(16'hD2BF,4);
TASK_PP(16'hD2C0,4);
TASK_PP(16'hD2C1,4);
TASK_PP(16'hD2C2,4);
TASK_PP(16'hD2C3,4);
TASK_PP(16'hD2C4,4);
TASK_PP(16'hD2C5,4);
TASK_PP(16'hD2C6,4);
TASK_PP(16'hD2C7,4);
TASK_PP(16'hD2C8,4);
TASK_PP(16'hD2C9,4);
TASK_PP(16'hD2CA,4);
TASK_PP(16'hD2CB,4);
TASK_PP(16'hD2CC,4);
TASK_PP(16'hD2CD,4);
TASK_PP(16'hD2CE,4);
TASK_PP(16'hD2CF,4);
TASK_PP(16'hD2D0,4);
TASK_PP(16'hD2D1,4);
TASK_PP(16'hD2D2,4);
TASK_PP(16'hD2D3,4);
TASK_PP(16'hD2D4,4);
TASK_PP(16'hD2D5,4);
TASK_PP(16'hD2D6,4);
TASK_PP(16'hD2D7,4);
TASK_PP(16'hD2D8,4);
TASK_PP(16'hD2D9,4);
TASK_PP(16'hD2DA,4);
TASK_PP(16'hD2DB,4);
TASK_PP(16'hD2DC,4);
TASK_PP(16'hD2DD,4);
TASK_PP(16'hD2DE,4);
TASK_PP(16'hD2DF,4);
TASK_PP(16'hD2E0,4);
TASK_PP(16'hD2E1,4);
TASK_PP(16'hD2E2,4);
TASK_PP(16'hD2E3,4);
TASK_PP(16'hD2E4,4);
TASK_PP(16'hD2E5,4);
TASK_PP(16'hD2E6,4);
TASK_PP(16'hD2E7,4);
TASK_PP(16'hD2E8,4);
TASK_PP(16'hD2E9,4);
TASK_PP(16'hD2EA,4);
TASK_PP(16'hD2EB,4);
TASK_PP(16'hD2EC,4);
TASK_PP(16'hD2ED,4);
TASK_PP(16'hD2EE,4);
TASK_PP(16'hD2EF,4);
TASK_PP(16'hD2F0,4);
TASK_PP(16'hD2F1,4);
TASK_PP(16'hD2F2,4);
TASK_PP(16'hD2F3,4);
TASK_PP(16'hD2F4,4);
TASK_PP(16'hD2F5,4);
TASK_PP(16'hD2F6,4);
TASK_PP(16'hD2F7,4);
TASK_PP(16'hD2F8,4);
TASK_PP(16'hD2F9,4);
TASK_PP(16'hD2FA,4);
TASK_PP(16'hD2FB,4);
TASK_PP(16'hD2FC,4);
TASK_PP(16'hD2FD,4);
TASK_PP(16'hD2FE,4);
TASK_PP(16'hD2FF,4);
TASK_PP(16'hD300,4);
TASK_PP(16'hD301,4);
TASK_PP(16'hD302,4);
TASK_PP(16'hD303,4);
TASK_PP(16'hD304,4);
TASK_PP(16'hD305,4);
TASK_PP(16'hD306,4);
TASK_PP(16'hD307,4);
TASK_PP(16'hD308,4);
TASK_PP(16'hD309,4);
TASK_PP(16'hD30A,4);
TASK_PP(16'hD30B,4);
TASK_PP(16'hD30C,4);
TASK_PP(16'hD30D,4);
TASK_PP(16'hD30E,4);
TASK_PP(16'hD30F,4);
TASK_PP(16'hD310,4);
TASK_PP(16'hD311,4);
TASK_PP(16'hD312,4);
TASK_PP(16'hD313,4);
TASK_PP(16'hD314,4);
TASK_PP(16'hD315,4);
TASK_PP(16'hD316,4);
TASK_PP(16'hD317,4);
TASK_PP(16'hD318,4);
TASK_PP(16'hD319,4);
TASK_PP(16'hD31A,4);
TASK_PP(16'hD31B,4);
TASK_PP(16'hD31C,4);
TASK_PP(16'hD31D,4);
TASK_PP(16'hD31E,4);
TASK_PP(16'hD31F,4);
TASK_PP(16'hD320,4);
TASK_PP(16'hD321,4);
TASK_PP(16'hD322,4);
TASK_PP(16'hD323,4);
TASK_PP(16'hD324,4);
TASK_PP(16'hD325,4);
TASK_PP(16'hD326,4);
TASK_PP(16'hD327,4);
TASK_PP(16'hD328,4);
TASK_PP(16'hD329,4);
TASK_PP(16'hD32A,4);
TASK_PP(16'hD32B,4);
TASK_PP(16'hD32C,4);
TASK_PP(16'hD32D,4);
TASK_PP(16'hD32E,4);
TASK_PP(16'hD32F,4);
TASK_PP(16'hD330,4);
TASK_PP(16'hD331,4);
TASK_PP(16'hD332,4);
TASK_PP(16'hD333,4);
TASK_PP(16'hD334,4);
TASK_PP(16'hD335,4);
TASK_PP(16'hD336,4);
TASK_PP(16'hD337,4);
TASK_PP(16'hD338,4);
TASK_PP(16'hD339,4);
TASK_PP(16'hD33A,4);
TASK_PP(16'hD33B,4);
TASK_PP(16'hD33C,4);
TASK_PP(16'hD33D,4);
TASK_PP(16'hD33E,4);
TASK_PP(16'hD33F,4);
TASK_PP(16'hD340,4);
TASK_PP(16'hD341,4);
TASK_PP(16'hD342,4);
TASK_PP(16'hD343,4);
TASK_PP(16'hD344,4);
TASK_PP(16'hD345,4);
TASK_PP(16'hD346,4);
TASK_PP(16'hD347,4);
TASK_PP(16'hD348,4);
TASK_PP(16'hD349,4);
TASK_PP(16'hD34A,4);
TASK_PP(16'hD34B,4);
TASK_PP(16'hD34C,4);
TASK_PP(16'hD34D,4);
TASK_PP(16'hD34E,4);
TASK_PP(16'hD34F,4);
TASK_PP(16'hD350,4);
TASK_PP(16'hD351,4);
TASK_PP(16'hD352,4);
TASK_PP(16'hD353,4);
TASK_PP(16'hD354,4);
TASK_PP(16'hD355,4);
TASK_PP(16'hD356,4);
TASK_PP(16'hD357,4);
TASK_PP(16'hD358,4);
TASK_PP(16'hD359,4);
TASK_PP(16'hD35A,4);
TASK_PP(16'hD35B,4);
TASK_PP(16'hD35C,4);
TASK_PP(16'hD35D,4);
TASK_PP(16'hD35E,4);
TASK_PP(16'hD35F,4);
TASK_PP(16'hD360,4);
TASK_PP(16'hD361,4);
TASK_PP(16'hD362,4);
TASK_PP(16'hD363,4);
TASK_PP(16'hD364,4);
TASK_PP(16'hD365,4);
TASK_PP(16'hD366,4);
TASK_PP(16'hD367,4);
TASK_PP(16'hD368,4);
TASK_PP(16'hD369,4);
TASK_PP(16'hD36A,4);
TASK_PP(16'hD36B,4);
TASK_PP(16'hD36C,4);
TASK_PP(16'hD36D,4);
TASK_PP(16'hD36E,4);
TASK_PP(16'hD36F,4);
TASK_PP(16'hD370,4);
TASK_PP(16'hD371,4);
TASK_PP(16'hD372,4);
TASK_PP(16'hD373,4);
TASK_PP(16'hD374,4);
TASK_PP(16'hD375,4);
TASK_PP(16'hD376,4);
TASK_PP(16'hD377,4);
TASK_PP(16'hD378,4);
TASK_PP(16'hD379,4);
TASK_PP(16'hD37A,4);
TASK_PP(16'hD37B,4);
TASK_PP(16'hD37C,4);
TASK_PP(16'hD37D,4);
TASK_PP(16'hD37E,4);
TASK_PP(16'hD37F,4);
TASK_PP(16'hD380,4);
TASK_PP(16'hD381,4);
TASK_PP(16'hD382,4);
TASK_PP(16'hD383,4);
TASK_PP(16'hD384,4);
TASK_PP(16'hD385,4);
TASK_PP(16'hD386,4);
TASK_PP(16'hD387,4);
TASK_PP(16'hD388,4);
TASK_PP(16'hD389,4);
TASK_PP(16'hD38A,4);
TASK_PP(16'hD38B,4);
TASK_PP(16'hD38C,4);
TASK_PP(16'hD38D,4);
TASK_PP(16'hD38E,4);
TASK_PP(16'hD38F,4);
TASK_PP(16'hD390,4);
TASK_PP(16'hD391,4);
TASK_PP(16'hD392,4);
TASK_PP(16'hD393,4);
TASK_PP(16'hD394,4);
TASK_PP(16'hD395,4);
TASK_PP(16'hD396,4);
TASK_PP(16'hD397,4);
TASK_PP(16'hD398,4);
TASK_PP(16'hD399,4);
TASK_PP(16'hD39A,4);
TASK_PP(16'hD39B,4);
TASK_PP(16'hD39C,4);
TASK_PP(16'hD39D,4);
TASK_PP(16'hD39E,4);
TASK_PP(16'hD39F,4);
TASK_PP(16'hD3A0,4);
TASK_PP(16'hD3A1,4);
TASK_PP(16'hD3A2,4);
TASK_PP(16'hD3A3,4);
TASK_PP(16'hD3A4,4);
TASK_PP(16'hD3A5,4);
TASK_PP(16'hD3A6,4);
TASK_PP(16'hD3A7,4);
TASK_PP(16'hD3A8,4);
TASK_PP(16'hD3A9,4);
TASK_PP(16'hD3AA,4);
TASK_PP(16'hD3AB,4);
TASK_PP(16'hD3AC,4);
TASK_PP(16'hD3AD,4);
TASK_PP(16'hD3AE,4);
TASK_PP(16'hD3AF,4);
TASK_PP(16'hD3B0,4);
TASK_PP(16'hD3B1,4);
TASK_PP(16'hD3B2,4);
TASK_PP(16'hD3B3,4);
TASK_PP(16'hD3B4,4);
TASK_PP(16'hD3B5,4);
TASK_PP(16'hD3B6,4);
TASK_PP(16'hD3B7,4);
TASK_PP(16'hD3B8,4);
TASK_PP(16'hD3B9,4);
TASK_PP(16'hD3BA,4);
TASK_PP(16'hD3BB,4);
TASK_PP(16'hD3BC,4);
TASK_PP(16'hD3BD,4);
TASK_PP(16'hD3BE,4);
TASK_PP(16'hD3BF,4);
TASK_PP(16'hD3C0,4);
TASK_PP(16'hD3C1,4);
TASK_PP(16'hD3C2,4);
TASK_PP(16'hD3C3,4);
TASK_PP(16'hD3C4,4);
TASK_PP(16'hD3C5,4);
TASK_PP(16'hD3C6,4);
TASK_PP(16'hD3C7,4);
TASK_PP(16'hD3C8,4);
TASK_PP(16'hD3C9,4);
TASK_PP(16'hD3CA,4);
TASK_PP(16'hD3CB,4);
TASK_PP(16'hD3CC,4);
TASK_PP(16'hD3CD,4);
TASK_PP(16'hD3CE,4);
TASK_PP(16'hD3CF,4);
TASK_PP(16'hD3D0,4);
TASK_PP(16'hD3D1,4);
TASK_PP(16'hD3D2,4);
TASK_PP(16'hD3D3,4);
TASK_PP(16'hD3D4,4);
TASK_PP(16'hD3D5,4);
TASK_PP(16'hD3D6,4);
TASK_PP(16'hD3D7,4);
TASK_PP(16'hD3D8,4);
TASK_PP(16'hD3D9,4);
TASK_PP(16'hD3DA,4);
TASK_PP(16'hD3DB,4);
TASK_PP(16'hD3DC,4);
TASK_PP(16'hD3DD,4);
TASK_PP(16'hD3DE,4);
TASK_PP(16'hD3DF,4);
TASK_PP(16'hD3E0,4);
TASK_PP(16'hD3E1,4);
TASK_PP(16'hD3E2,4);
TASK_PP(16'hD3E3,4);
TASK_PP(16'hD3E4,4);
TASK_PP(16'hD3E5,4);
TASK_PP(16'hD3E6,4);
TASK_PP(16'hD3E7,4);
TASK_PP(16'hD3E8,4);
TASK_PP(16'hD3E9,4);
TASK_PP(16'hD3EA,4);
TASK_PP(16'hD3EB,4);
TASK_PP(16'hD3EC,4);
TASK_PP(16'hD3ED,4);
TASK_PP(16'hD3EE,4);
TASK_PP(16'hD3EF,4);
TASK_PP(16'hD3F0,4);
TASK_PP(16'hD3F1,4);
TASK_PP(16'hD3F2,4);
TASK_PP(16'hD3F3,4);
TASK_PP(16'hD3F4,4);
TASK_PP(16'hD3F5,4);
TASK_PP(16'hD3F6,4);
TASK_PP(16'hD3F7,4);
TASK_PP(16'hD3F8,4);
TASK_PP(16'hD3F9,4);
TASK_PP(16'hD3FA,4);
TASK_PP(16'hD3FB,4);
TASK_PP(16'hD3FC,4);
TASK_PP(16'hD3FD,4);
TASK_PP(16'hD3FE,4);
TASK_PP(16'hD3FF,4);
TASK_PP(16'hD400,4);
TASK_PP(16'hD401,4);
TASK_PP(16'hD402,4);
TASK_PP(16'hD403,4);
TASK_PP(16'hD404,4);
TASK_PP(16'hD405,4);
TASK_PP(16'hD406,4);
TASK_PP(16'hD407,4);
TASK_PP(16'hD408,4);
TASK_PP(16'hD409,4);
TASK_PP(16'hD40A,4);
TASK_PP(16'hD40B,4);
TASK_PP(16'hD40C,4);
TASK_PP(16'hD40D,4);
TASK_PP(16'hD40E,4);
TASK_PP(16'hD40F,4);
TASK_PP(16'hD410,4);
TASK_PP(16'hD411,4);
TASK_PP(16'hD412,4);
TASK_PP(16'hD413,4);
TASK_PP(16'hD414,4);
TASK_PP(16'hD415,4);
TASK_PP(16'hD416,4);
TASK_PP(16'hD417,4);
TASK_PP(16'hD418,4);
TASK_PP(16'hD419,4);
TASK_PP(16'hD41A,4);
TASK_PP(16'hD41B,4);
TASK_PP(16'hD41C,4);
TASK_PP(16'hD41D,4);
TASK_PP(16'hD41E,4);
TASK_PP(16'hD41F,4);
TASK_PP(16'hD420,4);
TASK_PP(16'hD421,4);
TASK_PP(16'hD422,4);
TASK_PP(16'hD423,4);
TASK_PP(16'hD424,4);
TASK_PP(16'hD425,4);
TASK_PP(16'hD426,4);
TASK_PP(16'hD427,4);
TASK_PP(16'hD428,4);
TASK_PP(16'hD429,4);
TASK_PP(16'hD42A,4);
TASK_PP(16'hD42B,4);
TASK_PP(16'hD42C,4);
TASK_PP(16'hD42D,4);
TASK_PP(16'hD42E,4);
TASK_PP(16'hD42F,4);
TASK_PP(16'hD430,4);
TASK_PP(16'hD431,4);
TASK_PP(16'hD432,4);
TASK_PP(16'hD433,4);
TASK_PP(16'hD434,4);
TASK_PP(16'hD435,4);
TASK_PP(16'hD436,4);
TASK_PP(16'hD437,4);
TASK_PP(16'hD438,4);
TASK_PP(16'hD439,4);
TASK_PP(16'hD43A,4);
TASK_PP(16'hD43B,4);
TASK_PP(16'hD43C,4);
TASK_PP(16'hD43D,4);
TASK_PP(16'hD43E,4);
TASK_PP(16'hD43F,4);
TASK_PP(16'hD440,4);
TASK_PP(16'hD441,4);
TASK_PP(16'hD442,4);
TASK_PP(16'hD443,4);
TASK_PP(16'hD444,4);
TASK_PP(16'hD445,4);
TASK_PP(16'hD446,4);
TASK_PP(16'hD447,4);
TASK_PP(16'hD448,4);
TASK_PP(16'hD449,4);
TASK_PP(16'hD44A,4);
TASK_PP(16'hD44B,4);
TASK_PP(16'hD44C,4);
TASK_PP(16'hD44D,4);
TASK_PP(16'hD44E,4);
TASK_PP(16'hD44F,4);
TASK_PP(16'hD450,4);
TASK_PP(16'hD451,4);
TASK_PP(16'hD452,4);
TASK_PP(16'hD453,4);
TASK_PP(16'hD454,4);
TASK_PP(16'hD455,4);
TASK_PP(16'hD456,4);
TASK_PP(16'hD457,4);
TASK_PP(16'hD458,4);
TASK_PP(16'hD459,4);
TASK_PP(16'hD45A,4);
TASK_PP(16'hD45B,4);
TASK_PP(16'hD45C,4);
TASK_PP(16'hD45D,4);
TASK_PP(16'hD45E,4);
TASK_PP(16'hD45F,4);
TASK_PP(16'hD460,4);
TASK_PP(16'hD461,4);
TASK_PP(16'hD462,4);
TASK_PP(16'hD463,4);
TASK_PP(16'hD464,4);
TASK_PP(16'hD465,4);
TASK_PP(16'hD466,4);
TASK_PP(16'hD467,4);
TASK_PP(16'hD468,4);
TASK_PP(16'hD469,4);
TASK_PP(16'hD46A,4);
TASK_PP(16'hD46B,4);
TASK_PP(16'hD46C,4);
TASK_PP(16'hD46D,4);
TASK_PP(16'hD46E,4);
TASK_PP(16'hD46F,4);
TASK_PP(16'hD470,4);
TASK_PP(16'hD471,4);
TASK_PP(16'hD472,4);
TASK_PP(16'hD473,4);
TASK_PP(16'hD474,4);
TASK_PP(16'hD475,4);
TASK_PP(16'hD476,4);
TASK_PP(16'hD477,4);
TASK_PP(16'hD478,4);
TASK_PP(16'hD479,4);
TASK_PP(16'hD47A,4);
TASK_PP(16'hD47B,4);
TASK_PP(16'hD47C,4);
TASK_PP(16'hD47D,4);
TASK_PP(16'hD47E,4);
TASK_PP(16'hD47F,4);
TASK_PP(16'hD480,4);
TASK_PP(16'hD481,4);
TASK_PP(16'hD482,4);
TASK_PP(16'hD483,4);
TASK_PP(16'hD484,4);
TASK_PP(16'hD485,4);
TASK_PP(16'hD486,4);
TASK_PP(16'hD487,4);
TASK_PP(16'hD488,4);
TASK_PP(16'hD489,4);
TASK_PP(16'hD48A,4);
TASK_PP(16'hD48B,4);
TASK_PP(16'hD48C,4);
TASK_PP(16'hD48D,4);
TASK_PP(16'hD48E,4);
TASK_PP(16'hD48F,4);
TASK_PP(16'hD490,4);
TASK_PP(16'hD491,4);
TASK_PP(16'hD492,4);
TASK_PP(16'hD493,4);
TASK_PP(16'hD494,4);
TASK_PP(16'hD495,4);
TASK_PP(16'hD496,4);
TASK_PP(16'hD497,4);
TASK_PP(16'hD498,4);
TASK_PP(16'hD499,4);
TASK_PP(16'hD49A,4);
TASK_PP(16'hD49B,4);
TASK_PP(16'hD49C,4);
TASK_PP(16'hD49D,4);
TASK_PP(16'hD49E,4);
TASK_PP(16'hD49F,4);
TASK_PP(16'hD4A0,4);
TASK_PP(16'hD4A1,4);
TASK_PP(16'hD4A2,4);
TASK_PP(16'hD4A3,4);
TASK_PP(16'hD4A4,4);
TASK_PP(16'hD4A5,4);
TASK_PP(16'hD4A6,4);
TASK_PP(16'hD4A7,4);
TASK_PP(16'hD4A8,4);
TASK_PP(16'hD4A9,4);
TASK_PP(16'hD4AA,4);
TASK_PP(16'hD4AB,4);
TASK_PP(16'hD4AC,4);
TASK_PP(16'hD4AD,4);
TASK_PP(16'hD4AE,4);
TASK_PP(16'hD4AF,4);
TASK_PP(16'hD4B0,4);
TASK_PP(16'hD4B1,4);
TASK_PP(16'hD4B2,4);
TASK_PP(16'hD4B3,4);
TASK_PP(16'hD4B4,4);
TASK_PP(16'hD4B5,4);
TASK_PP(16'hD4B6,4);
TASK_PP(16'hD4B7,4);
TASK_PP(16'hD4B8,4);
TASK_PP(16'hD4B9,4);
TASK_PP(16'hD4BA,4);
TASK_PP(16'hD4BB,4);
TASK_PP(16'hD4BC,4);
TASK_PP(16'hD4BD,4);
TASK_PP(16'hD4BE,4);
TASK_PP(16'hD4BF,4);
TASK_PP(16'hD4C0,4);
TASK_PP(16'hD4C1,4);
TASK_PP(16'hD4C2,4);
TASK_PP(16'hD4C3,4);
TASK_PP(16'hD4C4,4);
TASK_PP(16'hD4C5,4);
TASK_PP(16'hD4C6,4);
TASK_PP(16'hD4C7,4);
TASK_PP(16'hD4C8,4);
TASK_PP(16'hD4C9,4);
TASK_PP(16'hD4CA,4);
TASK_PP(16'hD4CB,4);
TASK_PP(16'hD4CC,4);
TASK_PP(16'hD4CD,4);
TASK_PP(16'hD4CE,4);
TASK_PP(16'hD4CF,4);
TASK_PP(16'hD4D0,4);
TASK_PP(16'hD4D1,4);
TASK_PP(16'hD4D2,4);
TASK_PP(16'hD4D3,4);
TASK_PP(16'hD4D4,4);
TASK_PP(16'hD4D5,4);
TASK_PP(16'hD4D6,4);
TASK_PP(16'hD4D7,4);
TASK_PP(16'hD4D8,4);
TASK_PP(16'hD4D9,4);
TASK_PP(16'hD4DA,4);
TASK_PP(16'hD4DB,4);
TASK_PP(16'hD4DC,4);
TASK_PP(16'hD4DD,4);
TASK_PP(16'hD4DE,4);
TASK_PP(16'hD4DF,4);
TASK_PP(16'hD4E0,4);
TASK_PP(16'hD4E1,4);
TASK_PP(16'hD4E2,4);
TASK_PP(16'hD4E3,4);
TASK_PP(16'hD4E4,4);
TASK_PP(16'hD4E5,4);
TASK_PP(16'hD4E6,4);
TASK_PP(16'hD4E7,4);
TASK_PP(16'hD4E8,4);
TASK_PP(16'hD4E9,4);
TASK_PP(16'hD4EA,4);
TASK_PP(16'hD4EB,4);
TASK_PP(16'hD4EC,4);
TASK_PP(16'hD4ED,4);
TASK_PP(16'hD4EE,4);
TASK_PP(16'hD4EF,4);
TASK_PP(16'hD4F0,4);
TASK_PP(16'hD4F1,4);
TASK_PP(16'hD4F2,4);
TASK_PP(16'hD4F3,4);
TASK_PP(16'hD4F4,4);
TASK_PP(16'hD4F5,4);
TASK_PP(16'hD4F6,4);
TASK_PP(16'hD4F7,4);
TASK_PP(16'hD4F8,4);
TASK_PP(16'hD4F9,4);
TASK_PP(16'hD4FA,4);
TASK_PP(16'hD4FB,4);
TASK_PP(16'hD4FC,4);
TASK_PP(16'hD4FD,4);
TASK_PP(16'hD4FE,4);
TASK_PP(16'hD4FF,4);
TASK_PP(16'hD500,4);
TASK_PP(16'hD501,4);
TASK_PP(16'hD502,4);
TASK_PP(16'hD503,4);
TASK_PP(16'hD504,4);
TASK_PP(16'hD505,4);
TASK_PP(16'hD506,4);
TASK_PP(16'hD507,4);
TASK_PP(16'hD508,4);
TASK_PP(16'hD509,4);
TASK_PP(16'hD50A,4);
TASK_PP(16'hD50B,4);
TASK_PP(16'hD50C,4);
TASK_PP(16'hD50D,4);
TASK_PP(16'hD50E,4);
TASK_PP(16'hD50F,4);
TASK_PP(16'hD510,4);
TASK_PP(16'hD511,4);
TASK_PP(16'hD512,4);
TASK_PP(16'hD513,4);
TASK_PP(16'hD514,4);
TASK_PP(16'hD515,4);
TASK_PP(16'hD516,4);
TASK_PP(16'hD517,4);
TASK_PP(16'hD518,4);
TASK_PP(16'hD519,4);
TASK_PP(16'hD51A,4);
TASK_PP(16'hD51B,4);
TASK_PP(16'hD51C,4);
TASK_PP(16'hD51D,4);
TASK_PP(16'hD51E,4);
TASK_PP(16'hD51F,4);
TASK_PP(16'hD520,4);
TASK_PP(16'hD521,4);
TASK_PP(16'hD522,4);
TASK_PP(16'hD523,4);
TASK_PP(16'hD524,4);
TASK_PP(16'hD525,4);
TASK_PP(16'hD526,4);
TASK_PP(16'hD527,4);
TASK_PP(16'hD528,4);
TASK_PP(16'hD529,4);
TASK_PP(16'hD52A,4);
TASK_PP(16'hD52B,4);
TASK_PP(16'hD52C,4);
TASK_PP(16'hD52D,4);
TASK_PP(16'hD52E,4);
TASK_PP(16'hD52F,4);
TASK_PP(16'hD530,4);
TASK_PP(16'hD531,4);
TASK_PP(16'hD532,4);
TASK_PP(16'hD533,4);
TASK_PP(16'hD534,4);
TASK_PP(16'hD535,4);
TASK_PP(16'hD536,4);
TASK_PP(16'hD537,4);
TASK_PP(16'hD538,4);
TASK_PP(16'hD539,4);
TASK_PP(16'hD53A,4);
TASK_PP(16'hD53B,4);
TASK_PP(16'hD53C,4);
TASK_PP(16'hD53D,4);
TASK_PP(16'hD53E,4);
TASK_PP(16'hD53F,4);
TASK_PP(16'hD540,4);
TASK_PP(16'hD541,4);
TASK_PP(16'hD542,4);
TASK_PP(16'hD543,4);
TASK_PP(16'hD544,4);
TASK_PP(16'hD545,4);
TASK_PP(16'hD546,4);
TASK_PP(16'hD547,4);
TASK_PP(16'hD548,4);
TASK_PP(16'hD549,4);
TASK_PP(16'hD54A,4);
TASK_PP(16'hD54B,4);
TASK_PP(16'hD54C,4);
TASK_PP(16'hD54D,4);
TASK_PP(16'hD54E,4);
TASK_PP(16'hD54F,4);
TASK_PP(16'hD550,4);
TASK_PP(16'hD551,4);
TASK_PP(16'hD552,4);
TASK_PP(16'hD553,4);
TASK_PP(16'hD554,4);
TASK_PP(16'hD555,4);
TASK_PP(16'hD556,4);
TASK_PP(16'hD557,4);
TASK_PP(16'hD558,4);
TASK_PP(16'hD559,4);
TASK_PP(16'hD55A,4);
TASK_PP(16'hD55B,4);
TASK_PP(16'hD55C,4);
TASK_PP(16'hD55D,4);
TASK_PP(16'hD55E,4);
TASK_PP(16'hD55F,4);
TASK_PP(16'hD560,4);
TASK_PP(16'hD561,4);
TASK_PP(16'hD562,4);
TASK_PP(16'hD563,4);
TASK_PP(16'hD564,4);
TASK_PP(16'hD565,4);
TASK_PP(16'hD566,4);
TASK_PP(16'hD567,4);
TASK_PP(16'hD568,4);
TASK_PP(16'hD569,4);
TASK_PP(16'hD56A,4);
TASK_PP(16'hD56B,4);
TASK_PP(16'hD56C,4);
TASK_PP(16'hD56D,4);
TASK_PP(16'hD56E,4);
TASK_PP(16'hD56F,4);
TASK_PP(16'hD570,4);
TASK_PP(16'hD571,4);
TASK_PP(16'hD572,4);
TASK_PP(16'hD573,4);
TASK_PP(16'hD574,4);
TASK_PP(16'hD575,4);
TASK_PP(16'hD576,4);
TASK_PP(16'hD577,4);
TASK_PP(16'hD578,4);
TASK_PP(16'hD579,4);
TASK_PP(16'hD57A,4);
TASK_PP(16'hD57B,4);
TASK_PP(16'hD57C,4);
TASK_PP(16'hD57D,4);
TASK_PP(16'hD57E,4);
TASK_PP(16'hD57F,4);
TASK_PP(16'hD580,4);
TASK_PP(16'hD581,4);
TASK_PP(16'hD582,4);
TASK_PP(16'hD583,4);
TASK_PP(16'hD584,4);
TASK_PP(16'hD585,4);
TASK_PP(16'hD586,4);
TASK_PP(16'hD587,4);
TASK_PP(16'hD588,4);
TASK_PP(16'hD589,4);
TASK_PP(16'hD58A,4);
TASK_PP(16'hD58B,4);
TASK_PP(16'hD58C,4);
TASK_PP(16'hD58D,4);
TASK_PP(16'hD58E,4);
TASK_PP(16'hD58F,4);
TASK_PP(16'hD590,4);
TASK_PP(16'hD591,4);
TASK_PP(16'hD592,4);
TASK_PP(16'hD593,4);
TASK_PP(16'hD594,4);
TASK_PP(16'hD595,4);
TASK_PP(16'hD596,4);
TASK_PP(16'hD597,4);
TASK_PP(16'hD598,4);
TASK_PP(16'hD599,4);
TASK_PP(16'hD59A,4);
TASK_PP(16'hD59B,4);
TASK_PP(16'hD59C,4);
TASK_PP(16'hD59D,4);
TASK_PP(16'hD59E,4);
TASK_PP(16'hD59F,4);
TASK_PP(16'hD5A0,4);
TASK_PP(16'hD5A1,4);
TASK_PP(16'hD5A2,4);
TASK_PP(16'hD5A3,4);
TASK_PP(16'hD5A4,4);
TASK_PP(16'hD5A5,4);
TASK_PP(16'hD5A6,4);
TASK_PP(16'hD5A7,4);
TASK_PP(16'hD5A8,4);
TASK_PP(16'hD5A9,4);
TASK_PP(16'hD5AA,4);
TASK_PP(16'hD5AB,4);
TASK_PP(16'hD5AC,4);
TASK_PP(16'hD5AD,4);
TASK_PP(16'hD5AE,4);
TASK_PP(16'hD5AF,4);
TASK_PP(16'hD5B0,4);
TASK_PP(16'hD5B1,4);
TASK_PP(16'hD5B2,4);
TASK_PP(16'hD5B3,4);
TASK_PP(16'hD5B4,4);
TASK_PP(16'hD5B5,4);
TASK_PP(16'hD5B6,4);
TASK_PP(16'hD5B7,4);
TASK_PP(16'hD5B8,4);
TASK_PP(16'hD5B9,4);
TASK_PP(16'hD5BA,4);
TASK_PP(16'hD5BB,4);
TASK_PP(16'hD5BC,4);
TASK_PP(16'hD5BD,4);
TASK_PP(16'hD5BE,4);
TASK_PP(16'hD5BF,4);
TASK_PP(16'hD5C0,4);
TASK_PP(16'hD5C1,4);
TASK_PP(16'hD5C2,4);
TASK_PP(16'hD5C3,4);
TASK_PP(16'hD5C4,4);
TASK_PP(16'hD5C5,4);
TASK_PP(16'hD5C6,4);
TASK_PP(16'hD5C7,4);
TASK_PP(16'hD5C8,4);
TASK_PP(16'hD5C9,4);
TASK_PP(16'hD5CA,4);
TASK_PP(16'hD5CB,4);
TASK_PP(16'hD5CC,4);
TASK_PP(16'hD5CD,4);
TASK_PP(16'hD5CE,4);
TASK_PP(16'hD5CF,4);
TASK_PP(16'hD5D0,4);
TASK_PP(16'hD5D1,4);
TASK_PP(16'hD5D2,4);
TASK_PP(16'hD5D3,4);
TASK_PP(16'hD5D4,4);
TASK_PP(16'hD5D5,4);
TASK_PP(16'hD5D6,4);
TASK_PP(16'hD5D7,4);
TASK_PP(16'hD5D8,4);
TASK_PP(16'hD5D9,4);
TASK_PP(16'hD5DA,4);
TASK_PP(16'hD5DB,4);
TASK_PP(16'hD5DC,4);
TASK_PP(16'hD5DD,4);
TASK_PP(16'hD5DE,4);
TASK_PP(16'hD5DF,4);
TASK_PP(16'hD5E0,4);
TASK_PP(16'hD5E1,4);
TASK_PP(16'hD5E2,4);
TASK_PP(16'hD5E3,4);
TASK_PP(16'hD5E4,4);
TASK_PP(16'hD5E5,4);
TASK_PP(16'hD5E6,4);
TASK_PP(16'hD5E7,4);
TASK_PP(16'hD5E8,4);
TASK_PP(16'hD5E9,4);
TASK_PP(16'hD5EA,4);
TASK_PP(16'hD5EB,4);
TASK_PP(16'hD5EC,4);
TASK_PP(16'hD5ED,4);
TASK_PP(16'hD5EE,4);
TASK_PP(16'hD5EF,4);
TASK_PP(16'hD5F0,4);
TASK_PP(16'hD5F1,4);
TASK_PP(16'hD5F2,4);
TASK_PP(16'hD5F3,4);
TASK_PP(16'hD5F4,4);
TASK_PP(16'hD5F5,4);
TASK_PP(16'hD5F6,4);
TASK_PP(16'hD5F7,4);
TASK_PP(16'hD5F8,4);
TASK_PP(16'hD5F9,4);
TASK_PP(16'hD5FA,4);
TASK_PP(16'hD5FB,4);
TASK_PP(16'hD5FC,4);
TASK_PP(16'hD5FD,4);
TASK_PP(16'hD5FE,4);
TASK_PP(16'hD5FF,4);
TASK_PP(16'hD600,4);
TASK_PP(16'hD601,4);
TASK_PP(16'hD602,4);
TASK_PP(16'hD603,4);
TASK_PP(16'hD604,4);
TASK_PP(16'hD605,4);
TASK_PP(16'hD606,4);
TASK_PP(16'hD607,4);
TASK_PP(16'hD608,4);
TASK_PP(16'hD609,4);
TASK_PP(16'hD60A,4);
TASK_PP(16'hD60B,4);
TASK_PP(16'hD60C,4);
TASK_PP(16'hD60D,4);
TASK_PP(16'hD60E,4);
TASK_PP(16'hD60F,4);
TASK_PP(16'hD610,4);
TASK_PP(16'hD611,4);
TASK_PP(16'hD612,4);
TASK_PP(16'hD613,4);
TASK_PP(16'hD614,4);
TASK_PP(16'hD615,4);
TASK_PP(16'hD616,4);
TASK_PP(16'hD617,4);
TASK_PP(16'hD618,4);
TASK_PP(16'hD619,4);
TASK_PP(16'hD61A,4);
TASK_PP(16'hD61B,4);
TASK_PP(16'hD61C,4);
TASK_PP(16'hD61D,4);
TASK_PP(16'hD61E,4);
TASK_PP(16'hD61F,4);
TASK_PP(16'hD620,4);
TASK_PP(16'hD621,4);
TASK_PP(16'hD622,4);
TASK_PP(16'hD623,4);
TASK_PP(16'hD624,4);
TASK_PP(16'hD625,4);
TASK_PP(16'hD626,4);
TASK_PP(16'hD627,4);
TASK_PP(16'hD628,4);
TASK_PP(16'hD629,4);
TASK_PP(16'hD62A,4);
TASK_PP(16'hD62B,4);
TASK_PP(16'hD62C,4);
TASK_PP(16'hD62D,4);
TASK_PP(16'hD62E,4);
TASK_PP(16'hD62F,4);
TASK_PP(16'hD630,4);
TASK_PP(16'hD631,4);
TASK_PP(16'hD632,4);
TASK_PP(16'hD633,4);
TASK_PP(16'hD634,4);
TASK_PP(16'hD635,4);
TASK_PP(16'hD636,4);
TASK_PP(16'hD637,4);
TASK_PP(16'hD638,4);
TASK_PP(16'hD639,4);
TASK_PP(16'hD63A,4);
TASK_PP(16'hD63B,4);
TASK_PP(16'hD63C,4);
TASK_PP(16'hD63D,4);
TASK_PP(16'hD63E,4);
TASK_PP(16'hD63F,4);
TASK_PP(16'hD640,4);
TASK_PP(16'hD641,4);
TASK_PP(16'hD642,4);
TASK_PP(16'hD643,4);
TASK_PP(16'hD644,4);
TASK_PP(16'hD645,4);
TASK_PP(16'hD646,4);
TASK_PP(16'hD647,4);
TASK_PP(16'hD648,4);
TASK_PP(16'hD649,4);
TASK_PP(16'hD64A,4);
TASK_PP(16'hD64B,4);
TASK_PP(16'hD64C,4);
TASK_PP(16'hD64D,4);
TASK_PP(16'hD64E,4);
TASK_PP(16'hD64F,4);
TASK_PP(16'hD650,4);
TASK_PP(16'hD651,4);
TASK_PP(16'hD652,4);
TASK_PP(16'hD653,4);
TASK_PP(16'hD654,4);
TASK_PP(16'hD655,4);
TASK_PP(16'hD656,4);
TASK_PP(16'hD657,4);
TASK_PP(16'hD658,4);
TASK_PP(16'hD659,4);
TASK_PP(16'hD65A,4);
TASK_PP(16'hD65B,4);
TASK_PP(16'hD65C,4);
TASK_PP(16'hD65D,4);
TASK_PP(16'hD65E,4);
TASK_PP(16'hD65F,4);
TASK_PP(16'hD660,4);
TASK_PP(16'hD661,4);
TASK_PP(16'hD662,4);
TASK_PP(16'hD663,4);
TASK_PP(16'hD664,4);
TASK_PP(16'hD665,4);
TASK_PP(16'hD666,4);
TASK_PP(16'hD667,4);
TASK_PP(16'hD668,4);
TASK_PP(16'hD669,4);
TASK_PP(16'hD66A,4);
TASK_PP(16'hD66B,4);
TASK_PP(16'hD66C,4);
TASK_PP(16'hD66D,4);
TASK_PP(16'hD66E,4);
TASK_PP(16'hD66F,4);
TASK_PP(16'hD670,4);
TASK_PP(16'hD671,4);
TASK_PP(16'hD672,4);
TASK_PP(16'hD673,4);
TASK_PP(16'hD674,4);
TASK_PP(16'hD675,4);
TASK_PP(16'hD676,4);
TASK_PP(16'hD677,4);
TASK_PP(16'hD678,4);
TASK_PP(16'hD679,4);
TASK_PP(16'hD67A,4);
TASK_PP(16'hD67B,4);
TASK_PP(16'hD67C,4);
TASK_PP(16'hD67D,4);
TASK_PP(16'hD67E,4);
TASK_PP(16'hD67F,4);
TASK_PP(16'hD680,4);
TASK_PP(16'hD681,4);
TASK_PP(16'hD682,4);
TASK_PP(16'hD683,4);
TASK_PP(16'hD684,4);
TASK_PP(16'hD685,4);
TASK_PP(16'hD686,4);
TASK_PP(16'hD687,4);
TASK_PP(16'hD688,4);
TASK_PP(16'hD689,4);
TASK_PP(16'hD68A,4);
TASK_PP(16'hD68B,4);
TASK_PP(16'hD68C,4);
TASK_PP(16'hD68D,4);
TASK_PP(16'hD68E,4);
TASK_PP(16'hD68F,4);
TASK_PP(16'hD690,4);
TASK_PP(16'hD691,4);
TASK_PP(16'hD692,4);
TASK_PP(16'hD693,4);
TASK_PP(16'hD694,4);
TASK_PP(16'hD695,4);
TASK_PP(16'hD696,4);
TASK_PP(16'hD697,4);
TASK_PP(16'hD698,4);
TASK_PP(16'hD699,4);
TASK_PP(16'hD69A,4);
TASK_PP(16'hD69B,4);
TASK_PP(16'hD69C,4);
TASK_PP(16'hD69D,4);
TASK_PP(16'hD69E,4);
TASK_PP(16'hD69F,4);
TASK_PP(16'hD6A0,4);
TASK_PP(16'hD6A1,4);
TASK_PP(16'hD6A2,4);
TASK_PP(16'hD6A3,4);
TASK_PP(16'hD6A4,4);
TASK_PP(16'hD6A5,4);
TASK_PP(16'hD6A6,4);
TASK_PP(16'hD6A7,4);
TASK_PP(16'hD6A8,4);
TASK_PP(16'hD6A9,4);
TASK_PP(16'hD6AA,4);
TASK_PP(16'hD6AB,4);
TASK_PP(16'hD6AC,4);
TASK_PP(16'hD6AD,4);
TASK_PP(16'hD6AE,4);
TASK_PP(16'hD6AF,4);
TASK_PP(16'hD6B0,4);
TASK_PP(16'hD6B1,4);
TASK_PP(16'hD6B2,4);
TASK_PP(16'hD6B3,4);
TASK_PP(16'hD6B4,4);
TASK_PP(16'hD6B5,4);
TASK_PP(16'hD6B6,4);
TASK_PP(16'hD6B7,4);
TASK_PP(16'hD6B8,4);
TASK_PP(16'hD6B9,4);
TASK_PP(16'hD6BA,4);
TASK_PP(16'hD6BB,4);
TASK_PP(16'hD6BC,4);
TASK_PP(16'hD6BD,4);
TASK_PP(16'hD6BE,4);
TASK_PP(16'hD6BF,4);
TASK_PP(16'hD6C0,4);
TASK_PP(16'hD6C1,4);
TASK_PP(16'hD6C2,4);
TASK_PP(16'hD6C3,4);
TASK_PP(16'hD6C4,4);
TASK_PP(16'hD6C5,4);
TASK_PP(16'hD6C6,4);
TASK_PP(16'hD6C7,4);
TASK_PP(16'hD6C8,4);
TASK_PP(16'hD6C9,4);
TASK_PP(16'hD6CA,4);
TASK_PP(16'hD6CB,4);
TASK_PP(16'hD6CC,4);
TASK_PP(16'hD6CD,4);
TASK_PP(16'hD6CE,4);
TASK_PP(16'hD6CF,4);
TASK_PP(16'hD6D0,4);
TASK_PP(16'hD6D1,4);
TASK_PP(16'hD6D2,4);
TASK_PP(16'hD6D3,4);
TASK_PP(16'hD6D4,4);
TASK_PP(16'hD6D5,4);
TASK_PP(16'hD6D6,4);
TASK_PP(16'hD6D7,4);
TASK_PP(16'hD6D8,4);
TASK_PP(16'hD6D9,4);
TASK_PP(16'hD6DA,4);
TASK_PP(16'hD6DB,4);
TASK_PP(16'hD6DC,4);
TASK_PP(16'hD6DD,4);
TASK_PP(16'hD6DE,4);
TASK_PP(16'hD6DF,4);
TASK_PP(16'hD6E0,4);
TASK_PP(16'hD6E1,4);
TASK_PP(16'hD6E2,4);
TASK_PP(16'hD6E3,4);
TASK_PP(16'hD6E4,4);
TASK_PP(16'hD6E5,4);
TASK_PP(16'hD6E6,4);
TASK_PP(16'hD6E7,4);
TASK_PP(16'hD6E8,4);
TASK_PP(16'hD6E9,4);
TASK_PP(16'hD6EA,4);
TASK_PP(16'hD6EB,4);
TASK_PP(16'hD6EC,4);
TASK_PP(16'hD6ED,4);
TASK_PP(16'hD6EE,4);
TASK_PP(16'hD6EF,4);
TASK_PP(16'hD6F0,4);
TASK_PP(16'hD6F1,4);
TASK_PP(16'hD6F2,4);
TASK_PP(16'hD6F3,4);
TASK_PP(16'hD6F4,4);
TASK_PP(16'hD6F5,4);
TASK_PP(16'hD6F6,4);
TASK_PP(16'hD6F7,4);
TASK_PP(16'hD6F8,4);
TASK_PP(16'hD6F9,4);
TASK_PP(16'hD6FA,4);
TASK_PP(16'hD6FB,4);
TASK_PP(16'hD6FC,4);
TASK_PP(16'hD6FD,4);
TASK_PP(16'hD6FE,4);
TASK_PP(16'hD6FF,4);
TASK_PP(16'hD700,4);
TASK_PP(16'hD701,4);
TASK_PP(16'hD702,4);
TASK_PP(16'hD703,4);
TASK_PP(16'hD704,4);
TASK_PP(16'hD705,4);
TASK_PP(16'hD706,4);
TASK_PP(16'hD707,4);
TASK_PP(16'hD708,4);
TASK_PP(16'hD709,4);
TASK_PP(16'hD70A,4);
TASK_PP(16'hD70B,4);
TASK_PP(16'hD70C,4);
TASK_PP(16'hD70D,4);
TASK_PP(16'hD70E,4);
TASK_PP(16'hD70F,4);
TASK_PP(16'hD710,4);
TASK_PP(16'hD711,4);
TASK_PP(16'hD712,4);
TASK_PP(16'hD713,4);
TASK_PP(16'hD714,4);
TASK_PP(16'hD715,4);
TASK_PP(16'hD716,4);
TASK_PP(16'hD717,4);
TASK_PP(16'hD718,4);
TASK_PP(16'hD719,4);
TASK_PP(16'hD71A,4);
TASK_PP(16'hD71B,4);
TASK_PP(16'hD71C,4);
TASK_PP(16'hD71D,4);
TASK_PP(16'hD71E,4);
TASK_PP(16'hD71F,4);
TASK_PP(16'hD720,4);
TASK_PP(16'hD721,4);
TASK_PP(16'hD722,4);
TASK_PP(16'hD723,4);
TASK_PP(16'hD724,4);
TASK_PP(16'hD725,4);
TASK_PP(16'hD726,4);
TASK_PP(16'hD727,4);
TASK_PP(16'hD728,4);
TASK_PP(16'hD729,4);
TASK_PP(16'hD72A,4);
TASK_PP(16'hD72B,4);
TASK_PP(16'hD72C,4);
TASK_PP(16'hD72D,4);
TASK_PP(16'hD72E,4);
TASK_PP(16'hD72F,4);
TASK_PP(16'hD730,4);
TASK_PP(16'hD731,4);
TASK_PP(16'hD732,4);
TASK_PP(16'hD733,4);
TASK_PP(16'hD734,4);
TASK_PP(16'hD735,4);
TASK_PP(16'hD736,4);
TASK_PP(16'hD737,4);
TASK_PP(16'hD738,4);
TASK_PP(16'hD739,4);
TASK_PP(16'hD73A,4);
TASK_PP(16'hD73B,4);
TASK_PP(16'hD73C,4);
TASK_PP(16'hD73D,4);
TASK_PP(16'hD73E,4);
TASK_PP(16'hD73F,4);
TASK_PP(16'hD740,4);
TASK_PP(16'hD741,4);
TASK_PP(16'hD742,4);
TASK_PP(16'hD743,4);
TASK_PP(16'hD744,4);
TASK_PP(16'hD745,4);
TASK_PP(16'hD746,4);
TASK_PP(16'hD747,4);
TASK_PP(16'hD748,4);
TASK_PP(16'hD749,4);
TASK_PP(16'hD74A,4);
TASK_PP(16'hD74B,4);
TASK_PP(16'hD74C,4);
TASK_PP(16'hD74D,4);
TASK_PP(16'hD74E,4);
TASK_PP(16'hD74F,4);
TASK_PP(16'hD750,4);
TASK_PP(16'hD751,4);
TASK_PP(16'hD752,4);
TASK_PP(16'hD753,4);
TASK_PP(16'hD754,4);
TASK_PP(16'hD755,4);
TASK_PP(16'hD756,4);
TASK_PP(16'hD757,4);
TASK_PP(16'hD758,4);
TASK_PP(16'hD759,4);
TASK_PP(16'hD75A,4);
TASK_PP(16'hD75B,4);
TASK_PP(16'hD75C,4);
TASK_PP(16'hD75D,4);
TASK_PP(16'hD75E,4);
TASK_PP(16'hD75F,4);
TASK_PP(16'hD760,4);
TASK_PP(16'hD761,4);
TASK_PP(16'hD762,4);
TASK_PP(16'hD763,4);
TASK_PP(16'hD764,4);
TASK_PP(16'hD765,4);
TASK_PP(16'hD766,4);
TASK_PP(16'hD767,4);
TASK_PP(16'hD768,4);
TASK_PP(16'hD769,4);
TASK_PP(16'hD76A,4);
TASK_PP(16'hD76B,4);
TASK_PP(16'hD76C,4);
TASK_PP(16'hD76D,4);
TASK_PP(16'hD76E,4);
TASK_PP(16'hD76F,4);
TASK_PP(16'hD770,4);
TASK_PP(16'hD771,4);
TASK_PP(16'hD772,4);
TASK_PP(16'hD773,4);
TASK_PP(16'hD774,4);
TASK_PP(16'hD775,4);
TASK_PP(16'hD776,4);
TASK_PP(16'hD777,4);
TASK_PP(16'hD778,4);
TASK_PP(16'hD779,4);
TASK_PP(16'hD77A,4);
TASK_PP(16'hD77B,4);
TASK_PP(16'hD77C,4);
TASK_PP(16'hD77D,4);
TASK_PP(16'hD77E,4);
TASK_PP(16'hD77F,4);
TASK_PP(16'hD780,4);
TASK_PP(16'hD781,4);
TASK_PP(16'hD782,4);
TASK_PP(16'hD783,4);
TASK_PP(16'hD784,4);
TASK_PP(16'hD785,4);
TASK_PP(16'hD786,4);
TASK_PP(16'hD787,4);
TASK_PP(16'hD788,4);
TASK_PP(16'hD789,4);
TASK_PP(16'hD78A,4);
TASK_PP(16'hD78B,4);
TASK_PP(16'hD78C,4);
TASK_PP(16'hD78D,4);
TASK_PP(16'hD78E,4);
TASK_PP(16'hD78F,4);
TASK_PP(16'hD790,4);
TASK_PP(16'hD791,4);
TASK_PP(16'hD792,4);
TASK_PP(16'hD793,4);
TASK_PP(16'hD794,4);
TASK_PP(16'hD795,4);
TASK_PP(16'hD796,4);
TASK_PP(16'hD797,4);
TASK_PP(16'hD798,4);
TASK_PP(16'hD799,4);
TASK_PP(16'hD79A,4);
TASK_PP(16'hD79B,4);
TASK_PP(16'hD79C,4);
TASK_PP(16'hD79D,4);
TASK_PP(16'hD79E,4);
TASK_PP(16'hD79F,4);
TASK_PP(16'hD7A0,4);
TASK_PP(16'hD7A1,4);
TASK_PP(16'hD7A2,4);
TASK_PP(16'hD7A3,4);
TASK_PP(16'hD7A4,4);
TASK_PP(16'hD7A5,4);
TASK_PP(16'hD7A6,4);
TASK_PP(16'hD7A7,4);
TASK_PP(16'hD7A8,4);
TASK_PP(16'hD7A9,4);
TASK_PP(16'hD7AA,4);
TASK_PP(16'hD7AB,4);
TASK_PP(16'hD7AC,4);
TASK_PP(16'hD7AD,4);
TASK_PP(16'hD7AE,4);
TASK_PP(16'hD7AF,4);
TASK_PP(16'hD7B0,4);
TASK_PP(16'hD7B1,4);
TASK_PP(16'hD7B2,4);
TASK_PP(16'hD7B3,4);
TASK_PP(16'hD7B4,4);
TASK_PP(16'hD7B5,4);
TASK_PP(16'hD7B6,4);
TASK_PP(16'hD7B7,4);
TASK_PP(16'hD7B8,4);
TASK_PP(16'hD7B9,4);
TASK_PP(16'hD7BA,4);
TASK_PP(16'hD7BB,4);
TASK_PP(16'hD7BC,4);
TASK_PP(16'hD7BD,4);
TASK_PP(16'hD7BE,4);
TASK_PP(16'hD7BF,4);
TASK_PP(16'hD7C0,4);
TASK_PP(16'hD7C1,4);
TASK_PP(16'hD7C2,4);
TASK_PP(16'hD7C3,4);
TASK_PP(16'hD7C4,4);
TASK_PP(16'hD7C5,4);
TASK_PP(16'hD7C6,4);
TASK_PP(16'hD7C7,4);
TASK_PP(16'hD7C8,4);
TASK_PP(16'hD7C9,4);
TASK_PP(16'hD7CA,4);
TASK_PP(16'hD7CB,4);
TASK_PP(16'hD7CC,4);
TASK_PP(16'hD7CD,4);
TASK_PP(16'hD7CE,4);
TASK_PP(16'hD7CF,4);
TASK_PP(16'hD7D0,4);
TASK_PP(16'hD7D1,4);
TASK_PP(16'hD7D2,4);
TASK_PP(16'hD7D3,4);
TASK_PP(16'hD7D4,4);
TASK_PP(16'hD7D5,4);
TASK_PP(16'hD7D6,4);
TASK_PP(16'hD7D7,4);
TASK_PP(16'hD7D8,4);
TASK_PP(16'hD7D9,4);
TASK_PP(16'hD7DA,4);
TASK_PP(16'hD7DB,4);
TASK_PP(16'hD7DC,4);
TASK_PP(16'hD7DD,4);
TASK_PP(16'hD7DE,4);
TASK_PP(16'hD7DF,4);
TASK_PP(16'hD7E0,4);
TASK_PP(16'hD7E1,4);
TASK_PP(16'hD7E2,4);
TASK_PP(16'hD7E3,4);
TASK_PP(16'hD7E4,4);
TASK_PP(16'hD7E5,4);
TASK_PP(16'hD7E6,4);
TASK_PP(16'hD7E7,4);
TASK_PP(16'hD7E8,4);
TASK_PP(16'hD7E9,4);
TASK_PP(16'hD7EA,4);
TASK_PP(16'hD7EB,4);
TASK_PP(16'hD7EC,4);
TASK_PP(16'hD7ED,4);
TASK_PP(16'hD7EE,4);
TASK_PP(16'hD7EF,4);
TASK_PP(16'hD7F0,4);
TASK_PP(16'hD7F1,4);
TASK_PP(16'hD7F2,4);
TASK_PP(16'hD7F3,4);
TASK_PP(16'hD7F4,4);
TASK_PP(16'hD7F5,4);
TASK_PP(16'hD7F6,4);
TASK_PP(16'hD7F7,4);
TASK_PP(16'hD7F8,4);
TASK_PP(16'hD7F9,4);
TASK_PP(16'hD7FA,4);
TASK_PP(16'hD7FB,4);
TASK_PP(16'hD7FC,4);
TASK_PP(16'hD7FD,4);
TASK_PP(16'hD7FE,4);
TASK_PP(16'hD7FF,4);
TASK_PP(16'hD800,4);
TASK_PP(16'hD801,4);
TASK_PP(16'hD802,4);
TASK_PP(16'hD803,4);
TASK_PP(16'hD804,4);
TASK_PP(16'hD805,4);
TASK_PP(16'hD806,4);
TASK_PP(16'hD807,4);
TASK_PP(16'hD808,4);
TASK_PP(16'hD809,4);
TASK_PP(16'hD80A,4);
TASK_PP(16'hD80B,4);
TASK_PP(16'hD80C,4);
TASK_PP(16'hD80D,4);
TASK_PP(16'hD80E,4);
TASK_PP(16'hD80F,4);
TASK_PP(16'hD810,4);
TASK_PP(16'hD811,4);
TASK_PP(16'hD812,4);
TASK_PP(16'hD813,4);
TASK_PP(16'hD814,4);
TASK_PP(16'hD815,4);
TASK_PP(16'hD816,4);
TASK_PP(16'hD817,4);
TASK_PP(16'hD818,4);
TASK_PP(16'hD819,4);
TASK_PP(16'hD81A,4);
TASK_PP(16'hD81B,4);
TASK_PP(16'hD81C,4);
TASK_PP(16'hD81D,4);
TASK_PP(16'hD81E,4);
TASK_PP(16'hD81F,4);
TASK_PP(16'hD820,4);
TASK_PP(16'hD821,4);
TASK_PP(16'hD822,4);
TASK_PP(16'hD823,4);
TASK_PP(16'hD824,4);
TASK_PP(16'hD825,4);
TASK_PP(16'hD826,4);
TASK_PP(16'hD827,4);
TASK_PP(16'hD828,4);
TASK_PP(16'hD829,4);
TASK_PP(16'hD82A,4);
TASK_PP(16'hD82B,4);
TASK_PP(16'hD82C,4);
TASK_PP(16'hD82D,4);
TASK_PP(16'hD82E,4);
TASK_PP(16'hD82F,4);
TASK_PP(16'hD830,4);
TASK_PP(16'hD831,4);
TASK_PP(16'hD832,4);
TASK_PP(16'hD833,4);
TASK_PP(16'hD834,4);
TASK_PP(16'hD835,4);
TASK_PP(16'hD836,4);
TASK_PP(16'hD837,4);
TASK_PP(16'hD838,4);
TASK_PP(16'hD839,4);
TASK_PP(16'hD83A,4);
TASK_PP(16'hD83B,4);
TASK_PP(16'hD83C,4);
TASK_PP(16'hD83D,4);
TASK_PP(16'hD83E,4);
TASK_PP(16'hD83F,4);
TASK_PP(16'hD840,4);
TASK_PP(16'hD841,4);
TASK_PP(16'hD842,4);
TASK_PP(16'hD843,4);
TASK_PP(16'hD844,4);
TASK_PP(16'hD845,4);
TASK_PP(16'hD846,4);
TASK_PP(16'hD847,4);
TASK_PP(16'hD848,4);
TASK_PP(16'hD849,4);
TASK_PP(16'hD84A,4);
TASK_PP(16'hD84B,4);
TASK_PP(16'hD84C,4);
TASK_PP(16'hD84D,4);
TASK_PP(16'hD84E,4);
TASK_PP(16'hD84F,4);
TASK_PP(16'hD850,4);
TASK_PP(16'hD851,4);
TASK_PP(16'hD852,4);
TASK_PP(16'hD853,4);
TASK_PP(16'hD854,4);
TASK_PP(16'hD855,4);
TASK_PP(16'hD856,4);
TASK_PP(16'hD857,4);
TASK_PP(16'hD858,4);
TASK_PP(16'hD859,4);
TASK_PP(16'hD85A,4);
TASK_PP(16'hD85B,4);
TASK_PP(16'hD85C,4);
TASK_PP(16'hD85D,4);
TASK_PP(16'hD85E,4);
TASK_PP(16'hD85F,4);
TASK_PP(16'hD860,4);
TASK_PP(16'hD861,4);
TASK_PP(16'hD862,4);
TASK_PP(16'hD863,4);
TASK_PP(16'hD864,4);
TASK_PP(16'hD865,4);
TASK_PP(16'hD866,4);
TASK_PP(16'hD867,4);
TASK_PP(16'hD868,4);
TASK_PP(16'hD869,4);
TASK_PP(16'hD86A,4);
TASK_PP(16'hD86B,4);
TASK_PP(16'hD86C,4);
TASK_PP(16'hD86D,4);
TASK_PP(16'hD86E,4);
TASK_PP(16'hD86F,4);
TASK_PP(16'hD870,4);
TASK_PP(16'hD871,4);
TASK_PP(16'hD872,4);
TASK_PP(16'hD873,4);
TASK_PP(16'hD874,4);
TASK_PP(16'hD875,4);
TASK_PP(16'hD876,4);
TASK_PP(16'hD877,4);
TASK_PP(16'hD878,4);
TASK_PP(16'hD879,4);
TASK_PP(16'hD87A,4);
TASK_PP(16'hD87B,4);
TASK_PP(16'hD87C,4);
TASK_PP(16'hD87D,4);
TASK_PP(16'hD87E,4);
TASK_PP(16'hD87F,4);
TASK_PP(16'hD880,4);
TASK_PP(16'hD881,4);
TASK_PP(16'hD882,4);
TASK_PP(16'hD883,4);
TASK_PP(16'hD884,4);
TASK_PP(16'hD885,4);
TASK_PP(16'hD886,4);
TASK_PP(16'hD887,4);
TASK_PP(16'hD888,4);
TASK_PP(16'hD889,4);
TASK_PP(16'hD88A,4);
TASK_PP(16'hD88B,4);
TASK_PP(16'hD88C,4);
TASK_PP(16'hD88D,4);
TASK_PP(16'hD88E,4);
TASK_PP(16'hD88F,4);
TASK_PP(16'hD890,4);
TASK_PP(16'hD891,4);
TASK_PP(16'hD892,4);
TASK_PP(16'hD893,4);
TASK_PP(16'hD894,4);
TASK_PP(16'hD895,4);
TASK_PP(16'hD896,4);
TASK_PP(16'hD897,4);
TASK_PP(16'hD898,4);
TASK_PP(16'hD899,4);
TASK_PP(16'hD89A,4);
TASK_PP(16'hD89B,4);
TASK_PP(16'hD89C,4);
TASK_PP(16'hD89D,4);
TASK_PP(16'hD89E,4);
TASK_PP(16'hD89F,4);
TASK_PP(16'hD8A0,4);
TASK_PP(16'hD8A1,4);
TASK_PP(16'hD8A2,4);
TASK_PP(16'hD8A3,4);
TASK_PP(16'hD8A4,4);
TASK_PP(16'hD8A5,4);
TASK_PP(16'hD8A6,4);
TASK_PP(16'hD8A7,4);
TASK_PP(16'hD8A8,4);
TASK_PP(16'hD8A9,4);
TASK_PP(16'hD8AA,4);
TASK_PP(16'hD8AB,4);
TASK_PP(16'hD8AC,4);
TASK_PP(16'hD8AD,4);
TASK_PP(16'hD8AE,4);
TASK_PP(16'hD8AF,4);
TASK_PP(16'hD8B0,4);
TASK_PP(16'hD8B1,4);
TASK_PP(16'hD8B2,4);
TASK_PP(16'hD8B3,4);
TASK_PP(16'hD8B4,4);
TASK_PP(16'hD8B5,4);
TASK_PP(16'hD8B6,4);
TASK_PP(16'hD8B7,4);
TASK_PP(16'hD8B8,4);
TASK_PP(16'hD8B9,4);
TASK_PP(16'hD8BA,4);
TASK_PP(16'hD8BB,4);
TASK_PP(16'hD8BC,4);
TASK_PP(16'hD8BD,4);
TASK_PP(16'hD8BE,4);
TASK_PP(16'hD8BF,4);
TASK_PP(16'hD8C0,4);
TASK_PP(16'hD8C1,4);
TASK_PP(16'hD8C2,4);
TASK_PP(16'hD8C3,4);
TASK_PP(16'hD8C4,4);
TASK_PP(16'hD8C5,4);
TASK_PP(16'hD8C6,4);
TASK_PP(16'hD8C7,4);
TASK_PP(16'hD8C8,4);
TASK_PP(16'hD8C9,4);
TASK_PP(16'hD8CA,4);
TASK_PP(16'hD8CB,4);
TASK_PP(16'hD8CC,4);
TASK_PP(16'hD8CD,4);
TASK_PP(16'hD8CE,4);
TASK_PP(16'hD8CF,4);
TASK_PP(16'hD8D0,4);
TASK_PP(16'hD8D1,4);
TASK_PP(16'hD8D2,4);
TASK_PP(16'hD8D3,4);
TASK_PP(16'hD8D4,4);
TASK_PP(16'hD8D5,4);
TASK_PP(16'hD8D6,4);
TASK_PP(16'hD8D7,4);
TASK_PP(16'hD8D8,4);
TASK_PP(16'hD8D9,4);
TASK_PP(16'hD8DA,4);
TASK_PP(16'hD8DB,4);
TASK_PP(16'hD8DC,4);
TASK_PP(16'hD8DD,4);
TASK_PP(16'hD8DE,4);
TASK_PP(16'hD8DF,4);
TASK_PP(16'hD8E0,4);
TASK_PP(16'hD8E1,4);
TASK_PP(16'hD8E2,4);
TASK_PP(16'hD8E3,4);
TASK_PP(16'hD8E4,4);
TASK_PP(16'hD8E5,4);
TASK_PP(16'hD8E6,4);
TASK_PP(16'hD8E7,4);
TASK_PP(16'hD8E8,4);
TASK_PP(16'hD8E9,4);
TASK_PP(16'hD8EA,4);
TASK_PP(16'hD8EB,4);
TASK_PP(16'hD8EC,4);
TASK_PP(16'hD8ED,4);
TASK_PP(16'hD8EE,4);
TASK_PP(16'hD8EF,4);
TASK_PP(16'hD8F0,4);
TASK_PP(16'hD8F1,4);
TASK_PP(16'hD8F2,4);
TASK_PP(16'hD8F3,4);
TASK_PP(16'hD8F4,4);
TASK_PP(16'hD8F5,4);
TASK_PP(16'hD8F6,4);
TASK_PP(16'hD8F7,4);
TASK_PP(16'hD8F8,4);
TASK_PP(16'hD8F9,4);
TASK_PP(16'hD8FA,4);
TASK_PP(16'hD8FB,4);
TASK_PP(16'hD8FC,4);
TASK_PP(16'hD8FD,4);
TASK_PP(16'hD8FE,4);
TASK_PP(16'hD8FF,4);
TASK_PP(16'hD900,4);
TASK_PP(16'hD901,4);
TASK_PP(16'hD902,4);
TASK_PP(16'hD903,4);
TASK_PP(16'hD904,4);
TASK_PP(16'hD905,4);
TASK_PP(16'hD906,4);
TASK_PP(16'hD907,4);
TASK_PP(16'hD908,4);
TASK_PP(16'hD909,4);
TASK_PP(16'hD90A,4);
TASK_PP(16'hD90B,4);
TASK_PP(16'hD90C,4);
TASK_PP(16'hD90D,4);
TASK_PP(16'hD90E,4);
TASK_PP(16'hD90F,4);
TASK_PP(16'hD910,4);
TASK_PP(16'hD911,4);
TASK_PP(16'hD912,4);
TASK_PP(16'hD913,4);
TASK_PP(16'hD914,4);
TASK_PP(16'hD915,4);
TASK_PP(16'hD916,4);
TASK_PP(16'hD917,4);
TASK_PP(16'hD918,4);
TASK_PP(16'hD919,4);
TASK_PP(16'hD91A,4);
TASK_PP(16'hD91B,4);
TASK_PP(16'hD91C,4);
TASK_PP(16'hD91D,4);
TASK_PP(16'hD91E,4);
TASK_PP(16'hD91F,4);
TASK_PP(16'hD920,4);
TASK_PP(16'hD921,4);
TASK_PP(16'hD922,4);
TASK_PP(16'hD923,4);
TASK_PP(16'hD924,4);
TASK_PP(16'hD925,4);
TASK_PP(16'hD926,4);
TASK_PP(16'hD927,4);
TASK_PP(16'hD928,4);
TASK_PP(16'hD929,4);
TASK_PP(16'hD92A,4);
TASK_PP(16'hD92B,4);
TASK_PP(16'hD92C,4);
TASK_PP(16'hD92D,4);
TASK_PP(16'hD92E,4);
TASK_PP(16'hD92F,4);
TASK_PP(16'hD930,4);
TASK_PP(16'hD931,4);
TASK_PP(16'hD932,4);
TASK_PP(16'hD933,4);
TASK_PP(16'hD934,4);
TASK_PP(16'hD935,4);
TASK_PP(16'hD936,4);
TASK_PP(16'hD937,4);
TASK_PP(16'hD938,4);
TASK_PP(16'hD939,4);
TASK_PP(16'hD93A,4);
TASK_PP(16'hD93B,4);
TASK_PP(16'hD93C,4);
TASK_PP(16'hD93D,4);
TASK_PP(16'hD93E,4);
TASK_PP(16'hD93F,4);
TASK_PP(16'hD940,4);
TASK_PP(16'hD941,4);
TASK_PP(16'hD942,4);
TASK_PP(16'hD943,4);
TASK_PP(16'hD944,4);
TASK_PP(16'hD945,4);
TASK_PP(16'hD946,4);
TASK_PP(16'hD947,4);
TASK_PP(16'hD948,4);
TASK_PP(16'hD949,4);
TASK_PP(16'hD94A,4);
TASK_PP(16'hD94B,4);
TASK_PP(16'hD94C,4);
TASK_PP(16'hD94D,4);
TASK_PP(16'hD94E,4);
TASK_PP(16'hD94F,4);
TASK_PP(16'hD950,4);
TASK_PP(16'hD951,4);
TASK_PP(16'hD952,4);
TASK_PP(16'hD953,4);
TASK_PP(16'hD954,4);
TASK_PP(16'hD955,4);
TASK_PP(16'hD956,4);
TASK_PP(16'hD957,4);
TASK_PP(16'hD958,4);
TASK_PP(16'hD959,4);
TASK_PP(16'hD95A,4);
TASK_PP(16'hD95B,4);
TASK_PP(16'hD95C,4);
TASK_PP(16'hD95D,4);
TASK_PP(16'hD95E,4);
TASK_PP(16'hD95F,4);
TASK_PP(16'hD960,4);
TASK_PP(16'hD961,4);
TASK_PP(16'hD962,4);
TASK_PP(16'hD963,4);
TASK_PP(16'hD964,4);
TASK_PP(16'hD965,4);
TASK_PP(16'hD966,4);
TASK_PP(16'hD967,4);
TASK_PP(16'hD968,4);
TASK_PP(16'hD969,4);
TASK_PP(16'hD96A,4);
TASK_PP(16'hD96B,4);
TASK_PP(16'hD96C,4);
TASK_PP(16'hD96D,4);
TASK_PP(16'hD96E,4);
TASK_PP(16'hD96F,4);
TASK_PP(16'hD970,4);
TASK_PP(16'hD971,4);
TASK_PP(16'hD972,4);
TASK_PP(16'hD973,4);
TASK_PP(16'hD974,4);
TASK_PP(16'hD975,4);
TASK_PP(16'hD976,4);
TASK_PP(16'hD977,4);
TASK_PP(16'hD978,4);
TASK_PP(16'hD979,4);
TASK_PP(16'hD97A,4);
TASK_PP(16'hD97B,4);
TASK_PP(16'hD97C,4);
TASK_PP(16'hD97D,4);
TASK_PP(16'hD97E,4);
TASK_PP(16'hD97F,4);
TASK_PP(16'hD980,4);
TASK_PP(16'hD981,4);
TASK_PP(16'hD982,4);
TASK_PP(16'hD983,4);
TASK_PP(16'hD984,4);
TASK_PP(16'hD985,4);
TASK_PP(16'hD986,4);
TASK_PP(16'hD987,4);
TASK_PP(16'hD988,4);
TASK_PP(16'hD989,4);
TASK_PP(16'hD98A,4);
TASK_PP(16'hD98B,4);
TASK_PP(16'hD98C,4);
TASK_PP(16'hD98D,4);
TASK_PP(16'hD98E,4);
TASK_PP(16'hD98F,4);
TASK_PP(16'hD990,4);
TASK_PP(16'hD991,4);
TASK_PP(16'hD992,4);
TASK_PP(16'hD993,4);
TASK_PP(16'hD994,4);
TASK_PP(16'hD995,4);
TASK_PP(16'hD996,4);
TASK_PP(16'hD997,4);
TASK_PP(16'hD998,4);
TASK_PP(16'hD999,4);
TASK_PP(16'hD99A,4);
TASK_PP(16'hD99B,4);
TASK_PP(16'hD99C,4);
TASK_PP(16'hD99D,4);
TASK_PP(16'hD99E,4);
TASK_PP(16'hD99F,4);
TASK_PP(16'hD9A0,4);
TASK_PP(16'hD9A1,4);
TASK_PP(16'hD9A2,4);
TASK_PP(16'hD9A3,4);
TASK_PP(16'hD9A4,4);
TASK_PP(16'hD9A5,4);
TASK_PP(16'hD9A6,4);
TASK_PP(16'hD9A7,4);
TASK_PP(16'hD9A8,4);
TASK_PP(16'hD9A9,4);
TASK_PP(16'hD9AA,4);
TASK_PP(16'hD9AB,4);
TASK_PP(16'hD9AC,4);
TASK_PP(16'hD9AD,4);
TASK_PP(16'hD9AE,4);
TASK_PP(16'hD9AF,4);
TASK_PP(16'hD9B0,4);
TASK_PP(16'hD9B1,4);
TASK_PP(16'hD9B2,4);
TASK_PP(16'hD9B3,4);
TASK_PP(16'hD9B4,4);
TASK_PP(16'hD9B5,4);
TASK_PP(16'hD9B6,4);
TASK_PP(16'hD9B7,4);
TASK_PP(16'hD9B8,4);
TASK_PP(16'hD9B9,4);
TASK_PP(16'hD9BA,4);
TASK_PP(16'hD9BB,4);
TASK_PP(16'hD9BC,4);
TASK_PP(16'hD9BD,4);
TASK_PP(16'hD9BE,4);
TASK_PP(16'hD9BF,4);
TASK_PP(16'hD9C0,4);
TASK_PP(16'hD9C1,4);
TASK_PP(16'hD9C2,4);
TASK_PP(16'hD9C3,4);
TASK_PP(16'hD9C4,4);
TASK_PP(16'hD9C5,4);
TASK_PP(16'hD9C6,4);
TASK_PP(16'hD9C7,4);
TASK_PP(16'hD9C8,4);
TASK_PP(16'hD9C9,4);
TASK_PP(16'hD9CA,4);
TASK_PP(16'hD9CB,4);
TASK_PP(16'hD9CC,4);
TASK_PP(16'hD9CD,4);
TASK_PP(16'hD9CE,4);
TASK_PP(16'hD9CF,4);
TASK_PP(16'hD9D0,4);
TASK_PP(16'hD9D1,4);
TASK_PP(16'hD9D2,4);
TASK_PP(16'hD9D3,4);
TASK_PP(16'hD9D4,4);
TASK_PP(16'hD9D5,4);
TASK_PP(16'hD9D6,4);
TASK_PP(16'hD9D7,4);
TASK_PP(16'hD9D8,4);
TASK_PP(16'hD9D9,4);
TASK_PP(16'hD9DA,4);
TASK_PP(16'hD9DB,4);
TASK_PP(16'hD9DC,4);
TASK_PP(16'hD9DD,4);
TASK_PP(16'hD9DE,4);
TASK_PP(16'hD9DF,4);
TASK_PP(16'hD9E0,4);
TASK_PP(16'hD9E1,4);
TASK_PP(16'hD9E2,4);
TASK_PP(16'hD9E3,4);
TASK_PP(16'hD9E4,4);
TASK_PP(16'hD9E5,4);
TASK_PP(16'hD9E6,4);
TASK_PP(16'hD9E7,4);
TASK_PP(16'hD9E8,4);
TASK_PP(16'hD9E9,4);
TASK_PP(16'hD9EA,4);
TASK_PP(16'hD9EB,4);
TASK_PP(16'hD9EC,4);
TASK_PP(16'hD9ED,4);
TASK_PP(16'hD9EE,4);
TASK_PP(16'hD9EF,4);
TASK_PP(16'hD9F0,4);
TASK_PP(16'hD9F1,4);
TASK_PP(16'hD9F2,4);
TASK_PP(16'hD9F3,4);
TASK_PP(16'hD9F4,4);
TASK_PP(16'hD9F5,4);
TASK_PP(16'hD9F6,4);
TASK_PP(16'hD9F7,4);
TASK_PP(16'hD9F8,4);
TASK_PP(16'hD9F9,4);
TASK_PP(16'hD9FA,4);
TASK_PP(16'hD9FB,4);
TASK_PP(16'hD9FC,4);
TASK_PP(16'hD9FD,4);
TASK_PP(16'hD9FE,4);
TASK_PP(16'hD9FF,4);
TASK_PP(16'hDA00,4);
TASK_PP(16'hDA01,4);
TASK_PP(16'hDA02,4);
TASK_PP(16'hDA03,4);
TASK_PP(16'hDA04,4);
TASK_PP(16'hDA05,4);
TASK_PP(16'hDA06,4);
TASK_PP(16'hDA07,4);
TASK_PP(16'hDA08,4);
TASK_PP(16'hDA09,4);
TASK_PP(16'hDA0A,4);
TASK_PP(16'hDA0B,4);
TASK_PP(16'hDA0C,4);
TASK_PP(16'hDA0D,4);
TASK_PP(16'hDA0E,4);
TASK_PP(16'hDA0F,4);
TASK_PP(16'hDA10,4);
TASK_PP(16'hDA11,4);
TASK_PP(16'hDA12,4);
TASK_PP(16'hDA13,4);
TASK_PP(16'hDA14,4);
TASK_PP(16'hDA15,4);
TASK_PP(16'hDA16,4);
TASK_PP(16'hDA17,4);
TASK_PP(16'hDA18,4);
TASK_PP(16'hDA19,4);
TASK_PP(16'hDA1A,4);
TASK_PP(16'hDA1B,4);
TASK_PP(16'hDA1C,4);
TASK_PP(16'hDA1D,4);
TASK_PP(16'hDA1E,4);
TASK_PP(16'hDA1F,4);
TASK_PP(16'hDA20,4);
TASK_PP(16'hDA21,4);
TASK_PP(16'hDA22,4);
TASK_PP(16'hDA23,4);
TASK_PP(16'hDA24,4);
TASK_PP(16'hDA25,4);
TASK_PP(16'hDA26,4);
TASK_PP(16'hDA27,4);
TASK_PP(16'hDA28,4);
TASK_PP(16'hDA29,4);
TASK_PP(16'hDA2A,4);
TASK_PP(16'hDA2B,4);
TASK_PP(16'hDA2C,4);
TASK_PP(16'hDA2D,4);
TASK_PP(16'hDA2E,4);
TASK_PP(16'hDA2F,4);
TASK_PP(16'hDA30,4);
TASK_PP(16'hDA31,4);
TASK_PP(16'hDA32,4);
TASK_PP(16'hDA33,4);
TASK_PP(16'hDA34,4);
TASK_PP(16'hDA35,4);
TASK_PP(16'hDA36,4);
TASK_PP(16'hDA37,4);
TASK_PP(16'hDA38,4);
TASK_PP(16'hDA39,4);
TASK_PP(16'hDA3A,4);
TASK_PP(16'hDA3B,4);
TASK_PP(16'hDA3C,4);
TASK_PP(16'hDA3D,4);
TASK_PP(16'hDA3E,4);
TASK_PP(16'hDA3F,4);
TASK_PP(16'hDA40,4);
TASK_PP(16'hDA41,4);
TASK_PP(16'hDA42,4);
TASK_PP(16'hDA43,4);
TASK_PP(16'hDA44,4);
TASK_PP(16'hDA45,4);
TASK_PP(16'hDA46,4);
TASK_PP(16'hDA47,4);
TASK_PP(16'hDA48,4);
TASK_PP(16'hDA49,4);
TASK_PP(16'hDA4A,4);
TASK_PP(16'hDA4B,4);
TASK_PP(16'hDA4C,4);
TASK_PP(16'hDA4D,4);
TASK_PP(16'hDA4E,4);
TASK_PP(16'hDA4F,4);
TASK_PP(16'hDA50,4);
TASK_PP(16'hDA51,4);
TASK_PP(16'hDA52,4);
TASK_PP(16'hDA53,4);
TASK_PP(16'hDA54,4);
TASK_PP(16'hDA55,4);
TASK_PP(16'hDA56,4);
TASK_PP(16'hDA57,4);
TASK_PP(16'hDA58,4);
TASK_PP(16'hDA59,4);
TASK_PP(16'hDA5A,4);
TASK_PP(16'hDA5B,4);
TASK_PP(16'hDA5C,4);
TASK_PP(16'hDA5D,4);
TASK_PP(16'hDA5E,4);
TASK_PP(16'hDA5F,4);
TASK_PP(16'hDA60,4);
TASK_PP(16'hDA61,4);
TASK_PP(16'hDA62,4);
TASK_PP(16'hDA63,4);
TASK_PP(16'hDA64,4);
TASK_PP(16'hDA65,4);
TASK_PP(16'hDA66,4);
TASK_PP(16'hDA67,4);
TASK_PP(16'hDA68,4);
TASK_PP(16'hDA69,4);
TASK_PP(16'hDA6A,4);
TASK_PP(16'hDA6B,4);
TASK_PP(16'hDA6C,4);
TASK_PP(16'hDA6D,4);
TASK_PP(16'hDA6E,4);
TASK_PP(16'hDA6F,4);
TASK_PP(16'hDA70,4);
TASK_PP(16'hDA71,4);
TASK_PP(16'hDA72,4);
TASK_PP(16'hDA73,4);
TASK_PP(16'hDA74,4);
TASK_PP(16'hDA75,4);
TASK_PP(16'hDA76,4);
TASK_PP(16'hDA77,4);
TASK_PP(16'hDA78,4);
TASK_PP(16'hDA79,4);
TASK_PP(16'hDA7A,4);
TASK_PP(16'hDA7B,4);
TASK_PP(16'hDA7C,4);
TASK_PP(16'hDA7D,4);
TASK_PP(16'hDA7E,4);
TASK_PP(16'hDA7F,4);
TASK_PP(16'hDA80,4);
TASK_PP(16'hDA81,4);
TASK_PP(16'hDA82,4);
TASK_PP(16'hDA83,4);
TASK_PP(16'hDA84,4);
TASK_PP(16'hDA85,4);
TASK_PP(16'hDA86,4);
TASK_PP(16'hDA87,4);
TASK_PP(16'hDA88,4);
TASK_PP(16'hDA89,4);
TASK_PP(16'hDA8A,4);
TASK_PP(16'hDA8B,4);
TASK_PP(16'hDA8C,4);
TASK_PP(16'hDA8D,4);
TASK_PP(16'hDA8E,4);
TASK_PP(16'hDA8F,4);
TASK_PP(16'hDA90,4);
TASK_PP(16'hDA91,4);
TASK_PP(16'hDA92,4);
TASK_PP(16'hDA93,4);
TASK_PP(16'hDA94,4);
TASK_PP(16'hDA95,4);
TASK_PP(16'hDA96,4);
TASK_PP(16'hDA97,4);
TASK_PP(16'hDA98,4);
TASK_PP(16'hDA99,4);
TASK_PP(16'hDA9A,4);
TASK_PP(16'hDA9B,4);
TASK_PP(16'hDA9C,4);
TASK_PP(16'hDA9D,4);
TASK_PP(16'hDA9E,4);
TASK_PP(16'hDA9F,4);
TASK_PP(16'hDAA0,4);
TASK_PP(16'hDAA1,4);
TASK_PP(16'hDAA2,4);
TASK_PP(16'hDAA3,4);
TASK_PP(16'hDAA4,4);
TASK_PP(16'hDAA5,4);
TASK_PP(16'hDAA6,4);
TASK_PP(16'hDAA7,4);
TASK_PP(16'hDAA8,4);
TASK_PP(16'hDAA9,4);
TASK_PP(16'hDAAA,4);
TASK_PP(16'hDAAB,4);
TASK_PP(16'hDAAC,4);
TASK_PP(16'hDAAD,4);
TASK_PP(16'hDAAE,4);
TASK_PP(16'hDAAF,4);
TASK_PP(16'hDAB0,4);
TASK_PP(16'hDAB1,4);
TASK_PP(16'hDAB2,4);
TASK_PP(16'hDAB3,4);
TASK_PP(16'hDAB4,4);
TASK_PP(16'hDAB5,4);
TASK_PP(16'hDAB6,4);
TASK_PP(16'hDAB7,4);
TASK_PP(16'hDAB8,4);
TASK_PP(16'hDAB9,4);
TASK_PP(16'hDABA,4);
TASK_PP(16'hDABB,4);
TASK_PP(16'hDABC,4);
TASK_PP(16'hDABD,4);
TASK_PP(16'hDABE,4);
TASK_PP(16'hDABF,4);
TASK_PP(16'hDAC0,4);
TASK_PP(16'hDAC1,4);
TASK_PP(16'hDAC2,4);
TASK_PP(16'hDAC3,4);
TASK_PP(16'hDAC4,4);
TASK_PP(16'hDAC5,4);
TASK_PP(16'hDAC6,4);
TASK_PP(16'hDAC7,4);
TASK_PP(16'hDAC8,4);
TASK_PP(16'hDAC9,4);
TASK_PP(16'hDACA,4);
TASK_PP(16'hDACB,4);
TASK_PP(16'hDACC,4);
TASK_PP(16'hDACD,4);
TASK_PP(16'hDACE,4);
TASK_PP(16'hDACF,4);
TASK_PP(16'hDAD0,4);
TASK_PP(16'hDAD1,4);
TASK_PP(16'hDAD2,4);
TASK_PP(16'hDAD3,4);
TASK_PP(16'hDAD4,4);
TASK_PP(16'hDAD5,4);
TASK_PP(16'hDAD6,4);
TASK_PP(16'hDAD7,4);
TASK_PP(16'hDAD8,4);
TASK_PP(16'hDAD9,4);
TASK_PP(16'hDADA,4);
TASK_PP(16'hDADB,4);
TASK_PP(16'hDADC,4);
TASK_PP(16'hDADD,4);
TASK_PP(16'hDADE,4);
TASK_PP(16'hDADF,4);
TASK_PP(16'hDAE0,4);
TASK_PP(16'hDAE1,4);
TASK_PP(16'hDAE2,4);
TASK_PP(16'hDAE3,4);
TASK_PP(16'hDAE4,4);
TASK_PP(16'hDAE5,4);
TASK_PP(16'hDAE6,4);
TASK_PP(16'hDAE7,4);
TASK_PP(16'hDAE8,4);
TASK_PP(16'hDAE9,4);
TASK_PP(16'hDAEA,4);
TASK_PP(16'hDAEB,4);
TASK_PP(16'hDAEC,4);
TASK_PP(16'hDAED,4);
TASK_PP(16'hDAEE,4);
TASK_PP(16'hDAEF,4);
TASK_PP(16'hDAF0,4);
TASK_PP(16'hDAF1,4);
TASK_PP(16'hDAF2,4);
TASK_PP(16'hDAF3,4);
TASK_PP(16'hDAF4,4);
TASK_PP(16'hDAF5,4);
TASK_PP(16'hDAF6,4);
TASK_PP(16'hDAF7,4);
TASK_PP(16'hDAF8,4);
TASK_PP(16'hDAF9,4);
TASK_PP(16'hDAFA,4);
TASK_PP(16'hDAFB,4);
TASK_PP(16'hDAFC,4);
TASK_PP(16'hDAFD,4);
TASK_PP(16'hDAFE,4);
TASK_PP(16'hDAFF,4);
TASK_PP(16'hDB00,4);
TASK_PP(16'hDB01,4);
TASK_PP(16'hDB02,4);
TASK_PP(16'hDB03,4);
TASK_PP(16'hDB04,4);
TASK_PP(16'hDB05,4);
TASK_PP(16'hDB06,4);
TASK_PP(16'hDB07,4);
TASK_PP(16'hDB08,4);
TASK_PP(16'hDB09,4);
TASK_PP(16'hDB0A,4);
TASK_PP(16'hDB0B,4);
TASK_PP(16'hDB0C,4);
TASK_PP(16'hDB0D,4);
TASK_PP(16'hDB0E,4);
TASK_PP(16'hDB0F,4);
TASK_PP(16'hDB10,4);
TASK_PP(16'hDB11,4);
TASK_PP(16'hDB12,4);
TASK_PP(16'hDB13,4);
TASK_PP(16'hDB14,4);
TASK_PP(16'hDB15,4);
TASK_PP(16'hDB16,4);
TASK_PP(16'hDB17,4);
TASK_PP(16'hDB18,4);
TASK_PP(16'hDB19,4);
TASK_PP(16'hDB1A,4);
TASK_PP(16'hDB1B,4);
TASK_PP(16'hDB1C,4);
TASK_PP(16'hDB1D,4);
TASK_PP(16'hDB1E,4);
TASK_PP(16'hDB1F,4);
TASK_PP(16'hDB20,4);
TASK_PP(16'hDB21,4);
TASK_PP(16'hDB22,4);
TASK_PP(16'hDB23,4);
TASK_PP(16'hDB24,4);
TASK_PP(16'hDB25,4);
TASK_PP(16'hDB26,4);
TASK_PP(16'hDB27,4);
TASK_PP(16'hDB28,4);
TASK_PP(16'hDB29,4);
TASK_PP(16'hDB2A,4);
TASK_PP(16'hDB2B,4);
TASK_PP(16'hDB2C,4);
TASK_PP(16'hDB2D,4);
TASK_PP(16'hDB2E,4);
TASK_PP(16'hDB2F,4);
TASK_PP(16'hDB30,4);
TASK_PP(16'hDB31,4);
TASK_PP(16'hDB32,4);
TASK_PP(16'hDB33,4);
TASK_PP(16'hDB34,4);
TASK_PP(16'hDB35,4);
TASK_PP(16'hDB36,4);
TASK_PP(16'hDB37,4);
TASK_PP(16'hDB38,4);
TASK_PP(16'hDB39,4);
TASK_PP(16'hDB3A,4);
TASK_PP(16'hDB3B,4);
TASK_PP(16'hDB3C,4);
TASK_PP(16'hDB3D,4);
TASK_PP(16'hDB3E,4);
TASK_PP(16'hDB3F,4);
TASK_PP(16'hDB40,4);
TASK_PP(16'hDB41,4);
TASK_PP(16'hDB42,4);
TASK_PP(16'hDB43,4);
TASK_PP(16'hDB44,4);
TASK_PP(16'hDB45,4);
TASK_PP(16'hDB46,4);
TASK_PP(16'hDB47,4);
TASK_PP(16'hDB48,4);
TASK_PP(16'hDB49,4);
TASK_PP(16'hDB4A,4);
TASK_PP(16'hDB4B,4);
TASK_PP(16'hDB4C,4);
TASK_PP(16'hDB4D,4);
TASK_PP(16'hDB4E,4);
TASK_PP(16'hDB4F,4);
TASK_PP(16'hDB50,4);
TASK_PP(16'hDB51,4);
TASK_PP(16'hDB52,4);
TASK_PP(16'hDB53,4);
TASK_PP(16'hDB54,4);
TASK_PP(16'hDB55,4);
TASK_PP(16'hDB56,4);
TASK_PP(16'hDB57,4);
TASK_PP(16'hDB58,4);
TASK_PP(16'hDB59,4);
TASK_PP(16'hDB5A,4);
TASK_PP(16'hDB5B,4);
TASK_PP(16'hDB5C,4);
TASK_PP(16'hDB5D,4);
TASK_PP(16'hDB5E,4);
TASK_PP(16'hDB5F,4);
TASK_PP(16'hDB60,4);
TASK_PP(16'hDB61,4);
TASK_PP(16'hDB62,4);
TASK_PP(16'hDB63,4);
TASK_PP(16'hDB64,4);
TASK_PP(16'hDB65,4);
TASK_PP(16'hDB66,4);
TASK_PP(16'hDB67,4);
TASK_PP(16'hDB68,4);
TASK_PP(16'hDB69,4);
TASK_PP(16'hDB6A,4);
TASK_PP(16'hDB6B,4);
TASK_PP(16'hDB6C,4);
TASK_PP(16'hDB6D,4);
TASK_PP(16'hDB6E,4);
TASK_PP(16'hDB6F,4);
TASK_PP(16'hDB70,4);
TASK_PP(16'hDB71,4);
TASK_PP(16'hDB72,4);
TASK_PP(16'hDB73,4);
TASK_PP(16'hDB74,4);
TASK_PP(16'hDB75,4);
TASK_PP(16'hDB76,4);
TASK_PP(16'hDB77,4);
TASK_PP(16'hDB78,4);
TASK_PP(16'hDB79,4);
TASK_PP(16'hDB7A,4);
TASK_PP(16'hDB7B,4);
TASK_PP(16'hDB7C,4);
TASK_PP(16'hDB7D,4);
TASK_PP(16'hDB7E,4);
TASK_PP(16'hDB7F,4);
TASK_PP(16'hDB80,4);
TASK_PP(16'hDB81,4);
TASK_PP(16'hDB82,4);
TASK_PP(16'hDB83,4);
TASK_PP(16'hDB84,4);
TASK_PP(16'hDB85,4);
TASK_PP(16'hDB86,4);
TASK_PP(16'hDB87,4);
TASK_PP(16'hDB88,4);
TASK_PP(16'hDB89,4);
TASK_PP(16'hDB8A,4);
TASK_PP(16'hDB8B,4);
TASK_PP(16'hDB8C,4);
TASK_PP(16'hDB8D,4);
TASK_PP(16'hDB8E,4);
TASK_PP(16'hDB8F,4);
TASK_PP(16'hDB90,4);
TASK_PP(16'hDB91,4);
TASK_PP(16'hDB92,4);
TASK_PP(16'hDB93,4);
TASK_PP(16'hDB94,4);
TASK_PP(16'hDB95,4);
TASK_PP(16'hDB96,4);
TASK_PP(16'hDB97,4);
TASK_PP(16'hDB98,4);
TASK_PP(16'hDB99,4);
TASK_PP(16'hDB9A,4);
TASK_PP(16'hDB9B,4);
TASK_PP(16'hDB9C,4);
TASK_PP(16'hDB9D,4);
TASK_PP(16'hDB9E,4);
TASK_PP(16'hDB9F,4);
TASK_PP(16'hDBA0,4);
TASK_PP(16'hDBA1,4);
TASK_PP(16'hDBA2,4);
TASK_PP(16'hDBA3,4);
TASK_PP(16'hDBA4,4);
TASK_PP(16'hDBA5,4);
TASK_PP(16'hDBA6,4);
TASK_PP(16'hDBA7,4);
TASK_PP(16'hDBA8,4);
TASK_PP(16'hDBA9,4);
TASK_PP(16'hDBAA,4);
TASK_PP(16'hDBAB,4);
TASK_PP(16'hDBAC,4);
TASK_PP(16'hDBAD,4);
TASK_PP(16'hDBAE,4);
TASK_PP(16'hDBAF,4);
TASK_PP(16'hDBB0,4);
TASK_PP(16'hDBB1,4);
TASK_PP(16'hDBB2,4);
TASK_PP(16'hDBB3,4);
TASK_PP(16'hDBB4,4);
TASK_PP(16'hDBB5,4);
TASK_PP(16'hDBB6,4);
TASK_PP(16'hDBB7,4);
TASK_PP(16'hDBB8,4);
TASK_PP(16'hDBB9,4);
TASK_PP(16'hDBBA,4);
TASK_PP(16'hDBBB,4);
TASK_PP(16'hDBBC,4);
TASK_PP(16'hDBBD,4);
TASK_PP(16'hDBBE,4);
TASK_PP(16'hDBBF,4);
TASK_PP(16'hDBC0,4);
TASK_PP(16'hDBC1,4);
TASK_PP(16'hDBC2,4);
TASK_PP(16'hDBC3,4);
TASK_PP(16'hDBC4,4);
TASK_PP(16'hDBC5,4);
TASK_PP(16'hDBC6,4);
TASK_PP(16'hDBC7,4);
TASK_PP(16'hDBC8,4);
TASK_PP(16'hDBC9,4);
TASK_PP(16'hDBCA,4);
TASK_PP(16'hDBCB,4);
TASK_PP(16'hDBCC,4);
TASK_PP(16'hDBCD,4);
TASK_PP(16'hDBCE,4);
TASK_PP(16'hDBCF,4);
TASK_PP(16'hDBD0,4);
TASK_PP(16'hDBD1,4);
TASK_PP(16'hDBD2,4);
TASK_PP(16'hDBD3,4);
TASK_PP(16'hDBD4,4);
TASK_PP(16'hDBD5,4);
TASK_PP(16'hDBD6,4);
TASK_PP(16'hDBD7,4);
TASK_PP(16'hDBD8,4);
TASK_PP(16'hDBD9,4);
TASK_PP(16'hDBDA,4);
TASK_PP(16'hDBDB,4);
TASK_PP(16'hDBDC,4);
TASK_PP(16'hDBDD,4);
TASK_PP(16'hDBDE,4);
TASK_PP(16'hDBDF,4);
TASK_PP(16'hDBE0,4);
TASK_PP(16'hDBE1,4);
TASK_PP(16'hDBE2,4);
TASK_PP(16'hDBE3,4);
TASK_PP(16'hDBE4,4);
TASK_PP(16'hDBE5,4);
TASK_PP(16'hDBE6,4);
TASK_PP(16'hDBE7,4);
TASK_PP(16'hDBE8,4);
TASK_PP(16'hDBE9,4);
TASK_PP(16'hDBEA,4);
TASK_PP(16'hDBEB,4);
TASK_PP(16'hDBEC,4);
TASK_PP(16'hDBED,4);
TASK_PP(16'hDBEE,4);
TASK_PP(16'hDBEF,4);
TASK_PP(16'hDBF0,4);
TASK_PP(16'hDBF1,4);
TASK_PP(16'hDBF2,4);
TASK_PP(16'hDBF3,4);
TASK_PP(16'hDBF4,4);
TASK_PP(16'hDBF5,4);
TASK_PP(16'hDBF6,4);
TASK_PP(16'hDBF7,4);
TASK_PP(16'hDBF8,4);
TASK_PP(16'hDBF9,4);
TASK_PP(16'hDBFA,4);
TASK_PP(16'hDBFB,4);
TASK_PP(16'hDBFC,4);
TASK_PP(16'hDBFD,4);
TASK_PP(16'hDBFE,4);
TASK_PP(16'hDBFF,4);
TASK_PP(16'hDC00,4);
TASK_PP(16'hDC01,4);
TASK_PP(16'hDC02,4);
TASK_PP(16'hDC03,4);
TASK_PP(16'hDC04,4);
TASK_PP(16'hDC05,4);
TASK_PP(16'hDC06,4);
TASK_PP(16'hDC07,4);
TASK_PP(16'hDC08,4);
TASK_PP(16'hDC09,4);
TASK_PP(16'hDC0A,4);
TASK_PP(16'hDC0B,4);
TASK_PP(16'hDC0C,4);
TASK_PP(16'hDC0D,4);
TASK_PP(16'hDC0E,4);
TASK_PP(16'hDC0F,4);
TASK_PP(16'hDC10,4);
TASK_PP(16'hDC11,4);
TASK_PP(16'hDC12,4);
TASK_PP(16'hDC13,4);
TASK_PP(16'hDC14,4);
TASK_PP(16'hDC15,4);
TASK_PP(16'hDC16,4);
TASK_PP(16'hDC17,4);
TASK_PP(16'hDC18,4);
TASK_PP(16'hDC19,4);
TASK_PP(16'hDC1A,4);
TASK_PP(16'hDC1B,4);
TASK_PP(16'hDC1C,4);
TASK_PP(16'hDC1D,4);
TASK_PP(16'hDC1E,4);
TASK_PP(16'hDC1F,4);
TASK_PP(16'hDC20,4);
TASK_PP(16'hDC21,4);
TASK_PP(16'hDC22,4);
TASK_PP(16'hDC23,4);
TASK_PP(16'hDC24,4);
TASK_PP(16'hDC25,4);
TASK_PP(16'hDC26,4);
TASK_PP(16'hDC27,4);
TASK_PP(16'hDC28,4);
TASK_PP(16'hDC29,4);
TASK_PP(16'hDC2A,4);
TASK_PP(16'hDC2B,4);
TASK_PP(16'hDC2C,4);
TASK_PP(16'hDC2D,4);
TASK_PP(16'hDC2E,4);
TASK_PP(16'hDC2F,4);
TASK_PP(16'hDC30,4);
TASK_PP(16'hDC31,4);
TASK_PP(16'hDC32,4);
TASK_PP(16'hDC33,4);
TASK_PP(16'hDC34,4);
TASK_PP(16'hDC35,4);
TASK_PP(16'hDC36,4);
TASK_PP(16'hDC37,4);
TASK_PP(16'hDC38,4);
TASK_PP(16'hDC39,4);
TASK_PP(16'hDC3A,4);
TASK_PP(16'hDC3B,4);
TASK_PP(16'hDC3C,4);
TASK_PP(16'hDC3D,4);
TASK_PP(16'hDC3E,4);
TASK_PP(16'hDC3F,4);
TASK_PP(16'hDC40,4);
TASK_PP(16'hDC41,4);
TASK_PP(16'hDC42,4);
TASK_PP(16'hDC43,4);
TASK_PP(16'hDC44,4);
TASK_PP(16'hDC45,4);
TASK_PP(16'hDC46,4);
TASK_PP(16'hDC47,4);
TASK_PP(16'hDC48,4);
TASK_PP(16'hDC49,4);
TASK_PP(16'hDC4A,4);
TASK_PP(16'hDC4B,4);
TASK_PP(16'hDC4C,4);
TASK_PP(16'hDC4D,4);
TASK_PP(16'hDC4E,4);
TASK_PP(16'hDC4F,4);
TASK_PP(16'hDC50,4);
TASK_PP(16'hDC51,4);
TASK_PP(16'hDC52,4);
TASK_PP(16'hDC53,4);
TASK_PP(16'hDC54,4);
TASK_PP(16'hDC55,4);
TASK_PP(16'hDC56,4);
TASK_PP(16'hDC57,4);
TASK_PP(16'hDC58,4);
TASK_PP(16'hDC59,4);
TASK_PP(16'hDC5A,4);
TASK_PP(16'hDC5B,4);
TASK_PP(16'hDC5C,4);
TASK_PP(16'hDC5D,4);
TASK_PP(16'hDC5E,4);
TASK_PP(16'hDC5F,4);
TASK_PP(16'hDC60,4);
TASK_PP(16'hDC61,4);
TASK_PP(16'hDC62,4);
TASK_PP(16'hDC63,4);
TASK_PP(16'hDC64,4);
TASK_PP(16'hDC65,4);
TASK_PP(16'hDC66,4);
TASK_PP(16'hDC67,4);
TASK_PP(16'hDC68,4);
TASK_PP(16'hDC69,4);
TASK_PP(16'hDC6A,4);
TASK_PP(16'hDC6B,4);
TASK_PP(16'hDC6C,4);
TASK_PP(16'hDC6D,4);
TASK_PP(16'hDC6E,4);
TASK_PP(16'hDC6F,4);
TASK_PP(16'hDC70,4);
TASK_PP(16'hDC71,4);
TASK_PP(16'hDC72,4);
TASK_PP(16'hDC73,4);
TASK_PP(16'hDC74,4);
TASK_PP(16'hDC75,4);
TASK_PP(16'hDC76,4);
TASK_PP(16'hDC77,4);
TASK_PP(16'hDC78,4);
TASK_PP(16'hDC79,4);
TASK_PP(16'hDC7A,4);
TASK_PP(16'hDC7B,4);
TASK_PP(16'hDC7C,4);
TASK_PP(16'hDC7D,4);
TASK_PP(16'hDC7E,4);
TASK_PP(16'hDC7F,4);
TASK_PP(16'hDC80,4);
TASK_PP(16'hDC81,4);
TASK_PP(16'hDC82,4);
TASK_PP(16'hDC83,4);
TASK_PP(16'hDC84,4);
TASK_PP(16'hDC85,4);
TASK_PP(16'hDC86,4);
TASK_PP(16'hDC87,4);
TASK_PP(16'hDC88,4);
TASK_PP(16'hDC89,4);
TASK_PP(16'hDC8A,4);
TASK_PP(16'hDC8B,4);
TASK_PP(16'hDC8C,4);
TASK_PP(16'hDC8D,4);
TASK_PP(16'hDC8E,4);
TASK_PP(16'hDC8F,4);
TASK_PP(16'hDC90,4);
TASK_PP(16'hDC91,4);
TASK_PP(16'hDC92,4);
TASK_PP(16'hDC93,4);
TASK_PP(16'hDC94,4);
TASK_PP(16'hDC95,4);
TASK_PP(16'hDC96,4);
TASK_PP(16'hDC97,4);
TASK_PP(16'hDC98,4);
TASK_PP(16'hDC99,4);
TASK_PP(16'hDC9A,4);
TASK_PP(16'hDC9B,4);
TASK_PP(16'hDC9C,4);
TASK_PP(16'hDC9D,4);
TASK_PP(16'hDC9E,4);
TASK_PP(16'hDC9F,4);
TASK_PP(16'hDCA0,4);
TASK_PP(16'hDCA1,4);
TASK_PP(16'hDCA2,4);
TASK_PP(16'hDCA3,4);
TASK_PP(16'hDCA4,4);
TASK_PP(16'hDCA5,4);
TASK_PP(16'hDCA6,4);
TASK_PP(16'hDCA7,4);
TASK_PP(16'hDCA8,4);
TASK_PP(16'hDCA9,4);
TASK_PP(16'hDCAA,4);
TASK_PP(16'hDCAB,4);
TASK_PP(16'hDCAC,4);
TASK_PP(16'hDCAD,4);
TASK_PP(16'hDCAE,4);
TASK_PP(16'hDCAF,4);
TASK_PP(16'hDCB0,4);
TASK_PP(16'hDCB1,4);
TASK_PP(16'hDCB2,4);
TASK_PP(16'hDCB3,4);
TASK_PP(16'hDCB4,4);
TASK_PP(16'hDCB5,4);
TASK_PP(16'hDCB6,4);
TASK_PP(16'hDCB7,4);
TASK_PP(16'hDCB8,4);
TASK_PP(16'hDCB9,4);
TASK_PP(16'hDCBA,4);
TASK_PP(16'hDCBB,4);
TASK_PP(16'hDCBC,4);
TASK_PP(16'hDCBD,4);
TASK_PP(16'hDCBE,4);
TASK_PP(16'hDCBF,4);
TASK_PP(16'hDCC0,4);
TASK_PP(16'hDCC1,4);
TASK_PP(16'hDCC2,4);
TASK_PP(16'hDCC3,4);
TASK_PP(16'hDCC4,4);
TASK_PP(16'hDCC5,4);
TASK_PP(16'hDCC6,4);
TASK_PP(16'hDCC7,4);
TASK_PP(16'hDCC8,4);
TASK_PP(16'hDCC9,4);
TASK_PP(16'hDCCA,4);
TASK_PP(16'hDCCB,4);
TASK_PP(16'hDCCC,4);
TASK_PP(16'hDCCD,4);
TASK_PP(16'hDCCE,4);
TASK_PP(16'hDCCF,4);
TASK_PP(16'hDCD0,4);
TASK_PP(16'hDCD1,4);
TASK_PP(16'hDCD2,4);
TASK_PP(16'hDCD3,4);
TASK_PP(16'hDCD4,4);
TASK_PP(16'hDCD5,4);
TASK_PP(16'hDCD6,4);
TASK_PP(16'hDCD7,4);
TASK_PP(16'hDCD8,4);
TASK_PP(16'hDCD9,4);
TASK_PP(16'hDCDA,4);
TASK_PP(16'hDCDB,4);
TASK_PP(16'hDCDC,4);
TASK_PP(16'hDCDD,4);
TASK_PP(16'hDCDE,4);
TASK_PP(16'hDCDF,4);
TASK_PP(16'hDCE0,4);
TASK_PP(16'hDCE1,4);
TASK_PP(16'hDCE2,4);
TASK_PP(16'hDCE3,4);
TASK_PP(16'hDCE4,4);
TASK_PP(16'hDCE5,4);
TASK_PP(16'hDCE6,4);
TASK_PP(16'hDCE7,4);
TASK_PP(16'hDCE8,4);
TASK_PP(16'hDCE9,4);
TASK_PP(16'hDCEA,4);
TASK_PP(16'hDCEB,4);
TASK_PP(16'hDCEC,4);
TASK_PP(16'hDCED,4);
TASK_PP(16'hDCEE,4);
TASK_PP(16'hDCEF,4);
TASK_PP(16'hDCF0,4);
TASK_PP(16'hDCF1,4);
TASK_PP(16'hDCF2,4);
TASK_PP(16'hDCF3,4);
TASK_PP(16'hDCF4,4);
TASK_PP(16'hDCF5,4);
TASK_PP(16'hDCF6,4);
TASK_PP(16'hDCF7,4);
TASK_PP(16'hDCF8,4);
TASK_PP(16'hDCF9,4);
TASK_PP(16'hDCFA,4);
TASK_PP(16'hDCFB,4);
TASK_PP(16'hDCFC,4);
TASK_PP(16'hDCFD,4);
TASK_PP(16'hDCFE,4);
TASK_PP(16'hDCFF,4);
TASK_PP(16'hDD00,4);
TASK_PP(16'hDD01,4);
TASK_PP(16'hDD02,4);
TASK_PP(16'hDD03,4);
TASK_PP(16'hDD04,4);
TASK_PP(16'hDD05,4);
TASK_PP(16'hDD06,4);
TASK_PP(16'hDD07,4);
TASK_PP(16'hDD08,4);
TASK_PP(16'hDD09,4);
TASK_PP(16'hDD0A,4);
TASK_PP(16'hDD0B,4);
TASK_PP(16'hDD0C,4);
TASK_PP(16'hDD0D,4);
TASK_PP(16'hDD0E,4);
TASK_PP(16'hDD0F,4);
TASK_PP(16'hDD10,4);
TASK_PP(16'hDD11,4);
TASK_PP(16'hDD12,4);
TASK_PP(16'hDD13,4);
TASK_PP(16'hDD14,4);
TASK_PP(16'hDD15,4);
TASK_PP(16'hDD16,4);
TASK_PP(16'hDD17,4);
TASK_PP(16'hDD18,4);
TASK_PP(16'hDD19,4);
TASK_PP(16'hDD1A,4);
TASK_PP(16'hDD1B,4);
TASK_PP(16'hDD1C,4);
TASK_PP(16'hDD1D,4);
TASK_PP(16'hDD1E,4);
TASK_PP(16'hDD1F,4);
TASK_PP(16'hDD20,4);
TASK_PP(16'hDD21,4);
TASK_PP(16'hDD22,4);
TASK_PP(16'hDD23,4);
TASK_PP(16'hDD24,4);
TASK_PP(16'hDD25,4);
TASK_PP(16'hDD26,4);
TASK_PP(16'hDD27,4);
TASK_PP(16'hDD28,4);
TASK_PP(16'hDD29,4);
TASK_PP(16'hDD2A,4);
TASK_PP(16'hDD2B,4);
TASK_PP(16'hDD2C,4);
TASK_PP(16'hDD2D,4);
TASK_PP(16'hDD2E,4);
TASK_PP(16'hDD2F,4);
TASK_PP(16'hDD30,4);
TASK_PP(16'hDD31,4);
TASK_PP(16'hDD32,4);
TASK_PP(16'hDD33,4);
TASK_PP(16'hDD34,4);
TASK_PP(16'hDD35,4);
TASK_PP(16'hDD36,4);
TASK_PP(16'hDD37,4);
TASK_PP(16'hDD38,4);
TASK_PP(16'hDD39,4);
TASK_PP(16'hDD3A,4);
TASK_PP(16'hDD3B,4);
TASK_PP(16'hDD3C,4);
TASK_PP(16'hDD3D,4);
TASK_PP(16'hDD3E,4);
TASK_PP(16'hDD3F,4);
TASK_PP(16'hDD40,4);
TASK_PP(16'hDD41,4);
TASK_PP(16'hDD42,4);
TASK_PP(16'hDD43,4);
TASK_PP(16'hDD44,4);
TASK_PP(16'hDD45,4);
TASK_PP(16'hDD46,4);
TASK_PP(16'hDD47,4);
TASK_PP(16'hDD48,4);
TASK_PP(16'hDD49,4);
TASK_PP(16'hDD4A,4);
TASK_PP(16'hDD4B,4);
TASK_PP(16'hDD4C,4);
TASK_PP(16'hDD4D,4);
TASK_PP(16'hDD4E,4);
TASK_PP(16'hDD4F,4);
TASK_PP(16'hDD50,4);
TASK_PP(16'hDD51,4);
TASK_PP(16'hDD52,4);
TASK_PP(16'hDD53,4);
TASK_PP(16'hDD54,4);
TASK_PP(16'hDD55,4);
TASK_PP(16'hDD56,4);
TASK_PP(16'hDD57,4);
TASK_PP(16'hDD58,4);
TASK_PP(16'hDD59,4);
TASK_PP(16'hDD5A,4);
TASK_PP(16'hDD5B,4);
TASK_PP(16'hDD5C,4);
TASK_PP(16'hDD5D,4);
TASK_PP(16'hDD5E,4);
TASK_PP(16'hDD5F,4);
TASK_PP(16'hDD60,4);
TASK_PP(16'hDD61,4);
TASK_PP(16'hDD62,4);
TASK_PP(16'hDD63,4);
TASK_PP(16'hDD64,4);
TASK_PP(16'hDD65,4);
TASK_PP(16'hDD66,4);
TASK_PP(16'hDD67,4);
TASK_PP(16'hDD68,4);
TASK_PP(16'hDD69,4);
TASK_PP(16'hDD6A,4);
TASK_PP(16'hDD6B,4);
TASK_PP(16'hDD6C,4);
TASK_PP(16'hDD6D,4);
TASK_PP(16'hDD6E,4);
TASK_PP(16'hDD6F,4);
TASK_PP(16'hDD70,4);
TASK_PP(16'hDD71,4);
TASK_PP(16'hDD72,4);
TASK_PP(16'hDD73,4);
TASK_PP(16'hDD74,4);
TASK_PP(16'hDD75,4);
TASK_PP(16'hDD76,4);
TASK_PP(16'hDD77,4);
TASK_PP(16'hDD78,4);
TASK_PP(16'hDD79,4);
TASK_PP(16'hDD7A,4);
TASK_PP(16'hDD7B,4);
TASK_PP(16'hDD7C,4);
TASK_PP(16'hDD7D,4);
TASK_PP(16'hDD7E,4);
TASK_PP(16'hDD7F,4);
TASK_PP(16'hDD80,4);
TASK_PP(16'hDD81,4);
TASK_PP(16'hDD82,4);
TASK_PP(16'hDD83,4);
TASK_PP(16'hDD84,4);
TASK_PP(16'hDD85,4);
TASK_PP(16'hDD86,4);
TASK_PP(16'hDD87,4);
TASK_PP(16'hDD88,4);
TASK_PP(16'hDD89,4);
TASK_PP(16'hDD8A,4);
TASK_PP(16'hDD8B,4);
TASK_PP(16'hDD8C,4);
TASK_PP(16'hDD8D,4);
TASK_PP(16'hDD8E,4);
TASK_PP(16'hDD8F,4);
TASK_PP(16'hDD90,4);
TASK_PP(16'hDD91,4);
TASK_PP(16'hDD92,4);
TASK_PP(16'hDD93,4);
TASK_PP(16'hDD94,4);
TASK_PP(16'hDD95,4);
TASK_PP(16'hDD96,4);
TASK_PP(16'hDD97,4);
TASK_PP(16'hDD98,4);
TASK_PP(16'hDD99,4);
TASK_PP(16'hDD9A,4);
TASK_PP(16'hDD9B,4);
TASK_PP(16'hDD9C,4);
TASK_PP(16'hDD9D,4);
TASK_PP(16'hDD9E,4);
TASK_PP(16'hDD9F,4);
TASK_PP(16'hDDA0,4);
TASK_PP(16'hDDA1,4);
TASK_PP(16'hDDA2,4);
TASK_PP(16'hDDA3,4);
TASK_PP(16'hDDA4,4);
TASK_PP(16'hDDA5,4);
TASK_PP(16'hDDA6,4);
TASK_PP(16'hDDA7,4);
TASK_PP(16'hDDA8,4);
TASK_PP(16'hDDA9,4);
TASK_PP(16'hDDAA,4);
TASK_PP(16'hDDAB,4);
TASK_PP(16'hDDAC,4);
TASK_PP(16'hDDAD,4);
TASK_PP(16'hDDAE,4);
TASK_PP(16'hDDAF,4);
TASK_PP(16'hDDB0,4);
TASK_PP(16'hDDB1,4);
TASK_PP(16'hDDB2,4);
TASK_PP(16'hDDB3,4);
TASK_PP(16'hDDB4,4);
TASK_PP(16'hDDB5,4);
TASK_PP(16'hDDB6,4);
TASK_PP(16'hDDB7,4);
TASK_PP(16'hDDB8,4);
TASK_PP(16'hDDB9,4);
TASK_PP(16'hDDBA,4);
TASK_PP(16'hDDBB,4);
TASK_PP(16'hDDBC,4);
TASK_PP(16'hDDBD,4);
TASK_PP(16'hDDBE,4);
TASK_PP(16'hDDBF,4);
TASK_PP(16'hDDC0,4);
TASK_PP(16'hDDC1,4);
TASK_PP(16'hDDC2,4);
TASK_PP(16'hDDC3,4);
TASK_PP(16'hDDC4,4);
TASK_PP(16'hDDC5,4);
TASK_PP(16'hDDC6,4);
TASK_PP(16'hDDC7,4);
TASK_PP(16'hDDC8,4);
TASK_PP(16'hDDC9,4);
TASK_PP(16'hDDCA,4);
TASK_PP(16'hDDCB,4);
TASK_PP(16'hDDCC,4);
TASK_PP(16'hDDCD,4);
TASK_PP(16'hDDCE,4);
TASK_PP(16'hDDCF,4);
TASK_PP(16'hDDD0,4);
TASK_PP(16'hDDD1,4);
TASK_PP(16'hDDD2,4);
TASK_PP(16'hDDD3,4);
TASK_PP(16'hDDD4,4);
TASK_PP(16'hDDD5,4);
TASK_PP(16'hDDD6,4);
TASK_PP(16'hDDD7,4);
TASK_PP(16'hDDD8,4);
TASK_PP(16'hDDD9,4);
TASK_PP(16'hDDDA,4);
TASK_PP(16'hDDDB,4);
TASK_PP(16'hDDDC,4);
TASK_PP(16'hDDDD,4);
TASK_PP(16'hDDDE,4);
TASK_PP(16'hDDDF,4);
TASK_PP(16'hDDE0,4);
TASK_PP(16'hDDE1,4);
TASK_PP(16'hDDE2,4);
TASK_PP(16'hDDE3,4);
TASK_PP(16'hDDE4,4);
TASK_PP(16'hDDE5,4);
TASK_PP(16'hDDE6,4);
TASK_PP(16'hDDE7,4);
TASK_PP(16'hDDE8,4);
TASK_PP(16'hDDE9,4);
TASK_PP(16'hDDEA,4);
TASK_PP(16'hDDEB,4);
TASK_PP(16'hDDEC,4);
TASK_PP(16'hDDED,4);
TASK_PP(16'hDDEE,4);
TASK_PP(16'hDDEF,4);
TASK_PP(16'hDDF0,4);
TASK_PP(16'hDDF1,4);
TASK_PP(16'hDDF2,4);
TASK_PP(16'hDDF3,4);
TASK_PP(16'hDDF4,4);
TASK_PP(16'hDDF5,4);
TASK_PP(16'hDDF6,4);
TASK_PP(16'hDDF7,4);
TASK_PP(16'hDDF8,4);
TASK_PP(16'hDDF9,4);
TASK_PP(16'hDDFA,4);
TASK_PP(16'hDDFB,4);
TASK_PP(16'hDDFC,4);
TASK_PP(16'hDDFD,4);
TASK_PP(16'hDDFE,4);
TASK_PP(16'hDDFF,4);
TASK_PP(16'hDE00,4);
TASK_PP(16'hDE01,4);
TASK_PP(16'hDE02,4);
TASK_PP(16'hDE03,4);
TASK_PP(16'hDE04,4);
TASK_PP(16'hDE05,4);
TASK_PP(16'hDE06,4);
TASK_PP(16'hDE07,4);
TASK_PP(16'hDE08,4);
TASK_PP(16'hDE09,4);
TASK_PP(16'hDE0A,4);
TASK_PP(16'hDE0B,4);
TASK_PP(16'hDE0C,4);
TASK_PP(16'hDE0D,4);
TASK_PP(16'hDE0E,4);
TASK_PP(16'hDE0F,4);
TASK_PP(16'hDE10,4);
TASK_PP(16'hDE11,4);
TASK_PP(16'hDE12,4);
TASK_PP(16'hDE13,4);
TASK_PP(16'hDE14,4);
TASK_PP(16'hDE15,4);
TASK_PP(16'hDE16,4);
TASK_PP(16'hDE17,4);
TASK_PP(16'hDE18,4);
TASK_PP(16'hDE19,4);
TASK_PP(16'hDE1A,4);
TASK_PP(16'hDE1B,4);
TASK_PP(16'hDE1C,4);
TASK_PP(16'hDE1D,4);
TASK_PP(16'hDE1E,4);
TASK_PP(16'hDE1F,4);
TASK_PP(16'hDE20,4);
TASK_PP(16'hDE21,4);
TASK_PP(16'hDE22,4);
TASK_PP(16'hDE23,4);
TASK_PP(16'hDE24,4);
TASK_PP(16'hDE25,4);
TASK_PP(16'hDE26,4);
TASK_PP(16'hDE27,4);
TASK_PP(16'hDE28,4);
TASK_PP(16'hDE29,4);
TASK_PP(16'hDE2A,4);
TASK_PP(16'hDE2B,4);
TASK_PP(16'hDE2C,4);
TASK_PP(16'hDE2D,4);
TASK_PP(16'hDE2E,4);
TASK_PP(16'hDE2F,4);
TASK_PP(16'hDE30,4);
TASK_PP(16'hDE31,4);
TASK_PP(16'hDE32,4);
TASK_PP(16'hDE33,4);
TASK_PP(16'hDE34,4);
TASK_PP(16'hDE35,4);
TASK_PP(16'hDE36,4);
TASK_PP(16'hDE37,4);
TASK_PP(16'hDE38,4);
TASK_PP(16'hDE39,4);
TASK_PP(16'hDE3A,4);
TASK_PP(16'hDE3B,4);
TASK_PP(16'hDE3C,4);
TASK_PP(16'hDE3D,4);
TASK_PP(16'hDE3E,4);
TASK_PP(16'hDE3F,4);
TASK_PP(16'hDE40,4);
TASK_PP(16'hDE41,4);
TASK_PP(16'hDE42,4);
TASK_PP(16'hDE43,4);
TASK_PP(16'hDE44,4);
TASK_PP(16'hDE45,4);
TASK_PP(16'hDE46,4);
TASK_PP(16'hDE47,4);
TASK_PP(16'hDE48,4);
TASK_PP(16'hDE49,4);
TASK_PP(16'hDE4A,4);
TASK_PP(16'hDE4B,4);
TASK_PP(16'hDE4C,4);
TASK_PP(16'hDE4D,4);
TASK_PP(16'hDE4E,4);
TASK_PP(16'hDE4F,4);
TASK_PP(16'hDE50,4);
TASK_PP(16'hDE51,4);
TASK_PP(16'hDE52,4);
TASK_PP(16'hDE53,4);
TASK_PP(16'hDE54,4);
TASK_PP(16'hDE55,4);
TASK_PP(16'hDE56,4);
TASK_PP(16'hDE57,4);
TASK_PP(16'hDE58,4);
TASK_PP(16'hDE59,4);
TASK_PP(16'hDE5A,4);
TASK_PP(16'hDE5B,4);
TASK_PP(16'hDE5C,4);
TASK_PP(16'hDE5D,4);
TASK_PP(16'hDE5E,4);
TASK_PP(16'hDE5F,4);
TASK_PP(16'hDE60,4);
TASK_PP(16'hDE61,4);
TASK_PP(16'hDE62,4);
TASK_PP(16'hDE63,4);
TASK_PP(16'hDE64,4);
TASK_PP(16'hDE65,4);
TASK_PP(16'hDE66,4);
TASK_PP(16'hDE67,4);
TASK_PP(16'hDE68,4);
TASK_PP(16'hDE69,4);
TASK_PP(16'hDE6A,4);
TASK_PP(16'hDE6B,4);
TASK_PP(16'hDE6C,4);
TASK_PP(16'hDE6D,4);
TASK_PP(16'hDE6E,4);
TASK_PP(16'hDE6F,4);
TASK_PP(16'hDE70,4);
TASK_PP(16'hDE71,4);
TASK_PP(16'hDE72,4);
TASK_PP(16'hDE73,4);
TASK_PP(16'hDE74,4);
TASK_PP(16'hDE75,4);
TASK_PP(16'hDE76,4);
TASK_PP(16'hDE77,4);
TASK_PP(16'hDE78,4);
TASK_PP(16'hDE79,4);
TASK_PP(16'hDE7A,4);
TASK_PP(16'hDE7B,4);
TASK_PP(16'hDE7C,4);
TASK_PP(16'hDE7D,4);
TASK_PP(16'hDE7E,4);
TASK_PP(16'hDE7F,4);
TASK_PP(16'hDE80,4);
TASK_PP(16'hDE81,4);
TASK_PP(16'hDE82,4);
TASK_PP(16'hDE83,4);
TASK_PP(16'hDE84,4);
TASK_PP(16'hDE85,4);
TASK_PP(16'hDE86,4);
TASK_PP(16'hDE87,4);
TASK_PP(16'hDE88,4);
TASK_PP(16'hDE89,4);
TASK_PP(16'hDE8A,4);
TASK_PP(16'hDE8B,4);
TASK_PP(16'hDE8C,4);
TASK_PP(16'hDE8D,4);
TASK_PP(16'hDE8E,4);
TASK_PP(16'hDE8F,4);
TASK_PP(16'hDE90,4);
TASK_PP(16'hDE91,4);
TASK_PP(16'hDE92,4);
TASK_PP(16'hDE93,4);
TASK_PP(16'hDE94,4);
TASK_PP(16'hDE95,4);
TASK_PP(16'hDE96,4);
TASK_PP(16'hDE97,4);
TASK_PP(16'hDE98,4);
TASK_PP(16'hDE99,4);
TASK_PP(16'hDE9A,4);
TASK_PP(16'hDE9B,4);
TASK_PP(16'hDE9C,4);
TASK_PP(16'hDE9D,4);
TASK_PP(16'hDE9E,4);
TASK_PP(16'hDE9F,4);
TASK_PP(16'hDEA0,4);
TASK_PP(16'hDEA1,4);
TASK_PP(16'hDEA2,4);
TASK_PP(16'hDEA3,4);
TASK_PP(16'hDEA4,4);
TASK_PP(16'hDEA5,4);
TASK_PP(16'hDEA6,4);
TASK_PP(16'hDEA7,4);
TASK_PP(16'hDEA8,4);
TASK_PP(16'hDEA9,4);
TASK_PP(16'hDEAA,4);
TASK_PP(16'hDEAB,4);
TASK_PP(16'hDEAC,4);
TASK_PP(16'hDEAD,4);
TASK_PP(16'hDEAE,4);
TASK_PP(16'hDEAF,4);
TASK_PP(16'hDEB0,4);
TASK_PP(16'hDEB1,4);
TASK_PP(16'hDEB2,4);
TASK_PP(16'hDEB3,4);
TASK_PP(16'hDEB4,4);
TASK_PP(16'hDEB5,4);
TASK_PP(16'hDEB6,4);
TASK_PP(16'hDEB7,4);
TASK_PP(16'hDEB8,4);
TASK_PP(16'hDEB9,4);
TASK_PP(16'hDEBA,4);
TASK_PP(16'hDEBB,4);
TASK_PP(16'hDEBC,4);
TASK_PP(16'hDEBD,4);
TASK_PP(16'hDEBE,4);
TASK_PP(16'hDEBF,4);
TASK_PP(16'hDEC0,4);
TASK_PP(16'hDEC1,4);
TASK_PP(16'hDEC2,4);
TASK_PP(16'hDEC3,4);
TASK_PP(16'hDEC4,4);
TASK_PP(16'hDEC5,4);
TASK_PP(16'hDEC6,4);
TASK_PP(16'hDEC7,4);
TASK_PP(16'hDEC8,4);
TASK_PP(16'hDEC9,4);
TASK_PP(16'hDECA,4);
TASK_PP(16'hDECB,4);
TASK_PP(16'hDECC,4);
TASK_PP(16'hDECD,4);
TASK_PP(16'hDECE,4);
TASK_PP(16'hDECF,4);
TASK_PP(16'hDED0,4);
TASK_PP(16'hDED1,4);
TASK_PP(16'hDED2,4);
TASK_PP(16'hDED3,4);
TASK_PP(16'hDED4,4);
TASK_PP(16'hDED5,4);
TASK_PP(16'hDED6,4);
TASK_PP(16'hDED7,4);
TASK_PP(16'hDED8,4);
TASK_PP(16'hDED9,4);
TASK_PP(16'hDEDA,4);
TASK_PP(16'hDEDB,4);
TASK_PP(16'hDEDC,4);
TASK_PP(16'hDEDD,4);
TASK_PP(16'hDEDE,4);
TASK_PP(16'hDEDF,4);
TASK_PP(16'hDEE0,4);
TASK_PP(16'hDEE1,4);
TASK_PP(16'hDEE2,4);
TASK_PP(16'hDEE3,4);
TASK_PP(16'hDEE4,4);
TASK_PP(16'hDEE5,4);
TASK_PP(16'hDEE6,4);
TASK_PP(16'hDEE7,4);
TASK_PP(16'hDEE8,4);
TASK_PP(16'hDEE9,4);
TASK_PP(16'hDEEA,4);
TASK_PP(16'hDEEB,4);
TASK_PP(16'hDEEC,4);
TASK_PP(16'hDEED,4);
TASK_PP(16'hDEEE,4);
TASK_PP(16'hDEEF,4);
TASK_PP(16'hDEF0,4);
TASK_PP(16'hDEF1,4);
TASK_PP(16'hDEF2,4);
TASK_PP(16'hDEF3,4);
TASK_PP(16'hDEF4,4);
TASK_PP(16'hDEF5,4);
TASK_PP(16'hDEF6,4);
TASK_PP(16'hDEF7,4);
TASK_PP(16'hDEF8,4);
TASK_PP(16'hDEF9,4);
TASK_PP(16'hDEFA,4);
TASK_PP(16'hDEFB,4);
TASK_PP(16'hDEFC,4);
TASK_PP(16'hDEFD,4);
TASK_PP(16'hDEFE,4);
TASK_PP(16'hDEFF,4);
TASK_PP(16'hDF00,4);
TASK_PP(16'hDF01,4);
TASK_PP(16'hDF02,4);
TASK_PP(16'hDF03,4);
TASK_PP(16'hDF04,4);
TASK_PP(16'hDF05,4);
TASK_PP(16'hDF06,4);
TASK_PP(16'hDF07,4);
TASK_PP(16'hDF08,4);
TASK_PP(16'hDF09,4);
TASK_PP(16'hDF0A,4);
TASK_PP(16'hDF0B,4);
TASK_PP(16'hDF0C,4);
TASK_PP(16'hDF0D,4);
TASK_PP(16'hDF0E,4);
TASK_PP(16'hDF0F,4);
TASK_PP(16'hDF10,4);
TASK_PP(16'hDF11,4);
TASK_PP(16'hDF12,4);
TASK_PP(16'hDF13,4);
TASK_PP(16'hDF14,4);
TASK_PP(16'hDF15,4);
TASK_PP(16'hDF16,4);
TASK_PP(16'hDF17,4);
TASK_PP(16'hDF18,4);
TASK_PP(16'hDF19,4);
TASK_PP(16'hDF1A,4);
TASK_PP(16'hDF1B,4);
TASK_PP(16'hDF1C,4);
TASK_PP(16'hDF1D,4);
TASK_PP(16'hDF1E,4);
TASK_PP(16'hDF1F,4);
TASK_PP(16'hDF20,4);
TASK_PP(16'hDF21,4);
TASK_PP(16'hDF22,4);
TASK_PP(16'hDF23,4);
TASK_PP(16'hDF24,4);
TASK_PP(16'hDF25,4);
TASK_PP(16'hDF26,4);
TASK_PP(16'hDF27,4);
TASK_PP(16'hDF28,4);
TASK_PP(16'hDF29,4);
TASK_PP(16'hDF2A,4);
TASK_PP(16'hDF2B,4);
TASK_PP(16'hDF2C,4);
TASK_PP(16'hDF2D,4);
TASK_PP(16'hDF2E,4);
TASK_PP(16'hDF2F,4);
TASK_PP(16'hDF30,4);
TASK_PP(16'hDF31,4);
TASK_PP(16'hDF32,4);
TASK_PP(16'hDF33,4);
TASK_PP(16'hDF34,4);
TASK_PP(16'hDF35,4);
TASK_PP(16'hDF36,4);
TASK_PP(16'hDF37,4);
TASK_PP(16'hDF38,4);
TASK_PP(16'hDF39,4);
TASK_PP(16'hDF3A,4);
TASK_PP(16'hDF3B,4);
TASK_PP(16'hDF3C,4);
TASK_PP(16'hDF3D,4);
TASK_PP(16'hDF3E,4);
TASK_PP(16'hDF3F,4);
TASK_PP(16'hDF40,4);
TASK_PP(16'hDF41,4);
TASK_PP(16'hDF42,4);
TASK_PP(16'hDF43,4);
TASK_PP(16'hDF44,4);
TASK_PP(16'hDF45,4);
TASK_PP(16'hDF46,4);
TASK_PP(16'hDF47,4);
TASK_PP(16'hDF48,4);
TASK_PP(16'hDF49,4);
TASK_PP(16'hDF4A,4);
TASK_PP(16'hDF4B,4);
TASK_PP(16'hDF4C,4);
TASK_PP(16'hDF4D,4);
TASK_PP(16'hDF4E,4);
TASK_PP(16'hDF4F,4);
TASK_PP(16'hDF50,4);
TASK_PP(16'hDF51,4);
TASK_PP(16'hDF52,4);
TASK_PP(16'hDF53,4);
TASK_PP(16'hDF54,4);
TASK_PP(16'hDF55,4);
TASK_PP(16'hDF56,4);
TASK_PP(16'hDF57,4);
TASK_PP(16'hDF58,4);
TASK_PP(16'hDF59,4);
TASK_PP(16'hDF5A,4);
TASK_PP(16'hDF5B,4);
TASK_PP(16'hDF5C,4);
TASK_PP(16'hDF5D,4);
TASK_PP(16'hDF5E,4);
TASK_PP(16'hDF5F,4);
TASK_PP(16'hDF60,4);
TASK_PP(16'hDF61,4);
TASK_PP(16'hDF62,4);
TASK_PP(16'hDF63,4);
TASK_PP(16'hDF64,4);
TASK_PP(16'hDF65,4);
TASK_PP(16'hDF66,4);
TASK_PP(16'hDF67,4);
TASK_PP(16'hDF68,4);
TASK_PP(16'hDF69,4);
TASK_PP(16'hDF6A,4);
TASK_PP(16'hDF6B,4);
TASK_PP(16'hDF6C,4);
TASK_PP(16'hDF6D,4);
TASK_PP(16'hDF6E,4);
TASK_PP(16'hDF6F,4);
TASK_PP(16'hDF70,4);
TASK_PP(16'hDF71,4);
TASK_PP(16'hDF72,4);
TASK_PP(16'hDF73,4);
TASK_PP(16'hDF74,4);
TASK_PP(16'hDF75,4);
TASK_PP(16'hDF76,4);
TASK_PP(16'hDF77,4);
TASK_PP(16'hDF78,4);
TASK_PP(16'hDF79,4);
TASK_PP(16'hDF7A,4);
TASK_PP(16'hDF7B,4);
TASK_PP(16'hDF7C,4);
TASK_PP(16'hDF7D,4);
TASK_PP(16'hDF7E,4);
TASK_PP(16'hDF7F,4);
TASK_PP(16'hDF80,4);
TASK_PP(16'hDF81,4);
TASK_PP(16'hDF82,4);
TASK_PP(16'hDF83,4);
TASK_PP(16'hDF84,4);
TASK_PP(16'hDF85,4);
TASK_PP(16'hDF86,4);
TASK_PP(16'hDF87,4);
TASK_PP(16'hDF88,4);
TASK_PP(16'hDF89,4);
TASK_PP(16'hDF8A,4);
TASK_PP(16'hDF8B,4);
TASK_PP(16'hDF8C,4);
TASK_PP(16'hDF8D,4);
TASK_PP(16'hDF8E,4);
TASK_PP(16'hDF8F,4);
TASK_PP(16'hDF90,4);
TASK_PP(16'hDF91,4);
TASK_PP(16'hDF92,4);
TASK_PP(16'hDF93,4);
TASK_PP(16'hDF94,4);
TASK_PP(16'hDF95,4);
TASK_PP(16'hDF96,4);
TASK_PP(16'hDF97,4);
TASK_PP(16'hDF98,4);
TASK_PP(16'hDF99,4);
TASK_PP(16'hDF9A,4);
TASK_PP(16'hDF9B,4);
TASK_PP(16'hDF9C,4);
TASK_PP(16'hDF9D,4);
TASK_PP(16'hDF9E,4);
TASK_PP(16'hDF9F,4);
TASK_PP(16'hDFA0,4);
TASK_PP(16'hDFA1,4);
TASK_PP(16'hDFA2,4);
TASK_PP(16'hDFA3,4);
TASK_PP(16'hDFA4,4);
TASK_PP(16'hDFA5,4);
TASK_PP(16'hDFA6,4);
TASK_PP(16'hDFA7,4);
TASK_PP(16'hDFA8,4);
TASK_PP(16'hDFA9,4);
TASK_PP(16'hDFAA,4);
TASK_PP(16'hDFAB,4);
TASK_PP(16'hDFAC,4);
TASK_PP(16'hDFAD,4);
TASK_PP(16'hDFAE,4);
TASK_PP(16'hDFAF,4);
TASK_PP(16'hDFB0,4);
TASK_PP(16'hDFB1,4);
TASK_PP(16'hDFB2,4);
TASK_PP(16'hDFB3,4);
TASK_PP(16'hDFB4,4);
TASK_PP(16'hDFB5,4);
TASK_PP(16'hDFB6,4);
TASK_PP(16'hDFB7,4);
TASK_PP(16'hDFB8,4);
TASK_PP(16'hDFB9,4);
TASK_PP(16'hDFBA,4);
TASK_PP(16'hDFBB,4);
TASK_PP(16'hDFBC,4);
TASK_PP(16'hDFBD,4);
TASK_PP(16'hDFBE,4);
TASK_PP(16'hDFBF,4);
TASK_PP(16'hDFC0,4);
TASK_PP(16'hDFC1,4);
TASK_PP(16'hDFC2,4);
TASK_PP(16'hDFC3,4);
TASK_PP(16'hDFC4,4);
TASK_PP(16'hDFC5,4);
TASK_PP(16'hDFC6,4);
TASK_PP(16'hDFC7,4);
TASK_PP(16'hDFC8,4);
TASK_PP(16'hDFC9,4);
TASK_PP(16'hDFCA,4);
TASK_PP(16'hDFCB,4);
TASK_PP(16'hDFCC,4);
TASK_PP(16'hDFCD,4);
TASK_PP(16'hDFCE,4);
TASK_PP(16'hDFCF,4);
TASK_PP(16'hDFD0,4);
TASK_PP(16'hDFD1,4);
TASK_PP(16'hDFD2,4);
TASK_PP(16'hDFD3,4);
TASK_PP(16'hDFD4,4);
TASK_PP(16'hDFD5,4);
TASK_PP(16'hDFD6,4);
TASK_PP(16'hDFD7,4);
TASK_PP(16'hDFD8,4);
TASK_PP(16'hDFD9,4);
TASK_PP(16'hDFDA,4);
TASK_PP(16'hDFDB,4);
TASK_PP(16'hDFDC,4);
TASK_PP(16'hDFDD,4);
TASK_PP(16'hDFDE,4);
TASK_PP(16'hDFDF,4);
TASK_PP(16'hDFE0,4);
TASK_PP(16'hDFE1,4);
TASK_PP(16'hDFE2,4);
TASK_PP(16'hDFE3,4);
TASK_PP(16'hDFE4,4);
TASK_PP(16'hDFE5,4);
TASK_PP(16'hDFE6,4);
TASK_PP(16'hDFE7,4);
TASK_PP(16'hDFE8,4);
TASK_PP(16'hDFE9,4);
TASK_PP(16'hDFEA,4);
TASK_PP(16'hDFEB,4);
TASK_PP(16'hDFEC,4);
TASK_PP(16'hDFED,4);
TASK_PP(16'hDFEE,4);
TASK_PP(16'hDFEF,4);
TASK_PP(16'hDFF0,4);
TASK_PP(16'hDFF1,4);
TASK_PP(16'hDFF2,4);
TASK_PP(16'hDFF3,4);
TASK_PP(16'hDFF4,4);
TASK_PP(16'hDFF5,4);
TASK_PP(16'hDFF6,4);
TASK_PP(16'hDFF7,4);
TASK_PP(16'hDFF8,4);
TASK_PP(16'hDFF9,4);
TASK_PP(16'hDFFA,4);
TASK_PP(16'hDFFB,4);
TASK_PP(16'hDFFC,4);
TASK_PP(16'hDFFD,4);
TASK_PP(16'hDFFE,4);
TASK_PP(16'hDFFF,4);
TASK_PP(16'hE000,4);
TASK_PP(16'hE001,4);
TASK_PP(16'hE002,4);
TASK_PP(16'hE003,4);
TASK_PP(16'hE004,4);
TASK_PP(16'hE005,4);
TASK_PP(16'hE006,4);
TASK_PP(16'hE007,4);
TASK_PP(16'hE008,4);
TASK_PP(16'hE009,4);
TASK_PP(16'hE00A,4);
TASK_PP(16'hE00B,4);
TASK_PP(16'hE00C,4);
TASK_PP(16'hE00D,4);
TASK_PP(16'hE00E,4);
TASK_PP(16'hE00F,4);
TASK_PP(16'hE010,4);
TASK_PP(16'hE011,4);
TASK_PP(16'hE012,4);
TASK_PP(16'hE013,4);
TASK_PP(16'hE014,4);
TASK_PP(16'hE015,4);
TASK_PP(16'hE016,4);
TASK_PP(16'hE017,4);
TASK_PP(16'hE018,4);
TASK_PP(16'hE019,4);
TASK_PP(16'hE01A,4);
TASK_PP(16'hE01B,4);
TASK_PP(16'hE01C,4);
TASK_PP(16'hE01D,4);
TASK_PP(16'hE01E,4);
TASK_PP(16'hE01F,4);
TASK_PP(16'hE020,4);
TASK_PP(16'hE021,4);
TASK_PP(16'hE022,4);
TASK_PP(16'hE023,4);
TASK_PP(16'hE024,4);
TASK_PP(16'hE025,4);
TASK_PP(16'hE026,4);
TASK_PP(16'hE027,4);
TASK_PP(16'hE028,4);
TASK_PP(16'hE029,4);
TASK_PP(16'hE02A,4);
TASK_PP(16'hE02B,4);
TASK_PP(16'hE02C,4);
TASK_PP(16'hE02D,4);
TASK_PP(16'hE02E,4);
TASK_PP(16'hE02F,4);
TASK_PP(16'hE030,4);
TASK_PP(16'hE031,4);
TASK_PP(16'hE032,4);
TASK_PP(16'hE033,4);
TASK_PP(16'hE034,4);
TASK_PP(16'hE035,4);
TASK_PP(16'hE036,4);
TASK_PP(16'hE037,4);
TASK_PP(16'hE038,4);
TASK_PP(16'hE039,4);
TASK_PP(16'hE03A,4);
TASK_PP(16'hE03B,4);
TASK_PP(16'hE03C,4);
TASK_PP(16'hE03D,4);
TASK_PP(16'hE03E,4);
TASK_PP(16'hE03F,4);
TASK_PP(16'hE040,4);
TASK_PP(16'hE041,4);
TASK_PP(16'hE042,4);
TASK_PP(16'hE043,4);
TASK_PP(16'hE044,4);
TASK_PP(16'hE045,4);
TASK_PP(16'hE046,4);
TASK_PP(16'hE047,4);
TASK_PP(16'hE048,4);
TASK_PP(16'hE049,4);
TASK_PP(16'hE04A,4);
TASK_PP(16'hE04B,4);
TASK_PP(16'hE04C,4);
TASK_PP(16'hE04D,4);
TASK_PP(16'hE04E,4);
TASK_PP(16'hE04F,4);
TASK_PP(16'hE050,4);
TASK_PP(16'hE051,4);
TASK_PP(16'hE052,4);
TASK_PP(16'hE053,4);
TASK_PP(16'hE054,4);
TASK_PP(16'hE055,4);
TASK_PP(16'hE056,4);
TASK_PP(16'hE057,4);
TASK_PP(16'hE058,4);
TASK_PP(16'hE059,4);
TASK_PP(16'hE05A,4);
TASK_PP(16'hE05B,4);
TASK_PP(16'hE05C,4);
TASK_PP(16'hE05D,4);
TASK_PP(16'hE05E,4);
TASK_PP(16'hE05F,4);
TASK_PP(16'hE060,4);
TASK_PP(16'hE061,4);
TASK_PP(16'hE062,4);
TASK_PP(16'hE063,4);
TASK_PP(16'hE064,4);
TASK_PP(16'hE065,4);
TASK_PP(16'hE066,4);
TASK_PP(16'hE067,4);
TASK_PP(16'hE068,4);
TASK_PP(16'hE069,4);
TASK_PP(16'hE06A,4);
TASK_PP(16'hE06B,4);
TASK_PP(16'hE06C,4);
TASK_PP(16'hE06D,4);
TASK_PP(16'hE06E,4);
TASK_PP(16'hE06F,4);
TASK_PP(16'hE070,4);
TASK_PP(16'hE071,4);
TASK_PP(16'hE072,4);
TASK_PP(16'hE073,4);
TASK_PP(16'hE074,4);
TASK_PP(16'hE075,4);
TASK_PP(16'hE076,4);
TASK_PP(16'hE077,4);
TASK_PP(16'hE078,4);
TASK_PP(16'hE079,4);
TASK_PP(16'hE07A,4);
TASK_PP(16'hE07B,4);
TASK_PP(16'hE07C,4);
TASK_PP(16'hE07D,4);
TASK_PP(16'hE07E,4);
TASK_PP(16'hE07F,4);
TASK_PP(16'hE080,4);
TASK_PP(16'hE081,4);
TASK_PP(16'hE082,4);
TASK_PP(16'hE083,4);
TASK_PP(16'hE084,4);
TASK_PP(16'hE085,4);
TASK_PP(16'hE086,4);
TASK_PP(16'hE087,4);
TASK_PP(16'hE088,4);
TASK_PP(16'hE089,4);
TASK_PP(16'hE08A,4);
TASK_PP(16'hE08B,4);
TASK_PP(16'hE08C,4);
TASK_PP(16'hE08D,4);
TASK_PP(16'hE08E,4);
TASK_PP(16'hE08F,4);
TASK_PP(16'hE090,4);
TASK_PP(16'hE091,4);
TASK_PP(16'hE092,4);
TASK_PP(16'hE093,4);
TASK_PP(16'hE094,4);
TASK_PP(16'hE095,4);
TASK_PP(16'hE096,4);
TASK_PP(16'hE097,4);
TASK_PP(16'hE098,4);
TASK_PP(16'hE099,4);
TASK_PP(16'hE09A,4);
TASK_PP(16'hE09B,4);
TASK_PP(16'hE09C,4);
TASK_PP(16'hE09D,4);
TASK_PP(16'hE09E,4);
TASK_PP(16'hE09F,4);
TASK_PP(16'hE0A0,4);
TASK_PP(16'hE0A1,4);
TASK_PP(16'hE0A2,4);
TASK_PP(16'hE0A3,4);
TASK_PP(16'hE0A4,4);
TASK_PP(16'hE0A5,4);
TASK_PP(16'hE0A6,4);
TASK_PP(16'hE0A7,4);
TASK_PP(16'hE0A8,4);
TASK_PP(16'hE0A9,4);
TASK_PP(16'hE0AA,4);
TASK_PP(16'hE0AB,4);
TASK_PP(16'hE0AC,4);
TASK_PP(16'hE0AD,4);
TASK_PP(16'hE0AE,4);
TASK_PP(16'hE0AF,4);
TASK_PP(16'hE0B0,4);
TASK_PP(16'hE0B1,4);
TASK_PP(16'hE0B2,4);
TASK_PP(16'hE0B3,4);
TASK_PP(16'hE0B4,4);
TASK_PP(16'hE0B5,4);
TASK_PP(16'hE0B6,4);
TASK_PP(16'hE0B7,4);
TASK_PP(16'hE0B8,4);
TASK_PP(16'hE0B9,4);
TASK_PP(16'hE0BA,4);
TASK_PP(16'hE0BB,4);
TASK_PP(16'hE0BC,4);
TASK_PP(16'hE0BD,4);
TASK_PP(16'hE0BE,4);
TASK_PP(16'hE0BF,4);
TASK_PP(16'hE0C0,4);
TASK_PP(16'hE0C1,4);
TASK_PP(16'hE0C2,4);
TASK_PP(16'hE0C3,4);
TASK_PP(16'hE0C4,4);
TASK_PP(16'hE0C5,4);
TASK_PP(16'hE0C6,4);
TASK_PP(16'hE0C7,4);
TASK_PP(16'hE0C8,4);
TASK_PP(16'hE0C9,4);
TASK_PP(16'hE0CA,4);
TASK_PP(16'hE0CB,4);
TASK_PP(16'hE0CC,4);
TASK_PP(16'hE0CD,4);
TASK_PP(16'hE0CE,4);
TASK_PP(16'hE0CF,4);
TASK_PP(16'hE0D0,4);
TASK_PP(16'hE0D1,4);
TASK_PP(16'hE0D2,4);
TASK_PP(16'hE0D3,4);
TASK_PP(16'hE0D4,4);
TASK_PP(16'hE0D5,4);
TASK_PP(16'hE0D6,4);
TASK_PP(16'hE0D7,4);
TASK_PP(16'hE0D8,4);
TASK_PP(16'hE0D9,4);
TASK_PP(16'hE0DA,4);
TASK_PP(16'hE0DB,4);
TASK_PP(16'hE0DC,4);
TASK_PP(16'hE0DD,4);
TASK_PP(16'hE0DE,4);
TASK_PP(16'hE0DF,4);
TASK_PP(16'hE0E0,4);
TASK_PP(16'hE0E1,4);
TASK_PP(16'hE0E2,4);
TASK_PP(16'hE0E3,4);
TASK_PP(16'hE0E4,4);
TASK_PP(16'hE0E5,4);
TASK_PP(16'hE0E6,4);
TASK_PP(16'hE0E7,4);
TASK_PP(16'hE0E8,4);
TASK_PP(16'hE0E9,4);
TASK_PP(16'hE0EA,4);
TASK_PP(16'hE0EB,4);
TASK_PP(16'hE0EC,4);
TASK_PP(16'hE0ED,4);
TASK_PP(16'hE0EE,4);
TASK_PP(16'hE0EF,4);
TASK_PP(16'hE0F0,4);
TASK_PP(16'hE0F1,4);
TASK_PP(16'hE0F2,4);
TASK_PP(16'hE0F3,4);
TASK_PP(16'hE0F4,4);
TASK_PP(16'hE0F5,4);
TASK_PP(16'hE0F6,4);
TASK_PP(16'hE0F7,4);
TASK_PP(16'hE0F8,4);
TASK_PP(16'hE0F9,4);
TASK_PP(16'hE0FA,4);
TASK_PP(16'hE0FB,4);
TASK_PP(16'hE0FC,4);
TASK_PP(16'hE0FD,4);
TASK_PP(16'hE0FE,4);
TASK_PP(16'hE0FF,4);
TASK_PP(16'hE100,4);
TASK_PP(16'hE101,4);
TASK_PP(16'hE102,4);
TASK_PP(16'hE103,4);
TASK_PP(16'hE104,4);
TASK_PP(16'hE105,4);
TASK_PP(16'hE106,4);
TASK_PP(16'hE107,4);
TASK_PP(16'hE108,4);
TASK_PP(16'hE109,4);
TASK_PP(16'hE10A,4);
TASK_PP(16'hE10B,4);
TASK_PP(16'hE10C,4);
TASK_PP(16'hE10D,4);
TASK_PP(16'hE10E,4);
TASK_PP(16'hE10F,4);
TASK_PP(16'hE110,4);
TASK_PP(16'hE111,4);
TASK_PP(16'hE112,4);
TASK_PP(16'hE113,4);
TASK_PP(16'hE114,4);
TASK_PP(16'hE115,4);
TASK_PP(16'hE116,4);
TASK_PP(16'hE117,4);
TASK_PP(16'hE118,4);
TASK_PP(16'hE119,4);
TASK_PP(16'hE11A,4);
TASK_PP(16'hE11B,4);
TASK_PP(16'hE11C,4);
TASK_PP(16'hE11D,4);
TASK_PP(16'hE11E,4);
TASK_PP(16'hE11F,4);
TASK_PP(16'hE120,4);
TASK_PP(16'hE121,4);
TASK_PP(16'hE122,4);
TASK_PP(16'hE123,4);
TASK_PP(16'hE124,4);
TASK_PP(16'hE125,4);
TASK_PP(16'hE126,4);
TASK_PP(16'hE127,4);
TASK_PP(16'hE128,4);
TASK_PP(16'hE129,4);
TASK_PP(16'hE12A,4);
TASK_PP(16'hE12B,4);
TASK_PP(16'hE12C,4);
TASK_PP(16'hE12D,4);
TASK_PP(16'hE12E,4);
TASK_PP(16'hE12F,4);
TASK_PP(16'hE130,4);
TASK_PP(16'hE131,4);
TASK_PP(16'hE132,4);
TASK_PP(16'hE133,4);
TASK_PP(16'hE134,4);
TASK_PP(16'hE135,4);
TASK_PP(16'hE136,4);
TASK_PP(16'hE137,4);
TASK_PP(16'hE138,4);
TASK_PP(16'hE139,4);
TASK_PP(16'hE13A,4);
TASK_PP(16'hE13B,4);
TASK_PP(16'hE13C,4);
TASK_PP(16'hE13D,4);
TASK_PP(16'hE13E,4);
TASK_PP(16'hE13F,4);
TASK_PP(16'hE140,4);
TASK_PP(16'hE141,4);
TASK_PP(16'hE142,4);
TASK_PP(16'hE143,4);
TASK_PP(16'hE144,4);
TASK_PP(16'hE145,4);
TASK_PP(16'hE146,4);
TASK_PP(16'hE147,4);
TASK_PP(16'hE148,4);
TASK_PP(16'hE149,4);
TASK_PP(16'hE14A,4);
TASK_PP(16'hE14B,4);
TASK_PP(16'hE14C,4);
TASK_PP(16'hE14D,4);
TASK_PP(16'hE14E,4);
TASK_PP(16'hE14F,4);
TASK_PP(16'hE150,4);
TASK_PP(16'hE151,4);
TASK_PP(16'hE152,4);
TASK_PP(16'hE153,4);
TASK_PP(16'hE154,4);
TASK_PP(16'hE155,4);
TASK_PP(16'hE156,4);
TASK_PP(16'hE157,4);
TASK_PP(16'hE158,4);
TASK_PP(16'hE159,4);
TASK_PP(16'hE15A,4);
TASK_PP(16'hE15B,4);
TASK_PP(16'hE15C,4);
TASK_PP(16'hE15D,4);
TASK_PP(16'hE15E,4);
TASK_PP(16'hE15F,4);
TASK_PP(16'hE160,4);
TASK_PP(16'hE161,4);
TASK_PP(16'hE162,4);
TASK_PP(16'hE163,4);
TASK_PP(16'hE164,4);
TASK_PP(16'hE165,4);
TASK_PP(16'hE166,4);
TASK_PP(16'hE167,4);
TASK_PP(16'hE168,4);
TASK_PP(16'hE169,4);
TASK_PP(16'hE16A,4);
TASK_PP(16'hE16B,4);
TASK_PP(16'hE16C,4);
TASK_PP(16'hE16D,4);
TASK_PP(16'hE16E,4);
TASK_PP(16'hE16F,4);
TASK_PP(16'hE170,4);
TASK_PP(16'hE171,4);
TASK_PP(16'hE172,4);
TASK_PP(16'hE173,4);
TASK_PP(16'hE174,4);
TASK_PP(16'hE175,4);
TASK_PP(16'hE176,4);
TASK_PP(16'hE177,4);
TASK_PP(16'hE178,4);
TASK_PP(16'hE179,4);
TASK_PP(16'hE17A,4);
TASK_PP(16'hE17B,4);
TASK_PP(16'hE17C,4);
TASK_PP(16'hE17D,4);
TASK_PP(16'hE17E,4);
TASK_PP(16'hE17F,4);
TASK_PP(16'hE180,4);
TASK_PP(16'hE181,4);
TASK_PP(16'hE182,4);
TASK_PP(16'hE183,4);
TASK_PP(16'hE184,4);
TASK_PP(16'hE185,4);
TASK_PP(16'hE186,4);
TASK_PP(16'hE187,4);
TASK_PP(16'hE188,4);
TASK_PP(16'hE189,4);
TASK_PP(16'hE18A,4);
TASK_PP(16'hE18B,4);
TASK_PP(16'hE18C,4);
TASK_PP(16'hE18D,4);
TASK_PP(16'hE18E,4);
TASK_PP(16'hE18F,4);
TASK_PP(16'hE190,4);
TASK_PP(16'hE191,4);
TASK_PP(16'hE192,4);
TASK_PP(16'hE193,4);
TASK_PP(16'hE194,4);
TASK_PP(16'hE195,4);
TASK_PP(16'hE196,4);
TASK_PP(16'hE197,4);
TASK_PP(16'hE198,4);
TASK_PP(16'hE199,4);
TASK_PP(16'hE19A,4);
TASK_PP(16'hE19B,4);
TASK_PP(16'hE19C,4);
TASK_PP(16'hE19D,4);
TASK_PP(16'hE19E,4);
TASK_PP(16'hE19F,4);
TASK_PP(16'hE1A0,4);
TASK_PP(16'hE1A1,4);
TASK_PP(16'hE1A2,4);
TASK_PP(16'hE1A3,4);
TASK_PP(16'hE1A4,4);
TASK_PP(16'hE1A5,4);
TASK_PP(16'hE1A6,4);
TASK_PP(16'hE1A7,4);
TASK_PP(16'hE1A8,4);
TASK_PP(16'hE1A9,4);
TASK_PP(16'hE1AA,4);
TASK_PP(16'hE1AB,4);
TASK_PP(16'hE1AC,4);
TASK_PP(16'hE1AD,4);
TASK_PP(16'hE1AE,4);
TASK_PP(16'hE1AF,4);
TASK_PP(16'hE1B0,4);
TASK_PP(16'hE1B1,4);
TASK_PP(16'hE1B2,4);
TASK_PP(16'hE1B3,4);
TASK_PP(16'hE1B4,4);
TASK_PP(16'hE1B5,4);
TASK_PP(16'hE1B6,4);
TASK_PP(16'hE1B7,4);
TASK_PP(16'hE1B8,4);
TASK_PP(16'hE1B9,4);
TASK_PP(16'hE1BA,4);
TASK_PP(16'hE1BB,4);
TASK_PP(16'hE1BC,4);
TASK_PP(16'hE1BD,4);
TASK_PP(16'hE1BE,4);
TASK_PP(16'hE1BF,4);
TASK_PP(16'hE1C0,4);
TASK_PP(16'hE1C1,4);
TASK_PP(16'hE1C2,4);
TASK_PP(16'hE1C3,4);
TASK_PP(16'hE1C4,4);
TASK_PP(16'hE1C5,4);
TASK_PP(16'hE1C6,4);
TASK_PP(16'hE1C7,4);
TASK_PP(16'hE1C8,4);
TASK_PP(16'hE1C9,4);
TASK_PP(16'hE1CA,4);
TASK_PP(16'hE1CB,4);
TASK_PP(16'hE1CC,4);
TASK_PP(16'hE1CD,4);
TASK_PP(16'hE1CE,4);
TASK_PP(16'hE1CF,4);
TASK_PP(16'hE1D0,4);
TASK_PP(16'hE1D1,4);
TASK_PP(16'hE1D2,4);
TASK_PP(16'hE1D3,4);
TASK_PP(16'hE1D4,4);
TASK_PP(16'hE1D5,4);
TASK_PP(16'hE1D6,4);
TASK_PP(16'hE1D7,4);
TASK_PP(16'hE1D8,4);
TASK_PP(16'hE1D9,4);
TASK_PP(16'hE1DA,4);
TASK_PP(16'hE1DB,4);
TASK_PP(16'hE1DC,4);
TASK_PP(16'hE1DD,4);
TASK_PP(16'hE1DE,4);
TASK_PP(16'hE1DF,4);
TASK_PP(16'hE1E0,4);
TASK_PP(16'hE1E1,4);
TASK_PP(16'hE1E2,4);
TASK_PP(16'hE1E3,4);
TASK_PP(16'hE1E4,4);
TASK_PP(16'hE1E5,4);
TASK_PP(16'hE1E6,4);
TASK_PP(16'hE1E7,4);
TASK_PP(16'hE1E8,4);
TASK_PP(16'hE1E9,4);
TASK_PP(16'hE1EA,4);
TASK_PP(16'hE1EB,4);
TASK_PP(16'hE1EC,4);
TASK_PP(16'hE1ED,4);
TASK_PP(16'hE1EE,4);
TASK_PP(16'hE1EF,4);
TASK_PP(16'hE1F0,4);
TASK_PP(16'hE1F1,4);
TASK_PP(16'hE1F2,4);
TASK_PP(16'hE1F3,4);
TASK_PP(16'hE1F4,4);
TASK_PP(16'hE1F5,4);
TASK_PP(16'hE1F6,4);
TASK_PP(16'hE1F7,4);
TASK_PP(16'hE1F8,4);
TASK_PP(16'hE1F9,4);
TASK_PP(16'hE1FA,4);
TASK_PP(16'hE1FB,4);
TASK_PP(16'hE1FC,4);
TASK_PP(16'hE1FD,4);
TASK_PP(16'hE1FE,4);
TASK_PP(16'hE1FF,4);
TASK_PP(16'hE200,4);
TASK_PP(16'hE201,4);
TASK_PP(16'hE202,4);
TASK_PP(16'hE203,4);
TASK_PP(16'hE204,4);
TASK_PP(16'hE205,4);
TASK_PP(16'hE206,4);
TASK_PP(16'hE207,4);
TASK_PP(16'hE208,4);
TASK_PP(16'hE209,4);
TASK_PP(16'hE20A,4);
TASK_PP(16'hE20B,4);
TASK_PP(16'hE20C,4);
TASK_PP(16'hE20D,4);
TASK_PP(16'hE20E,4);
TASK_PP(16'hE20F,4);
TASK_PP(16'hE210,4);
TASK_PP(16'hE211,4);
TASK_PP(16'hE212,4);
TASK_PP(16'hE213,4);
TASK_PP(16'hE214,4);
TASK_PP(16'hE215,4);
TASK_PP(16'hE216,4);
TASK_PP(16'hE217,4);
TASK_PP(16'hE218,4);
TASK_PP(16'hE219,4);
TASK_PP(16'hE21A,4);
TASK_PP(16'hE21B,4);
TASK_PP(16'hE21C,4);
TASK_PP(16'hE21D,4);
TASK_PP(16'hE21E,4);
TASK_PP(16'hE21F,4);
TASK_PP(16'hE220,4);
TASK_PP(16'hE221,4);
TASK_PP(16'hE222,4);
TASK_PP(16'hE223,4);
TASK_PP(16'hE224,4);
TASK_PP(16'hE225,4);
TASK_PP(16'hE226,4);
TASK_PP(16'hE227,4);
TASK_PP(16'hE228,4);
TASK_PP(16'hE229,4);
TASK_PP(16'hE22A,4);
TASK_PP(16'hE22B,4);
TASK_PP(16'hE22C,4);
TASK_PP(16'hE22D,4);
TASK_PP(16'hE22E,4);
TASK_PP(16'hE22F,4);
TASK_PP(16'hE230,4);
TASK_PP(16'hE231,4);
TASK_PP(16'hE232,4);
TASK_PP(16'hE233,4);
TASK_PP(16'hE234,4);
TASK_PP(16'hE235,4);
TASK_PP(16'hE236,4);
TASK_PP(16'hE237,4);
TASK_PP(16'hE238,4);
TASK_PP(16'hE239,4);
TASK_PP(16'hE23A,4);
TASK_PP(16'hE23B,4);
TASK_PP(16'hE23C,4);
TASK_PP(16'hE23D,4);
TASK_PP(16'hE23E,4);
TASK_PP(16'hE23F,4);
TASK_PP(16'hE240,4);
TASK_PP(16'hE241,4);
TASK_PP(16'hE242,4);
TASK_PP(16'hE243,4);
TASK_PP(16'hE244,4);
TASK_PP(16'hE245,4);
TASK_PP(16'hE246,4);
TASK_PP(16'hE247,4);
TASK_PP(16'hE248,4);
TASK_PP(16'hE249,4);
TASK_PP(16'hE24A,4);
TASK_PP(16'hE24B,4);
TASK_PP(16'hE24C,4);
TASK_PP(16'hE24D,4);
TASK_PP(16'hE24E,4);
TASK_PP(16'hE24F,4);
TASK_PP(16'hE250,4);
TASK_PP(16'hE251,4);
TASK_PP(16'hE252,4);
TASK_PP(16'hE253,4);
TASK_PP(16'hE254,4);
TASK_PP(16'hE255,4);
TASK_PP(16'hE256,4);
TASK_PP(16'hE257,4);
TASK_PP(16'hE258,4);
TASK_PP(16'hE259,4);
TASK_PP(16'hE25A,4);
TASK_PP(16'hE25B,4);
TASK_PP(16'hE25C,4);
TASK_PP(16'hE25D,4);
TASK_PP(16'hE25E,4);
TASK_PP(16'hE25F,4);
TASK_PP(16'hE260,4);
TASK_PP(16'hE261,4);
TASK_PP(16'hE262,4);
TASK_PP(16'hE263,4);
TASK_PP(16'hE264,4);
TASK_PP(16'hE265,4);
TASK_PP(16'hE266,4);
TASK_PP(16'hE267,4);
TASK_PP(16'hE268,4);
TASK_PP(16'hE269,4);
TASK_PP(16'hE26A,4);
TASK_PP(16'hE26B,4);
TASK_PP(16'hE26C,4);
TASK_PP(16'hE26D,4);
TASK_PP(16'hE26E,4);
TASK_PP(16'hE26F,4);
TASK_PP(16'hE270,4);
TASK_PP(16'hE271,4);
TASK_PP(16'hE272,4);
TASK_PP(16'hE273,4);
TASK_PP(16'hE274,4);
TASK_PP(16'hE275,4);
TASK_PP(16'hE276,4);
TASK_PP(16'hE277,4);
TASK_PP(16'hE278,4);
TASK_PP(16'hE279,4);
TASK_PP(16'hE27A,4);
TASK_PP(16'hE27B,4);
TASK_PP(16'hE27C,4);
TASK_PP(16'hE27D,4);
TASK_PP(16'hE27E,4);
TASK_PP(16'hE27F,4);
TASK_PP(16'hE280,4);
TASK_PP(16'hE281,4);
TASK_PP(16'hE282,4);
TASK_PP(16'hE283,4);
TASK_PP(16'hE284,4);
TASK_PP(16'hE285,4);
TASK_PP(16'hE286,4);
TASK_PP(16'hE287,4);
TASK_PP(16'hE288,4);
TASK_PP(16'hE289,4);
TASK_PP(16'hE28A,4);
TASK_PP(16'hE28B,4);
TASK_PP(16'hE28C,4);
TASK_PP(16'hE28D,4);
TASK_PP(16'hE28E,4);
TASK_PP(16'hE28F,4);
TASK_PP(16'hE290,4);
TASK_PP(16'hE291,4);
TASK_PP(16'hE292,4);
TASK_PP(16'hE293,4);
TASK_PP(16'hE294,4);
TASK_PP(16'hE295,4);
TASK_PP(16'hE296,4);
TASK_PP(16'hE297,4);
TASK_PP(16'hE298,4);
TASK_PP(16'hE299,4);
TASK_PP(16'hE29A,4);
TASK_PP(16'hE29B,4);
TASK_PP(16'hE29C,4);
TASK_PP(16'hE29D,4);
TASK_PP(16'hE29E,4);
TASK_PP(16'hE29F,4);
TASK_PP(16'hE2A0,4);
TASK_PP(16'hE2A1,4);
TASK_PP(16'hE2A2,4);
TASK_PP(16'hE2A3,4);
TASK_PP(16'hE2A4,4);
TASK_PP(16'hE2A5,4);
TASK_PP(16'hE2A6,4);
TASK_PP(16'hE2A7,4);
TASK_PP(16'hE2A8,4);
TASK_PP(16'hE2A9,4);
TASK_PP(16'hE2AA,4);
TASK_PP(16'hE2AB,4);
TASK_PP(16'hE2AC,4);
TASK_PP(16'hE2AD,4);
TASK_PP(16'hE2AE,4);
TASK_PP(16'hE2AF,4);
TASK_PP(16'hE2B0,4);
TASK_PP(16'hE2B1,4);
TASK_PP(16'hE2B2,4);
TASK_PP(16'hE2B3,4);
TASK_PP(16'hE2B4,4);
TASK_PP(16'hE2B5,4);
TASK_PP(16'hE2B6,4);
TASK_PP(16'hE2B7,4);
TASK_PP(16'hE2B8,4);
TASK_PP(16'hE2B9,4);
TASK_PP(16'hE2BA,4);
TASK_PP(16'hE2BB,4);
TASK_PP(16'hE2BC,4);
TASK_PP(16'hE2BD,4);
TASK_PP(16'hE2BE,4);
TASK_PP(16'hE2BF,4);
TASK_PP(16'hE2C0,4);
TASK_PP(16'hE2C1,4);
TASK_PP(16'hE2C2,4);
TASK_PP(16'hE2C3,4);
TASK_PP(16'hE2C4,4);
TASK_PP(16'hE2C5,4);
TASK_PP(16'hE2C6,4);
TASK_PP(16'hE2C7,4);
TASK_PP(16'hE2C8,4);
TASK_PP(16'hE2C9,4);
TASK_PP(16'hE2CA,4);
TASK_PP(16'hE2CB,4);
TASK_PP(16'hE2CC,4);
TASK_PP(16'hE2CD,4);
TASK_PP(16'hE2CE,4);
TASK_PP(16'hE2CF,4);
TASK_PP(16'hE2D0,4);
TASK_PP(16'hE2D1,4);
TASK_PP(16'hE2D2,4);
TASK_PP(16'hE2D3,4);
TASK_PP(16'hE2D4,4);
TASK_PP(16'hE2D5,4);
TASK_PP(16'hE2D6,4);
TASK_PP(16'hE2D7,4);
TASK_PP(16'hE2D8,4);
TASK_PP(16'hE2D9,4);
TASK_PP(16'hE2DA,4);
TASK_PP(16'hE2DB,4);
TASK_PP(16'hE2DC,4);
TASK_PP(16'hE2DD,4);
TASK_PP(16'hE2DE,4);
TASK_PP(16'hE2DF,4);
TASK_PP(16'hE2E0,4);
TASK_PP(16'hE2E1,4);
TASK_PP(16'hE2E2,4);
TASK_PP(16'hE2E3,4);
TASK_PP(16'hE2E4,4);
TASK_PP(16'hE2E5,4);
TASK_PP(16'hE2E6,4);
TASK_PP(16'hE2E7,4);
TASK_PP(16'hE2E8,4);
TASK_PP(16'hE2E9,4);
TASK_PP(16'hE2EA,4);
TASK_PP(16'hE2EB,4);
TASK_PP(16'hE2EC,4);
TASK_PP(16'hE2ED,4);
TASK_PP(16'hE2EE,4);
TASK_PP(16'hE2EF,4);
TASK_PP(16'hE2F0,4);
TASK_PP(16'hE2F1,4);
TASK_PP(16'hE2F2,4);
TASK_PP(16'hE2F3,4);
TASK_PP(16'hE2F4,4);
TASK_PP(16'hE2F5,4);
TASK_PP(16'hE2F6,4);
TASK_PP(16'hE2F7,4);
TASK_PP(16'hE2F8,4);
TASK_PP(16'hE2F9,4);
TASK_PP(16'hE2FA,4);
TASK_PP(16'hE2FB,4);
TASK_PP(16'hE2FC,4);
TASK_PP(16'hE2FD,4);
TASK_PP(16'hE2FE,4);
TASK_PP(16'hE2FF,4);
TASK_PP(16'hE300,4);
TASK_PP(16'hE301,4);
TASK_PP(16'hE302,4);
TASK_PP(16'hE303,4);
TASK_PP(16'hE304,4);
TASK_PP(16'hE305,4);
TASK_PP(16'hE306,4);
TASK_PP(16'hE307,4);
TASK_PP(16'hE308,4);
TASK_PP(16'hE309,4);
TASK_PP(16'hE30A,4);
TASK_PP(16'hE30B,4);
TASK_PP(16'hE30C,4);
TASK_PP(16'hE30D,4);
TASK_PP(16'hE30E,4);
TASK_PP(16'hE30F,4);
TASK_PP(16'hE310,4);
TASK_PP(16'hE311,4);
TASK_PP(16'hE312,4);
TASK_PP(16'hE313,4);
TASK_PP(16'hE314,4);
TASK_PP(16'hE315,4);
TASK_PP(16'hE316,4);
TASK_PP(16'hE317,4);
TASK_PP(16'hE318,4);
TASK_PP(16'hE319,4);
TASK_PP(16'hE31A,4);
TASK_PP(16'hE31B,4);
TASK_PP(16'hE31C,4);
TASK_PP(16'hE31D,4);
TASK_PP(16'hE31E,4);
TASK_PP(16'hE31F,4);
TASK_PP(16'hE320,4);
TASK_PP(16'hE321,4);
TASK_PP(16'hE322,4);
TASK_PP(16'hE323,4);
TASK_PP(16'hE324,4);
TASK_PP(16'hE325,4);
TASK_PP(16'hE326,4);
TASK_PP(16'hE327,4);
TASK_PP(16'hE328,4);
TASK_PP(16'hE329,4);
TASK_PP(16'hE32A,4);
TASK_PP(16'hE32B,4);
TASK_PP(16'hE32C,4);
TASK_PP(16'hE32D,4);
TASK_PP(16'hE32E,4);
TASK_PP(16'hE32F,4);
TASK_PP(16'hE330,4);
TASK_PP(16'hE331,4);
TASK_PP(16'hE332,4);
TASK_PP(16'hE333,4);
TASK_PP(16'hE334,4);
TASK_PP(16'hE335,4);
TASK_PP(16'hE336,4);
TASK_PP(16'hE337,4);
TASK_PP(16'hE338,4);
TASK_PP(16'hE339,4);
TASK_PP(16'hE33A,4);
TASK_PP(16'hE33B,4);
TASK_PP(16'hE33C,4);
TASK_PP(16'hE33D,4);
TASK_PP(16'hE33E,4);
TASK_PP(16'hE33F,4);
TASK_PP(16'hE340,4);
TASK_PP(16'hE341,4);
TASK_PP(16'hE342,4);
TASK_PP(16'hE343,4);
TASK_PP(16'hE344,4);
TASK_PP(16'hE345,4);
TASK_PP(16'hE346,4);
TASK_PP(16'hE347,4);
TASK_PP(16'hE348,4);
TASK_PP(16'hE349,4);
TASK_PP(16'hE34A,4);
TASK_PP(16'hE34B,4);
TASK_PP(16'hE34C,4);
TASK_PP(16'hE34D,4);
TASK_PP(16'hE34E,4);
TASK_PP(16'hE34F,4);
TASK_PP(16'hE350,4);
TASK_PP(16'hE351,4);
TASK_PP(16'hE352,4);
TASK_PP(16'hE353,4);
TASK_PP(16'hE354,4);
TASK_PP(16'hE355,4);
TASK_PP(16'hE356,4);
TASK_PP(16'hE357,4);
TASK_PP(16'hE358,4);
TASK_PP(16'hE359,4);
TASK_PP(16'hE35A,4);
TASK_PP(16'hE35B,4);
TASK_PP(16'hE35C,4);
TASK_PP(16'hE35D,4);
TASK_PP(16'hE35E,4);
TASK_PP(16'hE35F,4);
TASK_PP(16'hE360,4);
TASK_PP(16'hE361,4);
TASK_PP(16'hE362,4);
TASK_PP(16'hE363,4);
TASK_PP(16'hE364,4);
TASK_PP(16'hE365,4);
TASK_PP(16'hE366,4);
TASK_PP(16'hE367,4);
TASK_PP(16'hE368,4);
TASK_PP(16'hE369,4);
TASK_PP(16'hE36A,4);
TASK_PP(16'hE36B,4);
TASK_PP(16'hE36C,4);
TASK_PP(16'hE36D,4);
TASK_PP(16'hE36E,4);
TASK_PP(16'hE36F,4);
TASK_PP(16'hE370,4);
TASK_PP(16'hE371,4);
TASK_PP(16'hE372,4);
TASK_PP(16'hE373,4);
TASK_PP(16'hE374,4);
TASK_PP(16'hE375,4);
TASK_PP(16'hE376,4);
TASK_PP(16'hE377,4);
TASK_PP(16'hE378,4);
TASK_PP(16'hE379,4);
TASK_PP(16'hE37A,4);
TASK_PP(16'hE37B,4);
TASK_PP(16'hE37C,4);
TASK_PP(16'hE37D,4);
TASK_PP(16'hE37E,4);
TASK_PP(16'hE37F,4);
TASK_PP(16'hE380,4);
TASK_PP(16'hE381,4);
TASK_PP(16'hE382,4);
TASK_PP(16'hE383,4);
TASK_PP(16'hE384,4);
TASK_PP(16'hE385,4);
TASK_PP(16'hE386,4);
TASK_PP(16'hE387,4);
TASK_PP(16'hE388,4);
TASK_PP(16'hE389,4);
TASK_PP(16'hE38A,4);
TASK_PP(16'hE38B,4);
TASK_PP(16'hE38C,4);
TASK_PP(16'hE38D,4);
TASK_PP(16'hE38E,4);
TASK_PP(16'hE38F,4);
TASK_PP(16'hE390,4);
TASK_PP(16'hE391,4);
TASK_PP(16'hE392,4);
TASK_PP(16'hE393,4);
TASK_PP(16'hE394,4);
TASK_PP(16'hE395,4);
TASK_PP(16'hE396,4);
TASK_PP(16'hE397,4);
TASK_PP(16'hE398,4);
TASK_PP(16'hE399,4);
TASK_PP(16'hE39A,4);
TASK_PP(16'hE39B,4);
TASK_PP(16'hE39C,4);
TASK_PP(16'hE39D,4);
TASK_PP(16'hE39E,4);
TASK_PP(16'hE39F,4);
TASK_PP(16'hE3A0,4);
TASK_PP(16'hE3A1,4);
TASK_PP(16'hE3A2,4);
TASK_PP(16'hE3A3,4);
TASK_PP(16'hE3A4,4);
TASK_PP(16'hE3A5,4);
TASK_PP(16'hE3A6,4);
TASK_PP(16'hE3A7,4);
TASK_PP(16'hE3A8,4);
TASK_PP(16'hE3A9,4);
TASK_PP(16'hE3AA,4);
TASK_PP(16'hE3AB,4);
TASK_PP(16'hE3AC,4);
TASK_PP(16'hE3AD,4);
TASK_PP(16'hE3AE,4);
TASK_PP(16'hE3AF,4);
TASK_PP(16'hE3B0,4);
TASK_PP(16'hE3B1,4);
TASK_PP(16'hE3B2,4);
TASK_PP(16'hE3B3,4);
TASK_PP(16'hE3B4,4);
TASK_PP(16'hE3B5,4);
TASK_PP(16'hE3B6,4);
TASK_PP(16'hE3B7,4);
TASK_PP(16'hE3B8,4);
TASK_PP(16'hE3B9,4);
TASK_PP(16'hE3BA,4);
TASK_PP(16'hE3BB,4);
TASK_PP(16'hE3BC,4);
TASK_PP(16'hE3BD,4);
TASK_PP(16'hE3BE,4);
TASK_PP(16'hE3BF,4);
TASK_PP(16'hE3C0,4);
TASK_PP(16'hE3C1,4);
TASK_PP(16'hE3C2,4);
TASK_PP(16'hE3C3,4);
TASK_PP(16'hE3C4,4);
TASK_PP(16'hE3C5,4);
TASK_PP(16'hE3C6,4);
TASK_PP(16'hE3C7,4);
TASK_PP(16'hE3C8,4);
TASK_PP(16'hE3C9,4);
TASK_PP(16'hE3CA,4);
TASK_PP(16'hE3CB,4);
TASK_PP(16'hE3CC,4);
TASK_PP(16'hE3CD,4);
TASK_PP(16'hE3CE,4);
TASK_PP(16'hE3CF,4);
TASK_PP(16'hE3D0,4);
TASK_PP(16'hE3D1,4);
TASK_PP(16'hE3D2,4);
TASK_PP(16'hE3D3,4);
TASK_PP(16'hE3D4,4);
TASK_PP(16'hE3D5,4);
TASK_PP(16'hE3D6,4);
TASK_PP(16'hE3D7,4);
TASK_PP(16'hE3D8,4);
TASK_PP(16'hE3D9,4);
TASK_PP(16'hE3DA,4);
TASK_PP(16'hE3DB,4);
TASK_PP(16'hE3DC,4);
TASK_PP(16'hE3DD,4);
TASK_PP(16'hE3DE,4);
TASK_PP(16'hE3DF,4);
TASK_PP(16'hE3E0,4);
TASK_PP(16'hE3E1,4);
TASK_PP(16'hE3E2,4);
TASK_PP(16'hE3E3,4);
TASK_PP(16'hE3E4,4);
TASK_PP(16'hE3E5,4);
TASK_PP(16'hE3E6,4);
TASK_PP(16'hE3E7,4);
TASK_PP(16'hE3E8,4);
TASK_PP(16'hE3E9,4);
TASK_PP(16'hE3EA,4);
TASK_PP(16'hE3EB,4);
TASK_PP(16'hE3EC,4);
TASK_PP(16'hE3ED,4);
TASK_PP(16'hE3EE,4);
TASK_PP(16'hE3EF,4);
TASK_PP(16'hE3F0,4);
TASK_PP(16'hE3F1,4);
TASK_PP(16'hE3F2,4);
TASK_PP(16'hE3F3,4);
TASK_PP(16'hE3F4,4);
TASK_PP(16'hE3F5,4);
TASK_PP(16'hE3F6,4);
TASK_PP(16'hE3F7,4);
TASK_PP(16'hE3F8,4);
TASK_PP(16'hE3F9,4);
TASK_PP(16'hE3FA,4);
TASK_PP(16'hE3FB,4);
TASK_PP(16'hE3FC,4);
TASK_PP(16'hE3FD,4);
TASK_PP(16'hE3FE,4);
TASK_PP(16'hE3FF,4);
TASK_PP(16'hE400,4);
TASK_PP(16'hE401,4);
TASK_PP(16'hE402,4);
TASK_PP(16'hE403,4);
TASK_PP(16'hE404,4);
TASK_PP(16'hE405,4);
TASK_PP(16'hE406,4);
TASK_PP(16'hE407,4);
TASK_PP(16'hE408,4);
TASK_PP(16'hE409,4);
TASK_PP(16'hE40A,4);
TASK_PP(16'hE40B,4);
TASK_PP(16'hE40C,4);
TASK_PP(16'hE40D,4);
TASK_PP(16'hE40E,4);
TASK_PP(16'hE40F,4);
TASK_PP(16'hE410,4);
TASK_PP(16'hE411,4);
TASK_PP(16'hE412,4);
TASK_PP(16'hE413,4);
TASK_PP(16'hE414,4);
TASK_PP(16'hE415,4);
TASK_PP(16'hE416,4);
TASK_PP(16'hE417,4);
TASK_PP(16'hE418,4);
TASK_PP(16'hE419,4);
TASK_PP(16'hE41A,4);
TASK_PP(16'hE41B,4);
TASK_PP(16'hE41C,4);
TASK_PP(16'hE41D,4);
TASK_PP(16'hE41E,4);
TASK_PP(16'hE41F,4);
TASK_PP(16'hE420,4);
TASK_PP(16'hE421,4);
TASK_PP(16'hE422,4);
TASK_PP(16'hE423,4);
TASK_PP(16'hE424,4);
TASK_PP(16'hE425,4);
TASK_PP(16'hE426,4);
TASK_PP(16'hE427,4);
TASK_PP(16'hE428,4);
TASK_PP(16'hE429,4);
TASK_PP(16'hE42A,4);
TASK_PP(16'hE42B,4);
TASK_PP(16'hE42C,4);
TASK_PP(16'hE42D,4);
TASK_PP(16'hE42E,4);
TASK_PP(16'hE42F,4);
TASK_PP(16'hE430,4);
TASK_PP(16'hE431,4);
TASK_PP(16'hE432,4);
TASK_PP(16'hE433,4);
TASK_PP(16'hE434,4);
TASK_PP(16'hE435,4);
TASK_PP(16'hE436,4);
TASK_PP(16'hE437,4);
TASK_PP(16'hE438,4);
TASK_PP(16'hE439,4);
TASK_PP(16'hE43A,4);
TASK_PP(16'hE43B,4);
TASK_PP(16'hE43C,4);
TASK_PP(16'hE43D,4);
TASK_PP(16'hE43E,4);
TASK_PP(16'hE43F,4);
TASK_PP(16'hE440,4);
TASK_PP(16'hE441,4);
TASK_PP(16'hE442,4);
TASK_PP(16'hE443,4);
TASK_PP(16'hE444,4);
TASK_PP(16'hE445,4);
TASK_PP(16'hE446,4);
TASK_PP(16'hE447,4);
TASK_PP(16'hE448,4);
TASK_PP(16'hE449,4);
TASK_PP(16'hE44A,4);
TASK_PP(16'hE44B,4);
TASK_PP(16'hE44C,4);
TASK_PP(16'hE44D,4);
TASK_PP(16'hE44E,4);
TASK_PP(16'hE44F,4);
TASK_PP(16'hE450,4);
TASK_PP(16'hE451,4);
TASK_PP(16'hE452,4);
TASK_PP(16'hE453,4);
TASK_PP(16'hE454,4);
TASK_PP(16'hE455,4);
TASK_PP(16'hE456,4);
TASK_PP(16'hE457,4);
TASK_PP(16'hE458,4);
TASK_PP(16'hE459,4);
TASK_PP(16'hE45A,4);
TASK_PP(16'hE45B,4);
TASK_PP(16'hE45C,4);
TASK_PP(16'hE45D,4);
TASK_PP(16'hE45E,4);
TASK_PP(16'hE45F,4);
TASK_PP(16'hE460,4);
TASK_PP(16'hE461,4);
TASK_PP(16'hE462,4);
TASK_PP(16'hE463,4);
TASK_PP(16'hE464,4);
TASK_PP(16'hE465,4);
TASK_PP(16'hE466,4);
TASK_PP(16'hE467,4);
TASK_PP(16'hE468,4);
TASK_PP(16'hE469,4);
TASK_PP(16'hE46A,4);
TASK_PP(16'hE46B,4);
TASK_PP(16'hE46C,4);
TASK_PP(16'hE46D,4);
TASK_PP(16'hE46E,4);
TASK_PP(16'hE46F,4);
TASK_PP(16'hE470,4);
TASK_PP(16'hE471,4);
TASK_PP(16'hE472,4);
TASK_PP(16'hE473,4);
TASK_PP(16'hE474,4);
TASK_PP(16'hE475,4);
TASK_PP(16'hE476,4);
TASK_PP(16'hE477,4);
TASK_PP(16'hE478,4);
TASK_PP(16'hE479,4);
TASK_PP(16'hE47A,4);
TASK_PP(16'hE47B,4);
TASK_PP(16'hE47C,4);
TASK_PP(16'hE47D,4);
TASK_PP(16'hE47E,4);
TASK_PP(16'hE47F,4);
TASK_PP(16'hE480,4);
TASK_PP(16'hE481,4);
TASK_PP(16'hE482,4);
TASK_PP(16'hE483,4);
TASK_PP(16'hE484,4);
TASK_PP(16'hE485,4);
TASK_PP(16'hE486,4);
TASK_PP(16'hE487,4);
TASK_PP(16'hE488,4);
TASK_PP(16'hE489,4);
TASK_PP(16'hE48A,4);
TASK_PP(16'hE48B,4);
TASK_PP(16'hE48C,4);
TASK_PP(16'hE48D,4);
TASK_PP(16'hE48E,4);
TASK_PP(16'hE48F,4);
TASK_PP(16'hE490,4);
TASK_PP(16'hE491,4);
TASK_PP(16'hE492,4);
TASK_PP(16'hE493,4);
TASK_PP(16'hE494,4);
TASK_PP(16'hE495,4);
TASK_PP(16'hE496,4);
TASK_PP(16'hE497,4);
TASK_PP(16'hE498,4);
TASK_PP(16'hE499,4);
TASK_PP(16'hE49A,4);
TASK_PP(16'hE49B,4);
TASK_PP(16'hE49C,4);
TASK_PP(16'hE49D,4);
TASK_PP(16'hE49E,4);
TASK_PP(16'hE49F,4);
TASK_PP(16'hE4A0,4);
TASK_PP(16'hE4A1,4);
TASK_PP(16'hE4A2,4);
TASK_PP(16'hE4A3,4);
TASK_PP(16'hE4A4,4);
TASK_PP(16'hE4A5,4);
TASK_PP(16'hE4A6,4);
TASK_PP(16'hE4A7,4);
TASK_PP(16'hE4A8,4);
TASK_PP(16'hE4A9,4);
TASK_PP(16'hE4AA,4);
TASK_PP(16'hE4AB,4);
TASK_PP(16'hE4AC,4);
TASK_PP(16'hE4AD,4);
TASK_PP(16'hE4AE,4);
TASK_PP(16'hE4AF,4);
TASK_PP(16'hE4B0,4);
TASK_PP(16'hE4B1,4);
TASK_PP(16'hE4B2,4);
TASK_PP(16'hE4B3,4);
TASK_PP(16'hE4B4,4);
TASK_PP(16'hE4B5,4);
TASK_PP(16'hE4B6,4);
TASK_PP(16'hE4B7,4);
TASK_PP(16'hE4B8,4);
TASK_PP(16'hE4B9,4);
TASK_PP(16'hE4BA,4);
TASK_PP(16'hE4BB,4);
TASK_PP(16'hE4BC,4);
TASK_PP(16'hE4BD,4);
TASK_PP(16'hE4BE,4);
TASK_PP(16'hE4BF,4);
TASK_PP(16'hE4C0,4);
TASK_PP(16'hE4C1,4);
TASK_PP(16'hE4C2,4);
TASK_PP(16'hE4C3,4);
TASK_PP(16'hE4C4,4);
TASK_PP(16'hE4C5,4);
TASK_PP(16'hE4C6,4);
TASK_PP(16'hE4C7,4);
TASK_PP(16'hE4C8,4);
TASK_PP(16'hE4C9,4);
TASK_PP(16'hE4CA,4);
TASK_PP(16'hE4CB,4);
TASK_PP(16'hE4CC,4);
TASK_PP(16'hE4CD,4);
TASK_PP(16'hE4CE,4);
TASK_PP(16'hE4CF,4);
TASK_PP(16'hE4D0,4);
TASK_PP(16'hE4D1,4);
TASK_PP(16'hE4D2,4);
TASK_PP(16'hE4D3,4);
TASK_PP(16'hE4D4,4);
TASK_PP(16'hE4D5,4);
TASK_PP(16'hE4D6,4);
TASK_PP(16'hE4D7,4);
TASK_PP(16'hE4D8,4);
TASK_PP(16'hE4D9,4);
TASK_PP(16'hE4DA,4);
TASK_PP(16'hE4DB,4);
TASK_PP(16'hE4DC,4);
TASK_PP(16'hE4DD,4);
TASK_PP(16'hE4DE,4);
TASK_PP(16'hE4DF,4);
TASK_PP(16'hE4E0,4);
TASK_PP(16'hE4E1,4);
TASK_PP(16'hE4E2,4);
TASK_PP(16'hE4E3,4);
TASK_PP(16'hE4E4,4);
TASK_PP(16'hE4E5,4);
TASK_PP(16'hE4E6,4);
TASK_PP(16'hE4E7,4);
TASK_PP(16'hE4E8,4);
TASK_PP(16'hE4E9,4);
TASK_PP(16'hE4EA,4);
TASK_PP(16'hE4EB,4);
TASK_PP(16'hE4EC,4);
TASK_PP(16'hE4ED,4);
TASK_PP(16'hE4EE,4);
TASK_PP(16'hE4EF,4);
TASK_PP(16'hE4F0,4);
TASK_PP(16'hE4F1,4);
TASK_PP(16'hE4F2,4);
TASK_PP(16'hE4F3,4);
TASK_PP(16'hE4F4,4);
TASK_PP(16'hE4F5,4);
TASK_PP(16'hE4F6,4);
TASK_PP(16'hE4F7,4);
TASK_PP(16'hE4F8,4);
TASK_PP(16'hE4F9,4);
TASK_PP(16'hE4FA,4);
TASK_PP(16'hE4FB,4);
TASK_PP(16'hE4FC,4);
TASK_PP(16'hE4FD,4);
TASK_PP(16'hE4FE,4);
TASK_PP(16'hE4FF,4);
TASK_PP(16'hE500,4);
TASK_PP(16'hE501,4);
TASK_PP(16'hE502,4);
TASK_PP(16'hE503,4);
TASK_PP(16'hE504,4);
TASK_PP(16'hE505,4);
TASK_PP(16'hE506,4);
TASK_PP(16'hE507,4);
TASK_PP(16'hE508,4);
TASK_PP(16'hE509,4);
TASK_PP(16'hE50A,4);
TASK_PP(16'hE50B,4);
TASK_PP(16'hE50C,4);
TASK_PP(16'hE50D,4);
TASK_PP(16'hE50E,4);
TASK_PP(16'hE50F,4);
TASK_PP(16'hE510,4);
TASK_PP(16'hE511,4);
TASK_PP(16'hE512,4);
TASK_PP(16'hE513,4);
TASK_PP(16'hE514,4);
TASK_PP(16'hE515,4);
TASK_PP(16'hE516,4);
TASK_PP(16'hE517,4);
TASK_PP(16'hE518,4);
TASK_PP(16'hE519,4);
TASK_PP(16'hE51A,4);
TASK_PP(16'hE51B,4);
TASK_PP(16'hE51C,4);
TASK_PP(16'hE51D,4);
TASK_PP(16'hE51E,4);
TASK_PP(16'hE51F,4);
TASK_PP(16'hE520,4);
TASK_PP(16'hE521,4);
TASK_PP(16'hE522,4);
TASK_PP(16'hE523,4);
TASK_PP(16'hE524,4);
TASK_PP(16'hE525,4);
TASK_PP(16'hE526,4);
TASK_PP(16'hE527,4);
TASK_PP(16'hE528,4);
TASK_PP(16'hE529,4);
TASK_PP(16'hE52A,4);
TASK_PP(16'hE52B,4);
TASK_PP(16'hE52C,4);
TASK_PP(16'hE52D,4);
TASK_PP(16'hE52E,4);
TASK_PP(16'hE52F,4);
TASK_PP(16'hE530,4);
TASK_PP(16'hE531,4);
TASK_PP(16'hE532,4);
TASK_PP(16'hE533,4);
TASK_PP(16'hE534,4);
TASK_PP(16'hE535,4);
TASK_PP(16'hE536,4);
TASK_PP(16'hE537,4);
TASK_PP(16'hE538,4);
TASK_PP(16'hE539,4);
TASK_PP(16'hE53A,4);
TASK_PP(16'hE53B,4);
TASK_PP(16'hE53C,4);
TASK_PP(16'hE53D,4);
TASK_PP(16'hE53E,4);
TASK_PP(16'hE53F,4);
TASK_PP(16'hE540,4);
TASK_PP(16'hE541,4);
TASK_PP(16'hE542,4);
TASK_PP(16'hE543,4);
TASK_PP(16'hE544,4);
TASK_PP(16'hE545,4);
TASK_PP(16'hE546,4);
TASK_PP(16'hE547,4);
TASK_PP(16'hE548,4);
TASK_PP(16'hE549,4);
TASK_PP(16'hE54A,4);
TASK_PP(16'hE54B,4);
TASK_PP(16'hE54C,4);
TASK_PP(16'hE54D,4);
TASK_PP(16'hE54E,4);
TASK_PP(16'hE54F,4);
TASK_PP(16'hE550,4);
TASK_PP(16'hE551,4);
TASK_PP(16'hE552,4);
TASK_PP(16'hE553,4);
TASK_PP(16'hE554,4);
TASK_PP(16'hE555,4);
TASK_PP(16'hE556,4);
TASK_PP(16'hE557,4);
TASK_PP(16'hE558,4);
TASK_PP(16'hE559,4);
TASK_PP(16'hE55A,4);
TASK_PP(16'hE55B,4);
TASK_PP(16'hE55C,4);
TASK_PP(16'hE55D,4);
TASK_PP(16'hE55E,4);
TASK_PP(16'hE55F,4);
TASK_PP(16'hE560,4);
TASK_PP(16'hE561,4);
TASK_PP(16'hE562,4);
TASK_PP(16'hE563,4);
TASK_PP(16'hE564,4);
TASK_PP(16'hE565,4);
TASK_PP(16'hE566,4);
TASK_PP(16'hE567,4);
TASK_PP(16'hE568,4);
TASK_PP(16'hE569,4);
TASK_PP(16'hE56A,4);
TASK_PP(16'hE56B,4);
TASK_PP(16'hE56C,4);
TASK_PP(16'hE56D,4);
TASK_PP(16'hE56E,4);
TASK_PP(16'hE56F,4);
TASK_PP(16'hE570,4);
TASK_PP(16'hE571,4);
TASK_PP(16'hE572,4);
TASK_PP(16'hE573,4);
TASK_PP(16'hE574,4);
TASK_PP(16'hE575,4);
TASK_PP(16'hE576,4);
TASK_PP(16'hE577,4);
TASK_PP(16'hE578,4);
TASK_PP(16'hE579,4);
TASK_PP(16'hE57A,4);
TASK_PP(16'hE57B,4);
TASK_PP(16'hE57C,4);
TASK_PP(16'hE57D,4);
TASK_PP(16'hE57E,4);
TASK_PP(16'hE57F,4);
TASK_PP(16'hE580,4);
TASK_PP(16'hE581,4);
TASK_PP(16'hE582,4);
TASK_PP(16'hE583,4);
TASK_PP(16'hE584,4);
TASK_PP(16'hE585,4);
TASK_PP(16'hE586,4);
TASK_PP(16'hE587,4);
TASK_PP(16'hE588,4);
TASK_PP(16'hE589,4);
TASK_PP(16'hE58A,4);
TASK_PP(16'hE58B,4);
TASK_PP(16'hE58C,4);
TASK_PP(16'hE58D,4);
TASK_PP(16'hE58E,4);
TASK_PP(16'hE58F,4);
TASK_PP(16'hE590,4);
TASK_PP(16'hE591,4);
TASK_PP(16'hE592,4);
TASK_PP(16'hE593,4);
TASK_PP(16'hE594,4);
TASK_PP(16'hE595,4);
TASK_PP(16'hE596,4);
TASK_PP(16'hE597,4);
TASK_PP(16'hE598,4);
TASK_PP(16'hE599,4);
TASK_PP(16'hE59A,4);
TASK_PP(16'hE59B,4);
TASK_PP(16'hE59C,4);
TASK_PP(16'hE59D,4);
TASK_PP(16'hE59E,4);
TASK_PP(16'hE59F,4);
TASK_PP(16'hE5A0,4);
TASK_PP(16'hE5A1,4);
TASK_PP(16'hE5A2,4);
TASK_PP(16'hE5A3,4);
TASK_PP(16'hE5A4,4);
TASK_PP(16'hE5A5,4);
TASK_PP(16'hE5A6,4);
TASK_PP(16'hE5A7,4);
TASK_PP(16'hE5A8,4);
TASK_PP(16'hE5A9,4);
TASK_PP(16'hE5AA,4);
TASK_PP(16'hE5AB,4);
TASK_PP(16'hE5AC,4);
TASK_PP(16'hE5AD,4);
TASK_PP(16'hE5AE,4);
TASK_PP(16'hE5AF,4);
TASK_PP(16'hE5B0,4);
TASK_PP(16'hE5B1,4);
TASK_PP(16'hE5B2,4);
TASK_PP(16'hE5B3,4);
TASK_PP(16'hE5B4,4);
TASK_PP(16'hE5B5,4);
TASK_PP(16'hE5B6,4);
TASK_PP(16'hE5B7,4);
TASK_PP(16'hE5B8,4);
TASK_PP(16'hE5B9,4);
TASK_PP(16'hE5BA,4);
TASK_PP(16'hE5BB,4);
TASK_PP(16'hE5BC,4);
TASK_PP(16'hE5BD,4);
TASK_PP(16'hE5BE,4);
TASK_PP(16'hE5BF,4);
TASK_PP(16'hE5C0,4);
TASK_PP(16'hE5C1,4);
TASK_PP(16'hE5C2,4);
TASK_PP(16'hE5C3,4);
TASK_PP(16'hE5C4,4);
TASK_PP(16'hE5C5,4);
TASK_PP(16'hE5C6,4);
TASK_PP(16'hE5C7,4);
TASK_PP(16'hE5C8,4);
TASK_PP(16'hE5C9,4);
TASK_PP(16'hE5CA,4);
TASK_PP(16'hE5CB,4);
TASK_PP(16'hE5CC,4);
TASK_PP(16'hE5CD,4);
TASK_PP(16'hE5CE,4);
TASK_PP(16'hE5CF,4);
TASK_PP(16'hE5D0,4);
TASK_PP(16'hE5D1,4);
TASK_PP(16'hE5D2,4);
TASK_PP(16'hE5D3,4);
TASK_PP(16'hE5D4,4);
TASK_PP(16'hE5D5,4);
TASK_PP(16'hE5D6,4);
TASK_PP(16'hE5D7,4);
TASK_PP(16'hE5D8,4);
TASK_PP(16'hE5D9,4);
TASK_PP(16'hE5DA,4);
TASK_PP(16'hE5DB,4);
TASK_PP(16'hE5DC,4);
TASK_PP(16'hE5DD,4);
TASK_PP(16'hE5DE,4);
TASK_PP(16'hE5DF,4);
TASK_PP(16'hE5E0,4);
TASK_PP(16'hE5E1,4);
TASK_PP(16'hE5E2,4);
TASK_PP(16'hE5E3,4);
TASK_PP(16'hE5E4,4);
TASK_PP(16'hE5E5,4);
TASK_PP(16'hE5E6,4);
TASK_PP(16'hE5E7,4);
TASK_PP(16'hE5E8,4);
TASK_PP(16'hE5E9,4);
TASK_PP(16'hE5EA,4);
TASK_PP(16'hE5EB,4);
TASK_PP(16'hE5EC,4);
TASK_PP(16'hE5ED,4);
TASK_PP(16'hE5EE,4);
TASK_PP(16'hE5EF,4);
TASK_PP(16'hE5F0,4);
TASK_PP(16'hE5F1,4);
TASK_PP(16'hE5F2,4);
TASK_PP(16'hE5F3,4);
TASK_PP(16'hE5F4,4);
TASK_PP(16'hE5F5,4);
TASK_PP(16'hE5F6,4);
TASK_PP(16'hE5F7,4);
TASK_PP(16'hE5F8,4);
TASK_PP(16'hE5F9,4);
TASK_PP(16'hE5FA,4);
TASK_PP(16'hE5FB,4);
TASK_PP(16'hE5FC,4);
TASK_PP(16'hE5FD,4);
TASK_PP(16'hE5FE,4);
TASK_PP(16'hE5FF,4);
TASK_PP(16'hE600,4);
TASK_PP(16'hE601,4);
TASK_PP(16'hE602,4);
TASK_PP(16'hE603,4);
TASK_PP(16'hE604,4);
TASK_PP(16'hE605,4);
TASK_PP(16'hE606,4);
TASK_PP(16'hE607,4);
TASK_PP(16'hE608,4);
TASK_PP(16'hE609,4);
TASK_PP(16'hE60A,4);
TASK_PP(16'hE60B,4);
TASK_PP(16'hE60C,4);
TASK_PP(16'hE60D,4);
TASK_PP(16'hE60E,4);
TASK_PP(16'hE60F,4);
TASK_PP(16'hE610,4);
TASK_PP(16'hE611,4);
TASK_PP(16'hE612,4);
TASK_PP(16'hE613,4);
TASK_PP(16'hE614,4);
TASK_PP(16'hE615,4);
TASK_PP(16'hE616,4);
TASK_PP(16'hE617,4);
TASK_PP(16'hE618,4);
TASK_PP(16'hE619,4);
TASK_PP(16'hE61A,4);
TASK_PP(16'hE61B,4);
TASK_PP(16'hE61C,4);
TASK_PP(16'hE61D,4);
TASK_PP(16'hE61E,4);
TASK_PP(16'hE61F,4);
TASK_PP(16'hE620,4);
TASK_PP(16'hE621,4);
TASK_PP(16'hE622,4);
TASK_PP(16'hE623,4);
TASK_PP(16'hE624,4);
TASK_PP(16'hE625,4);
TASK_PP(16'hE626,4);
TASK_PP(16'hE627,4);
TASK_PP(16'hE628,4);
TASK_PP(16'hE629,4);
TASK_PP(16'hE62A,4);
TASK_PP(16'hE62B,4);
TASK_PP(16'hE62C,4);
TASK_PP(16'hE62D,4);
TASK_PP(16'hE62E,4);
TASK_PP(16'hE62F,4);
TASK_PP(16'hE630,4);
TASK_PP(16'hE631,4);
TASK_PP(16'hE632,4);
TASK_PP(16'hE633,4);
TASK_PP(16'hE634,4);
TASK_PP(16'hE635,4);
TASK_PP(16'hE636,4);
TASK_PP(16'hE637,4);
TASK_PP(16'hE638,4);
TASK_PP(16'hE639,4);
TASK_PP(16'hE63A,4);
TASK_PP(16'hE63B,4);
TASK_PP(16'hE63C,4);
TASK_PP(16'hE63D,4);
TASK_PP(16'hE63E,4);
TASK_PP(16'hE63F,4);
TASK_PP(16'hE640,4);
TASK_PP(16'hE641,4);
TASK_PP(16'hE642,4);
TASK_PP(16'hE643,4);
TASK_PP(16'hE644,4);
TASK_PP(16'hE645,4);
TASK_PP(16'hE646,4);
TASK_PP(16'hE647,4);
TASK_PP(16'hE648,4);
TASK_PP(16'hE649,4);
TASK_PP(16'hE64A,4);
TASK_PP(16'hE64B,4);
TASK_PP(16'hE64C,4);
TASK_PP(16'hE64D,4);
TASK_PP(16'hE64E,4);
TASK_PP(16'hE64F,4);
TASK_PP(16'hE650,4);
TASK_PP(16'hE651,4);
TASK_PP(16'hE652,4);
TASK_PP(16'hE653,4);
TASK_PP(16'hE654,4);
TASK_PP(16'hE655,4);
TASK_PP(16'hE656,4);
TASK_PP(16'hE657,4);
TASK_PP(16'hE658,4);
TASK_PP(16'hE659,4);
TASK_PP(16'hE65A,4);
TASK_PP(16'hE65B,4);
TASK_PP(16'hE65C,4);
TASK_PP(16'hE65D,4);
TASK_PP(16'hE65E,4);
TASK_PP(16'hE65F,4);
TASK_PP(16'hE660,4);
TASK_PP(16'hE661,4);
TASK_PP(16'hE662,4);
TASK_PP(16'hE663,4);
TASK_PP(16'hE664,4);
TASK_PP(16'hE665,4);
TASK_PP(16'hE666,4);
TASK_PP(16'hE667,4);
TASK_PP(16'hE668,4);
TASK_PP(16'hE669,4);
TASK_PP(16'hE66A,4);
TASK_PP(16'hE66B,4);
TASK_PP(16'hE66C,4);
TASK_PP(16'hE66D,4);
TASK_PP(16'hE66E,4);
TASK_PP(16'hE66F,4);
TASK_PP(16'hE670,4);
TASK_PP(16'hE671,4);
TASK_PP(16'hE672,4);
TASK_PP(16'hE673,4);
TASK_PP(16'hE674,4);
TASK_PP(16'hE675,4);
TASK_PP(16'hE676,4);
TASK_PP(16'hE677,4);
TASK_PP(16'hE678,4);
TASK_PP(16'hE679,4);
TASK_PP(16'hE67A,4);
TASK_PP(16'hE67B,4);
TASK_PP(16'hE67C,4);
TASK_PP(16'hE67D,4);
TASK_PP(16'hE67E,4);
TASK_PP(16'hE67F,4);
TASK_PP(16'hE680,4);
TASK_PP(16'hE681,4);
TASK_PP(16'hE682,4);
TASK_PP(16'hE683,4);
TASK_PP(16'hE684,4);
TASK_PP(16'hE685,4);
TASK_PP(16'hE686,4);
TASK_PP(16'hE687,4);
TASK_PP(16'hE688,4);
TASK_PP(16'hE689,4);
TASK_PP(16'hE68A,4);
TASK_PP(16'hE68B,4);
TASK_PP(16'hE68C,4);
TASK_PP(16'hE68D,4);
TASK_PP(16'hE68E,4);
TASK_PP(16'hE68F,4);
TASK_PP(16'hE690,4);
TASK_PP(16'hE691,4);
TASK_PP(16'hE692,4);
TASK_PP(16'hE693,4);
TASK_PP(16'hE694,4);
TASK_PP(16'hE695,4);
TASK_PP(16'hE696,4);
TASK_PP(16'hE697,4);
TASK_PP(16'hE698,4);
TASK_PP(16'hE699,4);
TASK_PP(16'hE69A,4);
TASK_PP(16'hE69B,4);
TASK_PP(16'hE69C,4);
TASK_PP(16'hE69D,4);
TASK_PP(16'hE69E,4);
TASK_PP(16'hE69F,4);
TASK_PP(16'hE6A0,4);
TASK_PP(16'hE6A1,4);
TASK_PP(16'hE6A2,4);
TASK_PP(16'hE6A3,4);
TASK_PP(16'hE6A4,4);
TASK_PP(16'hE6A5,4);
TASK_PP(16'hE6A6,4);
TASK_PP(16'hE6A7,4);
TASK_PP(16'hE6A8,4);
TASK_PP(16'hE6A9,4);
TASK_PP(16'hE6AA,4);
TASK_PP(16'hE6AB,4);
TASK_PP(16'hE6AC,4);
TASK_PP(16'hE6AD,4);
TASK_PP(16'hE6AE,4);
TASK_PP(16'hE6AF,4);
TASK_PP(16'hE6B0,4);
TASK_PP(16'hE6B1,4);
TASK_PP(16'hE6B2,4);
TASK_PP(16'hE6B3,4);
TASK_PP(16'hE6B4,4);
TASK_PP(16'hE6B5,4);
TASK_PP(16'hE6B6,4);
TASK_PP(16'hE6B7,4);
TASK_PP(16'hE6B8,4);
TASK_PP(16'hE6B9,4);
TASK_PP(16'hE6BA,4);
TASK_PP(16'hE6BB,4);
TASK_PP(16'hE6BC,4);
TASK_PP(16'hE6BD,4);
TASK_PP(16'hE6BE,4);
TASK_PP(16'hE6BF,4);
TASK_PP(16'hE6C0,4);
TASK_PP(16'hE6C1,4);
TASK_PP(16'hE6C2,4);
TASK_PP(16'hE6C3,4);
TASK_PP(16'hE6C4,4);
TASK_PP(16'hE6C5,4);
TASK_PP(16'hE6C6,4);
TASK_PP(16'hE6C7,4);
TASK_PP(16'hE6C8,4);
TASK_PP(16'hE6C9,4);
TASK_PP(16'hE6CA,4);
TASK_PP(16'hE6CB,4);
TASK_PP(16'hE6CC,4);
TASK_PP(16'hE6CD,4);
TASK_PP(16'hE6CE,4);
TASK_PP(16'hE6CF,4);
TASK_PP(16'hE6D0,4);
TASK_PP(16'hE6D1,4);
TASK_PP(16'hE6D2,4);
TASK_PP(16'hE6D3,4);
TASK_PP(16'hE6D4,4);
TASK_PP(16'hE6D5,4);
TASK_PP(16'hE6D6,4);
TASK_PP(16'hE6D7,4);
TASK_PP(16'hE6D8,4);
TASK_PP(16'hE6D9,4);
TASK_PP(16'hE6DA,4);
TASK_PP(16'hE6DB,4);
TASK_PP(16'hE6DC,4);
TASK_PP(16'hE6DD,4);
TASK_PP(16'hE6DE,4);
TASK_PP(16'hE6DF,4);
TASK_PP(16'hE6E0,4);
TASK_PP(16'hE6E1,4);
TASK_PP(16'hE6E2,4);
TASK_PP(16'hE6E3,4);
TASK_PP(16'hE6E4,4);
TASK_PP(16'hE6E5,4);
TASK_PP(16'hE6E6,4);
TASK_PP(16'hE6E7,4);
TASK_PP(16'hE6E8,4);
TASK_PP(16'hE6E9,4);
TASK_PP(16'hE6EA,4);
TASK_PP(16'hE6EB,4);
TASK_PP(16'hE6EC,4);
TASK_PP(16'hE6ED,4);
TASK_PP(16'hE6EE,4);
TASK_PP(16'hE6EF,4);
TASK_PP(16'hE6F0,4);
TASK_PP(16'hE6F1,4);
TASK_PP(16'hE6F2,4);
TASK_PP(16'hE6F3,4);
TASK_PP(16'hE6F4,4);
TASK_PP(16'hE6F5,4);
TASK_PP(16'hE6F6,4);
TASK_PP(16'hE6F7,4);
TASK_PP(16'hE6F8,4);
TASK_PP(16'hE6F9,4);
TASK_PP(16'hE6FA,4);
TASK_PP(16'hE6FB,4);
TASK_PP(16'hE6FC,4);
TASK_PP(16'hE6FD,4);
TASK_PP(16'hE6FE,4);
TASK_PP(16'hE6FF,4);
TASK_PP(16'hE700,4);
TASK_PP(16'hE701,4);
TASK_PP(16'hE702,4);
TASK_PP(16'hE703,4);
TASK_PP(16'hE704,4);
TASK_PP(16'hE705,4);
TASK_PP(16'hE706,4);
TASK_PP(16'hE707,4);
TASK_PP(16'hE708,4);
TASK_PP(16'hE709,4);
TASK_PP(16'hE70A,4);
TASK_PP(16'hE70B,4);
TASK_PP(16'hE70C,4);
TASK_PP(16'hE70D,4);
TASK_PP(16'hE70E,4);
TASK_PP(16'hE70F,4);
TASK_PP(16'hE710,4);
TASK_PP(16'hE711,4);
TASK_PP(16'hE712,4);
TASK_PP(16'hE713,4);
TASK_PP(16'hE714,4);
TASK_PP(16'hE715,4);
TASK_PP(16'hE716,4);
TASK_PP(16'hE717,4);
TASK_PP(16'hE718,4);
TASK_PP(16'hE719,4);
TASK_PP(16'hE71A,4);
TASK_PP(16'hE71B,4);
TASK_PP(16'hE71C,4);
TASK_PP(16'hE71D,4);
TASK_PP(16'hE71E,4);
TASK_PP(16'hE71F,4);
TASK_PP(16'hE720,4);
TASK_PP(16'hE721,4);
TASK_PP(16'hE722,4);
TASK_PP(16'hE723,4);
TASK_PP(16'hE724,4);
TASK_PP(16'hE725,4);
TASK_PP(16'hE726,4);
TASK_PP(16'hE727,4);
TASK_PP(16'hE728,4);
TASK_PP(16'hE729,4);
TASK_PP(16'hE72A,4);
TASK_PP(16'hE72B,4);
TASK_PP(16'hE72C,4);
TASK_PP(16'hE72D,4);
TASK_PP(16'hE72E,4);
TASK_PP(16'hE72F,4);
TASK_PP(16'hE730,4);
TASK_PP(16'hE731,4);
TASK_PP(16'hE732,4);
TASK_PP(16'hE733,4);
TASK_PP(16'hE734,4);
TASK_PP(16'hE735,4);
TASK_PP(16'hE736,4);
TASK_PP(16'hE737,4);
TASK_PP(16'hE738,4);
TASK_PP(16'hE739,4);
TASK_PP(16'hE73A,4);
TASK_PP(16'hE73B,4);
TASK_PP(16'hE73C,4);
TASK_PP(16'hE73D,4);
TASK_PP(16'hE73E,4);
TASK_PP(16'hE73F,4);
TASK_PP(16'hE740,4);
TASK_PP(16'hE741,4);
TASK_PP(16'hE742,4);
TASK_PP(16'hE743,4);
TASK_PP(16'hE744,4);
TASK_PP(16'hE745,4);
TASK_PP(16'hE746,4);
TASK_PP(16'hE747,4);
TASK_PP(16'hE748,4);
TASK_PP(16'hE749,4);
TASK_PP(16'hE74A,4);
TASK_PP(16'hE74B,4);
TASK_PP(16'hE74C,4);
TASK_PP(16'hE74D,4);
TASK_PP(16'hE74E,4);
TASK_PP(16'hE74F,4);
TASK_PP(16'hE750,4);
TASK_PP(16'hE751,4);
TASK_PP(16'hE752,4);
TASK_PP(16'hE753,4);
TASK_PP(16'hE754,4);
TASK_PP(16'hE755,4);
TASK_PP(16'hE756,4);
TASK_PP(16'hE757,4);
TASK_PP(16'hE758,4);
TASK_PP(16'hE759,4);
TASK_PP(16'hE75A,4);
TASK_PP(16'hE75B,4);
TASK_PP(16'hE75C,4);
TASK_PP(16'hE75D,4);
TASK_PP(16'hE75E,4);
TASK_PP(16'hE75F,4);
TASK_PP(16'hE760,4);
TASK_PP(16'hE761,4);
TASK_PP(16'hE762,4);
TASK_PP(16'hE763,4);
TASK_PP(16'hE764,4);
TASK_PP(16'hE765,4);
TASK_PP(16'hE766,4);
TASK_PP(16'hE767,4);
TASK_PP(16'hE768,4);
TASK_PP(16'hE769,4);
TASK_PP(16'hE76A,4);
TASK_PP(16'hE76B,4);
TASK_PP(16'hE76C,4);
TASK_PP(16'hE76D,4);
TASK_PP(16'hE76E,4);
TASK_PP(16'hE76F,4);
TASK_PP(16'hE770,4);
TASK_PP(16'hE771,4);
TASK_PP(16'hE772,4);
TASK_PP(16'hE773,4);
TASK_PP(16'hE774,4);
TASK_PP(16'hE775,4);
TASK_PP(16'hE776,4);
TASK_PP(16'hE777,4);
TASK_PP(16'hE778,4);
TASK_PP(16'hE779,4);
TASK_PP(16'hE77A,4);
TASK_PP(16'hE77B,4);
TASK_PP(16'hE77C,4);
TASK_PP(16'hE77D,4);
TASK_PP(16'hE77E,4);
TASK_PP(16'hE77F,4);
TASK_PP(16'hE780,4);
TASK_PP(16'hE781,4);
TASK_PP(16'hE782,4);
TASK_PP(16'hE783,4);
TASK_PP(16'hE784,4);
TASK_PP(16'hE785,4);
TASK_PP(16'hE786,4);
TASK_PP(16'hE787,4);
TASK_PP(16'hE788,4);
TASK_PP(16'hE789,4);
TASK_PP(16'hE78A,4);
TASK_PP(16'hE78B,4);
TASK_PP(16'hE78C,4);
TASK_PP(16'hE78D,4);
TASK_PP(16'hE78E,4);
TASK_PP(16'hE78F,4);
TASK_PP(16'hE790,4);
TASK_PP(16'hE791,4);
TASK_PP(16'hE792,4);
TASK_PP(16'hE793,4);
TASK_PP(16'hE794,4);
TASK_PP(16'hE795,4);
TASK_PP(16'hE796,4);
TASK_PP(16'hE797,4);
TASK_PP(16'hE798,4);
TASK_PP(16'hE799,4);
TASK_PP(16'hE79A,4);
TASK_PP(16'hE79B,4);
TASK_PP(16'hE79C,4);
TASK_PP(16'hE79D,4);
TASK_PP(16'hE79E,4);
TASK_PP(16'hE79F,4);
TASK_PP(16'hE7A0,4);
TASK_PP(16'hE7A1,4);
TASK_PP(16'hE7A2,4);
TASK_PP(16'hE7A3,4);
TASK_PP(16'hE7A4,4);
TASK_PP(16'hE7A5,4);
TASK_PP(16'hE7A6,4);
TASK_PP(16'hE7A7,4);
TASK_PP(16'hE7A8,4);
TASK_PP(16'hE7A9,4);
TASK_PP(16'hE7AA,4);
TASK_PP(16'hE7AB,4);
TASK_PP(16'hE7AC,4);
TASK_PP(16'hE7AD,4);
TASK_PP(16'hE7AE,4);
TASK_PP(16'hE7AF,4);
TASK_PP(16'hE7B0,4);
TASK_PP(16'hE7B1,4);
TASK_PP(16'hE7B2,4);
TASK_PP(16'hE7B3,4);
TASK_PP(16'hE7B4,4);
TASK_PP(16'hE7B5,4);
TASK_PP(16'hE7B6,4);
TASK_PP(16'hE7B7,4);
TASK_PP(16'hE7B8,4);
TASK_PP(16'hE7B9,4);
TASK_PP(16'hE7BA,4);
TASK_PP(16'hE7BB,4);
TASK_PP(16'hE7BC,4);
TASK_PP(16'hE7BD,4);
TASK_PP(16'hE7BE,4);
TASK_PP(16'hE7BF,4);
TASK_PP(16'hE7C0,4);
TASK_PP(16'hE7C1,4);
TASK_PP(16'hE7C2,4);
TASK_PP(16'hE7C3,4);
TASK_PP(16'hE7C4,4);
TASK_PP(16'hE7C5,4);
TASK_PP(16'hE7C6,4);
TASK_PP(16'hE7C7,4);
TASK_PP(16'hE7C8,4);
TASK_PP(16'hE7C9,4);
TASK_PP(16'hE7CA,4);
TASK_PP(16'hE7CB,4);
TASK_PP(16'hE7CC,4);
TASK_PP(16'hE7CD,4);
TASK_PP(16'hE7CE,4);
TASK_PP(16'hE7CF,4);
TASK_PP(16'hE7D0,4);
TASK_PP(16'hE7D1,4);
TASK_PP(16'hE7D2,4);
TASK_PP(16'hE7D3,4);
TASK_PP(16'hE7D4,4);
TASK_PP(16'hE7D5,4);
TASK_PP(16'hE7D6,4);
TASK_PP(16'hE7D7,4);
TASK_PP(16'hE7D8,4);
TASK_PP(16'hE7D9,4);
TASK_PP(16'hE7DA,4);
TASK_PP(16'hE7DB,4);
TASK_PP(16'hE7DC,4);
TASK_PP(16'hE7DD,4);
TASK_PP(16'hE7DE,4);
TASK_PP(16'hE7DF,4);
TASK_PP(16'hE7E0,4);
TASK_PP(16'hE7E1,4);
TASK_PP(16'hE7E2,4);
TASK_PP(16'hE7E3,4);
TASK_PP(16'hE7E4,4);
TASK_PP(16'hE7E5,4);
TASK_PP(16'hE7E6,4);
TASK_PP(16'hE7E7,4);
TASK_PP(16'hE7E8,4);
TASK_PP(16'hE7E9,4);
TASK_PP(16'hE7EA,4);
TASK_PP(16'hE7EB,4);
TASK_PP(16'hE7EC,4);
TASK_PP(16'hE7ED,4);
TASK_PP(16'hE7EE,4);
TASK_PP(16'hE7EF,4);
TASK_PP(16'hE7F0,4);
TASK_PP(16'hE7F1,4);
TASK_PP(16'hE7F2,4);
TASK_PP(16'hE7F3,4);
TASK_PP(16'hE7F4,4);
TASK_PP(16'hE7F5,4);
TASK_PP(16'hE7F6,4);
TASK_PP(16'hE7F7,4);
TASK_PP(16'hE7F8,4);
TASK_PP(16'hE7F9,4);
TASK_PP(16'hE7FA,4);
TASK_PP(16'hE7FB,4);
TASK_PP(16'hE7FC,4);
TASK_PP(16'hE7FD,4);
TASK_PP(16'hE7FE,4);
TASK_PP(16'hE7FF,4);
TASK_PP(16'hE800,4);
TASK_PP(16'hE801,4);
TASK_PP(16'hE802,4);
TASK_PP(16'hE803,4);
TASK_PP(16'hE804,4);
TASK_PP(16'hE805,4);
TASK_PP(16'hE806,4);
TASK_PP(16'hE807,4);
TASK_PP(16'hE808,4);
TASK_PP(16'hE809,4);
TASK_PP(16'hE80A,4);
TASK_PP(16'hE80B,4);
TASK_PP(16'hE80C,4);
TASK_PP(16'hE80D,4);
TASK_PP(16'hE80E,4);
TASK_PP(16'hE80F,4);
TASK_PP(16'hE810,4);
TASK_PP(16'hE811,4);
TASK_PP(16'hE812,4);
TASK_PP(16'hE813,4);
TASK_PP(16'hE814,4);
TASK_PP(16'hE815,4);
TASK_PP(16'hE816,4);
TASK_PP(16'hE817,4);
TASK_PP(16'hE818,4);
TASK_PP(16'hE819,4);
TASK_PP(16'hE81A,4);
TASK_PP(16'hE81B,4);
TASK_PP(16'hE81C,4);
TASK_PP(16'hE81D,4);
TASK_PP(16'hE81E,4);
TASK_PP(16'hE81F,4);
TASK_PP(16'hE820,4);
TASK_PP(16'hE821,4);
TASK_PP(16'hE822,4);
TASK_PP(16'hE823,4);
TASK_PP(16'hE824,4);
TASK_PP(16'hE825,4);
TASK_PP(16'hE826,4);
TASK_PP(16'hE827,4);
TASK_PP(16'hE828,4);
TASK_PP(16'hE829,4);
TASK_PP(16'hE82A,4);
TASK_PP(16'hE82B,4);
TASK_PP(16'hE82C,4);
TASK_PP(16'hE82D,4);
TASK_PP(16'hE82E,4);
TASK_PP(16'hE82F,4);
TASK_PP(16'hE830,4);
TASK_PP(16'hE831,4);
TASK_PP(16'hE832,4);
TASK_PP(16'hE833,4);
TASK_PP(16'hE834,4);
TASK_PP(16'hE835,4);
TASK_PP(16'hE836,4);
TASK_PP(16'hE837,4);
TASK_PP(16'hE838,4);
TASK_PP(16'hE839,4);
TASK_PP(16'hE83A,4);
TASK_PP(16'hE83B,4);
TASK_PP(16'hE83C,4);
TASK_PP(16'hE83D,4);
TASK_PP(16'hE83E,4);
TASK_PP(16'hE83F,4);
TASK_PP(16'hE840,4);
TASK_PP(16'hE841,4);
TASK_PP(16'hE842,4);
TASK_PP(16'hE843,4);
TASK_PP(16'hE844,4);
TASK_PP(16'hE845,4);
TASK_PP(16'hE846,4);
TASK_PP(16'hE847,4);
TASK_PP(16'hE848,4);
TASK_PP(16'hE849,4);
TASK_PP(16'hE84A,4);
TASK_PP(16'hE84B,4);
TASK_PP(16'hE84C,4);
TASK_PP(16'hE84D,4);
TASK_PP(16'hE84E,4);
TASK_PP(16'hE84F,4);
TASK_PP(16'hE850,4);
TASK_PP(16'hE851,4);
TASK_PP(16'hE852,4);
TASK_PP(16'hE853,4);
TASK_PP(16'hE854,4);
TASK_PP(16'hE855,4);
TASK_PP(16'hE856,4);
TASK_PP(16'hE857,4);
TASK_PP(16'hE858,4);
TASK_PP(16'hE859,4);
TASK_PP(16'hE85A,4);
TASK_PP(16'hE85B,4);
TASK_PP(16'hE85C,4);
TASK_PP(16'hE85D,4);
TASK_PP(16'hE85E,4);
TASK_PP(16'hE85F,4);
TASK_PP(16'hE860,4);
TASK_PP(16'hE861,4);
TASK_PP(16'hE862,4);
TASK_PP(16'hE863,4);
TASK_PP(16'hE864,4);
TASK_PP(16'hE865,4);
TASK_PP(16'hE866,4);
TASK_PP(16'hE867,4);
TASK_PP(16'hE868,4);
TASK_PP(16'hE869,4);
TASK_PP(16'hE86A,4);
TASK_PP(16'hE86B,4);
TASK_PP(16'hE86C,4);
TASK_PP(16'hE86D,4);
TASK_PP(16'hE86E,4);
TASK_PP(16'hE86F,4);
TASK_PP(16'hE870,4);
TASK_PP(16'hE871,4);
TASK_PP(16'hE872,4);
TASK_PP(16'hE873,4);
TASK_PP(16'hE874,4);
TASK_PP(16'hE875,4);
TASK_PP(16'hE876,4);
TASK_PP(16'hE877,4);
TASK_PP(16'hE878,4);
TASK_PP(16'hE879,4);
TASK_PP(16'hE87A,4);
TASK_PP(16'hE87B,4);
TASK_PP(16'hE87C,4);
TASK_PP(16'hE87D,4);
TASK_PP(16'hE87E,4);
TASK_PP(16'hE87F,4);
TASK_PP(16'hE880,4);
TASK_PP(16'hE881,4);
TASK_PP(16'hE882,4);
TASK_PP(16'hE883,4);
TASK_PP(16'hE884,4);
TASK_PP(16'hE885,4);
TASK_PP(16'hE886,4);
TASK_PP(16'hE887,4);
TASK_PP(16'hE888,4);
TASK_PP(16'hE889,4);
TASK_PP(16'hE88A,4);
TASK_PP(16'hE88B,4);
TASK_PP(16'hE88C,4);
TASK_PP(16'hE88D,4);
TASK_PP(16'hE88E,4);
TASK_PP(16'hE88F,4);
TASK_PP(16'hE890,4);
TASK_PP(16'hE891,4);
TASK_PP(16'hE892,4);
TASK_PP(16'hE893,4);
TASK_PP(16'hE894,4);
TASK_PP(16'hE895,4);
TASK_PP(16'hE896,4);
TASK_PP(16'hE897,4);
TASK_PP(16'hE898,4);
TASK_PP(16'hE899,4);
TASK_PP(16'hE89A,4);
TASK_PP(16'hE89B,4);
TASK_PP(16'hE89C,4);
TASK_PP(16'hE89D,4);
TASK_PP(16'hE89E,4);
TASK_PP(16'hE89F,4);
TASK_PP(16'hE8A0,4);
TASK_PP(16'hE8A1,4);
TASK_PP(16'hE8A2,4);
TASK_PP(16'hE8A3,4);
TASK_PP(16'hE8A4,4);
TASK_PP(16'hE8A5,4);
TASK_PP(16'hE8A6,4);
TASK_PP(16'hE8A7,4);
TASK_PP(16'hE8A8,4);
TASK_PP(16'hE8A9,4);
TASK_PP(16'hE8AA,4);
TASK_PP(16'hE8AB,4);
TASK_PP(16'hE8AC,4);
TASK_PP(16'hE8AD,4);
TASK_PP(16'hE8AE,4);
TASK_PP(16'hE8AF,4);
TASK_PP(16'hE8B0,4);
TASK_PP(16'hE8B1,4);
TASK_PP(16'hE8B2,4);
TASK_PP(16'hE8B3,4);
TASK_PP(16'hE8B4,4);
TASK_PP(16'hE8B5,4);
TASK_PP(16'hE8B6,4);
TASK_PP(16'hE8B7,4);
TASK_PP(16'hE8B8,4);
TASK_PP(16'hE8B9,4);
TASK_PP(16'hE8BA,4);
TASK_PP(16'hE8BB,4);
TASK_PP(16'hE8BC,4);
TASK_PP(16'hE8BD,4);
TASK_PP(16'hE8BE,4);
TASK_PP(16'hE8BF,4);
TASK_PP(16'hE8C0,4);
TASK_PP(16'hE8C1,4);
TASK_PP(16'hE8C2,4);
TASK_PP(16'hE8C3,4);
TASK_PP(16'hE8C4,4);
TASK_PP(16'hE8C5,4);
TASK_PP(16'hE8C6,4);
TASK_PP(16'hE8C7,4);
TASK_PP(16'hE8C8,4);
TASK_PP(16'hE8C9,4);
TASK_PP(16'hE8CA,4);
TASK_PP(16'hE8CB,4);
TASK_PP(16'hE8CC,4);
TASK_PP(16'hE8CD,4);
TASK_PP(16'hE8CE,4);
TASK_PP(16'hE8CF,4);
TASK_PP(16'hE8D0,4);
TASK_PP(16'hE8D1,4);
TASK_PP(16'hE8D2,4);
TASK_PP(16'hE8D3,4);
TASK_PP(16'hE8D4,4);
TASK_PP(16'hE8D5,4);
TASK_PP(16'hE8D6,4);
TASK_PP(16'hE8D7,4);
TASK_PP(16'hE8D8,4);
TASK_PP(16'hE8D9,4);
TASK_PP(16'hE8DA,4);
TASK_PP(16'hE8DB,4);
TASK_PP(16'hE8DC,4);
TASK_PP(16'hE8DD,4);
TASK_PP(16'hE8DE,4);
TASK_PP(16'hE8DF,4);
TASK_PP(16'hE8E0,4);
TASK_PP(16'hE8E1,4);
TASK_PP(16'hE8E2,4);
TASK_PP(16'hE8E3,4);
TASK_PP(16'hE8E4,4);
TASK_PP(16'hE8E5,4);
TASK_PP(16'hE8E6,4);
TASK_PP(16'hE8E7,4);
TASK_PP(16'hE8E8,4);
TASK_PP(16'hE8E9,4);
TASK_PP(16'hE8EA,4);
TASK_PP(16'hE8EB,4);
TASK_PP(16'hE8EC,4);
TASK_PP(16'hE8ED,4);
TASK_PP(16'hE8EE,4);
TASK_PP(16'hE8EF,4);
TASK_PP(16'hE8F0,4);
TASK_PP(16'hE8F1,4);
TASK_PP(16'hE8F2,4);
TASK_PP(16'hE8F3,4);
TASK_PP(16'hE8F4,4);
TASK_PP(16'hE8F5,4);
TASK_PP(16'hE8F6,4);
TASK_PP(16'hE8F7,4);
TASK_PP(16'hE8F8,4);
TASK_PP(16'hE8F9,4);
TASK_PP(16'hE8FA,4);
TASK_PP(16'hE8FB,4);
TASK_PP(16'hE8FC,4);
TASK_PP(16'hE8FD,4);
TASK_PP(16'hE8FE,4);
TASK_PP(16'hE8FF,4);
TASK_PP(16'hE900,4);
TASK_PP(16'hE901,4);
TASK_PP(16'hE902,4);
TASK_PP(16'hE903,4);
TASK_PP(16'hE904,4);
TASK_PP(16'hE905,4);
TASK_PP(16'hE906,4);
TASK_PP(16'hE907,4);
TASK_PP(16'hE908,4);
TASK_PP(16'hE909,4);
TASK_PP(16'hE90A,4);
TASK_PP(16'hE90B,4);
TASK_PP(16'hE90C,4);
TASK_PP(16'hE90D,4);
TASK_PP(16'hE90E,4);
TASK_PP(16'hE90F,4);
TASK_PP(16'hE910,4);
TASK_PP(16'hE911,4);
TASK_PP(16'hE912,4);
TASK_PP(16'hE913,4);
TASK_PP(16'hE914,4);
TASK_PP(16'hE915,4);
TASK_PP(16'hE916,4);
TASK_PP(16'hE917,4);
TASK_PP(16'hE918,4);
TASK_PP(16'hE919,4);
TASK_PP(16'hE91A,4);
TASK_PP(16'hE91B,4);
TASK_PP(16'hE91C,4);
TASK_PP(16'hE91D,4);
TASK_PP(16'hE91E,4);
TASK_PP(16'hE91F,4);
TASK_PP(16'hE920,4);
TASK_PP(16'hE921,4);
TASK_PP(16'hE922,4);
TASK_PP(16'hE923,4);
TASK_PP(16'hE924,4);
TASK_PP(16'hE925,4);
TASK_PP(16'hE926,4);
TASK_PP(16'hE927,4);
TASK_PP(16'hE928,4);
TASK_PP(16'hE929,4);
TASK_PP(16'hE92A,4);
TASK_PP(16'hE92B,4);
TASK_PP(16'hE92C,4);
TASK_PP(16'hE92D,4);
TASK_PP(16'hE92E,4);
TASK_PP(16'hE92F,4);
TASK_PP(16'hE930,4);
TASK_PP(16'hE931,4);
TASK_PP(16'hE932,4);
TASK_PP(16'hE933,4);
TASK_PP(16'hE934,4);
TASK_PP(16'hE935,4);
TASK_PP(16'hE936,4);
TASK_PP(16'hE937,4);
TASK_PP(16'hE938,4);
TASK_PP(16'hE939,4);
TASK_PP(16'hE93A,4);
TASK_PP(16'hE93B,4);
TASK_PP(16'hE93C,4);
TASK_PP(16'hE93D,4);
TASK_PP(16'hE93E,4);
TASK_PP(16'hE93F,4);
TASK_PP(16'hE940,4);
TASK_PP(16'hE941,4);
TASK_PP(16'hE942,4);
TASK_PP(16'hE943,4);
TASK_PP(16'hE944,4);
TASK_PP(16'hE945,4);
TASK_PP(16'hE946,4);
TASK_PP(16'hE947,4);
TASK_PP(16'hE948,4);
TASK_PP(16'hE949,4);
TASK_PP(16'hE94A,4);
TASK_PP(16'hE94B,4);
TASK_PP(16'hE94C,4);
TASK_PP(16'hE94D,4);
TASK_PP(16'hE94E,4);
TASK_PP(16'hE94F,4);
TASK_PP(16'hE950,4);
TASK_PP(16'hE951,4);
TASK_PP(16'hE952,4);
TASK_PP(16'hE953,4);
TASK_PP(16'hE954,4);
TASK_PP(16'hE955,4);
TASK_PP(16'hE956,4);
TASK_PP(16'hE957,4);
TASK_PP(16'hE958,4);
TASK_PP(16'hE959,4);
TASK_PP(16'hE95A,4);
TASK_PP(16'hE95B,4);
TASK_PP(16'hE95C,4);
TASK_PP(16'hE95D,4);
TASK_PP(16'hE95E,4);
TASK_PP(16'hE95F,4);
TASK_PP(16'hE960,4);
TASK_PP(16'hE961,4);
TASK_PP(16'hE962,4);
TASK_PP(16'hE963,4);
TASK_PP(16'hE964,4);
TASK_PP(16'hE965,4);
TASK_PP(16'hE966,4);
TASK_PP(16'hE967,4);
TASK_PP(16'hE968,4);
TASK_PP(16'hE969,4);
TASK_PP(16'hE96A,4);
TASK_PP(16'hE96B,4);
TASK_PP(16'hE96C,4);
TASK_PP(16'hE96D,4);
TASK_PP(16'hE96E,4);
TASK_PP(16'hE96F,4);
TASK_PP(16'hE970,4);
TASK_PP(16'hE971,4);
TASK_PP(16'hE972,4);
TASK_PP(16'hE973,4);
TASK_PP(16'hE974,4);
TASK_PP(16'hE975,4);
TASK_PP(16'hE976,4);
TASK_PP(16'hE977,4);
TASK_PP(16'hE978,4);
TASK_PP(16'hE979,4);
TASK_PP(16'hE97A,4);
TASK_PP(16'hE97B,4);
TASK_PP(16'hE97C,4);
TASK_PP(16'hE97D,4);
TASK_PP(16'hE97E,4);
TASK_PP(16'hE97F,4);
TASK_PP(16'hE980,4);
TASK_PP(16'hE981,4);
TASK_PP(16'hE982,4);
TASK_PP(16'hE983,4);
TASK_PP(16'hE984,4);
TASK_PP(16'hE985,4);
TASK_PP(16'hE986,4);
TASK_PP(16'hE987,4);
TASK_PP(16'hE988,4);
TASK_PP(16'hE989,4);
TASK_PP(16'hE98A,4);
TASK_PP(16'hE98B,4);
TASK_PP(16'hE98C,4);
TASK_PP(16'hE98D,4);
TASK_PP(16'hE98E,4);
TASK_PP(16'hE98F,4);
TASK_PP(16'hE990,4);
TASK_PP(16'hE991,4);
TASK_PP(16'hE992,4);
TASK_PP(16'hE993,4);
TASK_PP(16'hE994,4);
TASK_PP(16'hE995,4);
TASK_PP(16'hE996,4);
TASK_PP(16'hE997,4);
TASK_PP(16'hE998,4);
TASK_PP(16'hE999,4);
TASK_PP(16'hE99A,4);
TASK_PP(16'hE99B,4);
TASK_PP(16'hE99C,4);
TASK_PP(16'hE99D,4);
TASK_PP(16'hE99E,4);
TASK_PP(16'hE99F,4);
TASK_PP(16'hE9A0,4);
TASK_PP(16'hE9A1,4);
TASK_PP(16'hE9A2,4);
TASK_PP(16'hE9A3,4);
TASK_PP(16'hE9A4,4);
TASK_PP(16'hE9A5,4);
TASK_PP(16'hE9A6,4);
TASK_PP(16'hE9A7,4);
TASK_PP(16'hE9A8,4);
TASK_PP(16'hE9A9,4);
TASK_PP(16'hE9AA,4);
TASK_PP(16'hE9AB,4);
TASK_PP(16'hE9AC,4);
TASK_PP(16'hE9AD,4);
TASK_PP(16'hE9AE,4);
TASK_PP(16'hE9AF,4);
TASK_PP(16'hE9B0,4);
TASK_PP(16'hE9B1,4);
TASK_PP(16'hE9B2,4);
TASK_PP(16'hE9B3,4);
TASK_PP(16'hE9B4,4);
TASK_PP(16'hE9B5,4);
TASK_PP(16'hE9B6,4);
TASK_PP(16'hE9B7,4);
TASK_PP(16'hE9B8,4);
TASK_PP(16'hE9B9,4);
TASK_PP(16'hE9BA,4);
TASK_PP(16'hE9BB,4);
TASK_PP(16'hE9BC,4);
TASK_PP(16'hE9BD,4);
TASK_PP(16'hE9BE,4);
TASK_PP(16'hE9BF,4);
TASK_PP(16'hE9C0,4);
TASK_PP(16'hE9C1,4);
TASK_PP(16'hE9C2,4);
TASK_PP(16'hE9C3,4);
TASK_PP(16'hE9C4,4);
TASK_PP(16'hE9C5,4);
TASK_PP(16'hE9C6,4);
TASK_PP(16'hE9C7,4);
TASK_PP(16'hE9C8,4);
TASK_PP(16'hE9C9,4);
TASK_PP(16'hE9CA,4);
TASK_PP(16'hE9CB,4);
TASK_PP(16'hE9CC,4);
TASK_PP(16'hE9CD,4);
TASK_PP(16'hE9CE,4);
TASK_PP(16'hE9CF,4);
TASK_PP(16'hE9D0,4);
TASK_PP(16'hE9D1,4);
TASK_PP(16'hE9D2,4);
TASK_PP(16'hE9D3,4);
TASK_PP(16'hE9D4,4);
TASK_PP(16'hE9D5,4);
TASK_PP(16'hE9D6,4);
TASK_PP(16'hE9D7,4);
TASK_PP(16'hE9D8,4);
TASK_PP(16'hE9D9,4);
TASK_PP(16'hE9DA,4);
TASK_PP(16'hE9DB,4);
TASK_PP(16'hE9DC,4);
TASK_PP(16'hE9DD,4);
TASK_PP(16'hE9DE,4);
TASK_PP(16'hE9DF,4);
TASK_PP(16'hE9E0,4);
TASK_PP(16'hE9E1,4);
TASK_PP(16'hE9E2,4);
TASK_PP(16'hE9E3,4);
TASK_PP(16'hE9E4,4);
TASK_PP(16'hE9E5,4);
TASK_PP(16'hE9E6,4);
TASK_PP(16'hE9E7,4);
TASK_PP(16'hE9E8,4);
TASK_PP(16'hE9E9,4);
TASK_PP(16'hE9EA,4);
TASK_PP(16'hE9EB,4);
TASK_PP(16'hE9EC,4);
TASK_PP(16'hE9ED,4);
TASK_PP(16'hE9EE,4);
TASK_PP(16'hE9EF,4);
TASK_PP(16'hE9F0,4);
TASK_PP(16'hE9F1,4);
TASK_PP(16'hE9F2,4);
TASK_PP(16'hE9F3,4);
TASK_PP(16'hE9F4,4);
TASK_PP(16'hE9F5,4);
TASK_PP(16'hE9F6,4);
TASK_PP(16'hE9F7,4);
TASK_PP(16'hE9F8,4);
TASK_PP(16'hE9F9,4);
TASK_PP(16'hE9FA,4);
TASK_PP(16'hE9FB,4);
TASK_PP(16'hE9FC,4);
TASK_PP(16'hE9FD,4);
TASK_PP(16'hE9FE,4);
TASK_PP(16'hE9FF,4);
TASK_PP(16'hEA00,4);
TASK_PP(16'hEA01,4);
TASK_PP(16'hEA02,4);
TASK_PP(16'hEA03,4);
TASK_PP(16'hEA04,4);
TASK_PP(16'hEA05,4);
TASK_PP(16'hEA06,4);
TASK_PP(16'hEA07,4);
TASK_PP(16'hEA08,4);
TASK_PP(16'hEA09,4);
TASK_PP(16'hEA0A,4);
TASK_PP(16'hEA0B,4);
TASK_PP(16'hEA0C,4);
TASK_PP(16'hEA0D,4);
TASK_PP(16'hEA0E,4);
TASK_PP(16'hEA0F,4);
TASK_PP(16'hEA10,4);
TASK_PP(16'hEA11,4);
TASK_PP(16'hEA12,4);
TASK_PP(16'hEA13,4);
TASK_PP(16'hEA14,4);
TASK_PP(16'hEA15,4);
TASK_PP(16'hEA16,4);
TASK_PP(16'hEA17,4);
TASK_PP(16'hEA18,4);
TASK_PP(16'hEA19,4);
TASK_PP(16'hEA1A,4);
TASK_PP(16'hEA1B,4);
TASK_PP(16'hEA1C,4);
TASK_PP(16'hEA1D,4);
TASK_PP(16'hEA1E,4);
TASK_PP(16'hEA1F,4);
TASK_PP(16'hEA20,4);
TASK_PP(16'hEA21,4);
TASK_PP(16'hEA22,4);
TASK_PP(16'hEA23,4);
TASK_PP(16'hEA24,4);
TASK_PP(16'hEA25,4);
TASK_PP(16'hEA26,4);
TASK_PP(16'hEA27,4);
TASK_PP(16'hEA28,4);
TASK_PP(16'hEA29,4);
TASK_PP(16'hEA2A,4);
TASK_PP(16'hEA2B,4);
TASK_PP(16'hEA2C,4);
TASK_PP(16'hEA2D,4);
TASK_PP(16'hEA2E,4);
TASK_PP(16'hEA2F,4);
TASK_PP(16'hEA30,4);
TASK_PP(16'hEA31,4);
TASK_PP(16'hEA32,4);
TASK_PP(16'hEA33,4);
TASK_PP(16'hEA34,4);
TASK_PP(16'hEA35,4);
TASK_PP(16'hEA36,4);
TASK_PP(16'hEA37,4);
TASK_PP(16'hEA38,4);
TASK_PP(16'hEA39,4);
TASK_PP(16'hEA3A,4);
TASK_PP(16'hEA3B,4);
TASK_PP(16'hEA3C,4);
TASK_PP(16'hEA3D,4);
TASK_PP(16'hEA3E,4);
TASK_PP(16'hEA3F,4);
TASK_PP(16'hEA40,4);
TASK_PP(16'hEA41,4);
TASK_PP(16'hEA42,4);
TASK_PP(16'hEA43,4);
TASK_PP(16'hEA44,4);
TASK_PP(16'hEA45,4);
TASK_PP(16'hEA46,4);
TASK_PP(16'hEA47,4);
TASK_PP(16'hEA48,4);
TASK_PP(16'hEA49,4);
TASK_PP(16'hEA4A,4);
TASK_PP(16'hEA4B,4);
TASK_PP(16'hEA4C,4);
TASK_PP(16'hEA4D,4);
TASK_PP(16'hEA4E,4);
TASK_PP(16'hEA4F,4);
TASK_PP(16'hEA50,4);
TASK_PP(16'hEA51,4);
TASK_PP(16'hEA52,4);
TASK_PP(16'hEA53,4);
TASK_PP(16'hEA54,4);
TASK_PP(16'hEA55,4);
TASK_PP(16'hEA56,4);
TASK_PP(16'hEA57,4);
TASK_PP(16'hEA58,4);
TASK_PP(16'hEA59,4);
TASK_PP(16'hEA5A,4);
TASK_PP(16'hEA5B,4);
TASK_PP(16'hEA5C,4);
TASK_PP(16'hEA5D,4);
TASK_PP(16'hEA5E,4);
TASK_PP(16'hEA5F,4);
TASK_PP(16'hEA60,4);
TASK_PP(16'hEA61,4);
TASK_PP(16'hEA62,4);
TASK_PP(16'hEA63,4);
TASK_PP(16'hEA64,4);
TASK_PP(16'hEA65,4);
TASK_PP(16'hEA66,4);
TASK_PP(16'hEA67,4);
TASK_PP(16'hEA68,4);
TASK_PP(16'hEA69,4);
TASK_PP(16'hEA6A,4);
TASK_PP(16'hEA6B,4);
TASK_PP(16'hEA6C,4);
TASK_PP(16'hEA6D,4);
TASK_PP(16'hEA6E,4);
TASK_PP(16'hEA6F,4);
TASK_PP(16'hEA70,4);
TASK_PP(16'hEA71,4);
TASK_PP(16'hEA72,4);
TASK_PP(16'hEA73,4);
TASK_PP(16'hEA74,4);
TASK_PP(16'hEA75,4);
TASK_PP(16'hEA76,4);
TASK_PP(16'hEA77,4);
TASK_PP(16'hEA78,4);
TASK_PP(16'hEA79,4);
TASK_PP(16'hEA7A,4);
TASK_PP(16'hEA7B,4);
TASK_PP(16'hEA7C,4);
TASK_PP(16'hEA7D,4);
TASK_PP(16'hEA7E,4);
TASK_PP(16'hEA7F,4);
TASK_PP(16'hEA80,4);
TASK_PP(16'hEA81,4);
TASK_PP(16'hEA82,4);
TASK_PP(16'hEA83,4);
TASK_PP(16'hEA84,4);
TASK_PP(16'hEA85,4);
TASK_PP(16'hEA86,4);
TASK_PP(16'hEA87,4);
TASK_PP(16'hEA88,4);
TASK_PP(16'hEA89,4);
TASK_PP(16'hEA8A,4);
TASK_PP(16'hEA8B,4);
TASK_PP(16'hEA8C,4);
TASK_PP(16'hEA8D,4);
TASK_PP(16'hEA8E,4);
TASK_PP(16'hEA8F,4);
TASK_PP(16'hEA90,4);
TASK_PP(16'hEA91,4);
TASK_PP(16'hEA92,4);
TASK_PP(16'hEA93,4);
TASK_PP(16'hEA94,4);
TASK_PP(16'hEA95,4);
TASK_PP(16'hEA96,4);
TASK_PP(16'hEA97,4);
TASK_PP(16'hEA98,4);
TASK_PP(16'hEA99,4);
TASK_PP(16'hEA9A,4);
TASK_PP(16'hEA9B,4);
TASK_PP(16'hEA9C,4);
TASK_PP(16'hEA9D,4);
TASK_PP(16'hEA9E,4);
TASK_PP(16'hEA9F,4);
TASK_PP(16'hEAA0,4);
TASK_PP(16'hEAA1,4);
TASK_PP(16'hEAA2,4);
TASK_PP(16'hEAA3,4);
TASK_PP(16'hEAA4,4);
TASK_PP(16'hEAA5,4);
TASK_PP(16'hEAA6,4);
TASK_PP(16'hEAA7,4);
TASK_PP(16'hEAA8,4);
TASK_PP(16'hEAA9,4);
TASK_PP(16'hEAAA,4);
TASK_PP(16'hEAAB,4);
TASK_PP(16'hEAAC,4);
TASK_PP(16'hEAAD,4);
TASK_PP(16'hEAAE,4);
TASK_PP(16'hEAAF,4);
TASK_PP(16'hEAB0,4);
TASK_PP(16'hEAB1,4);
TASK_PP(16'hEAB2,4);
TASK_PP(16'hEAB3,4);
TASK_PP(16'hEAB4,4);
TASK_PP(16'hEAB5,4);
TASK_PP(16'hEAB6,4);
TASK_PP(16'hEAB7,4);
TASK_PP(16'hEAB8,4);
TASK_PP(16'hEAB9,4);
TASK_PP(16'hEABA,4);
TASK_PP(16'hEABB,4);
TASK_PP(16'hEABC,4);
TASK_PP(16'hEABD,4);
TASK_PP(16'hEABE,4);
TASK_PP(16'hEABF,4);
TASK_PP(16'hEAC0,4);
TASK_PP(16'hEAC1,4);
TASK_PP(16'hEAC2,4);
TASK_PP(16'hEAC3,4);
TASK_PP(16'hEAC4,4);
TASK_PP(16'hEAC5,4);
TASK_PP(16'hEAC6,4);
TASK_PP(16'hEAC7,4);
TASK_PP(16'hEAC8,4);
TASK_PP(16'hEAC9,4);
TASK_PP(16'hEACA,4);
TASK_PP(16'hEACB,4);
TASK_PP(16'hEACC,4);
TASK_PP(16'hEACD,4);
TASK_PP(16'hEACE,4);
TASK_PP(16'hEACF,4);
TASK_PP(16'hEAD0,4);
TASK_PP(16'hEAD1,4);
TASK_PP(16'hEAD2,4);
TASK_PP(16'hEAD3,4);
TASK_PP(16'hEAD4,4);
TASK_PP(16'hEAD5,4);
TASK_PP(16'hEAD6,4);
TASK_PP(16'hEAD7,4);
TASK_PP(16'hEAD8,4);
TASK_PP(16'hEAD9,4);
TASK_PP(16'hEADA,4);
TASK_PP(16'hEADB,4);
TASK_PP(16'hEADC,4);
TASK_PP(16'hEADD,4);
TASK_PP(16'hEADE,4);
TASK_PP(16'hEADF,4);
TASK_PP(16'hEAE0,4);
TASK_PP(16'hEAE1,4);
TASK_PP(16'hEAE2,4);
TASK_PP(16'hEAE3,4);
TASK_PP(16'hEAE4,4);
TASK_PP(16'hEAE5,4);
TASK_PP(16'hEAE6,4);
TASK_PP(16'hEAE7,4);
TASK_PP(16'hEAE8,4);
TASK_PP(16'hEAE9,4);
TASK_PP(16'hEAEA,4);
TASK_PP(16'hEAEB,4);
TASK_PP(16'hEAEC,4);
TASK_PP(16'hEAED,4);
TASK_PP(16'hEAEE,4);
TASK_PP(16'hEAEF,4);
TASK_PP(16'hEAF0,4);
TASK_PP(16'hEAF1,4);
TASK_PP(16'hEAF2,4);
TASK_PP(16'hEAF3,4);
TASK_PP(16'hEAF4,4);
TASK_PP(16'hEAF5,4);
TASK_PP(16'hEAF6,4);
TASK_PP(16'hEAF7,4);
TASK_PP(16'hEAF8,4);
TASK_PP(16'hEAF9,4);
TASK_PP(16'hEAFA,4);
TASK_PP(16'hEAFB,4);
TASK_PP(16'hEAFC,4);
TASK_PP(16'hEAFD,4);
TASK_PP(16'hEAFE,4);
TASK_PP(16'hEAFF,4);
TASK_PP(16'hEB00,4);
TASK_PP(16'hEB01,4);
TASK_PP(16'hEB02,4);
TASK_PP(16'hEB03,4);
TASK_PP(16'hEB04,4);
TASK_PP(16'hEB05,4);
TASK_PP(16'hEB06,4);
TASK_PP(16'hEB07,4);
TASK_PP(16'hEB08,4);
TASK_PP(16'hEB09,4);
TASK_PP(16'hEB0A,4);
TASK_PP(16'hEB0B,4);
TASK_PP(16'hEB0C,4);
TASK_PP(16'hEB0D,4);
TASK_PP(16'hEB0E,4);
TASK_PP(16'hEB0F,4);
TASK_PP(16'hEB10,4);
TASK_PP(16'hEB11,4);
TASK_PP(16'hEB12,4);
TASK_PP(16'hEB13,4);
TASK_PP(16'hEB14,4);
TASK_PP(16'hEB15,4);
TASK_PP(16'hEB16,4);
TASK_PP(16'hEB17,4);
TASK_PP(16'hEB18,4);
TASK_PP(16'hEB19,4);
TASK_PP(16'hEB1A,4);
TASK_PP(16'hEB1B,4);
TASK_PP(16'hEB1C,4);
TASK_PP(16'hEB1D,4);
TASK_PP(16'hEB1E,4);
TASK_PP(16'hEB1F,4);
TASK_PP(16'hEB20,4);
TASK_PP(16'hEB21,4);
TASK_PP(16'hEB22,4);
TASK_PP(16'hEB23,4);
TASK_PP(16'hEB24,4);
TASK_PP(16'hEB25,4);
TASK_PP(16'hEB26,4);
TASK_PP(16'hEB27,4);
TASK_PP(16'hEB28,4);
TASK_PP(16'hEB29,4);
TASK_PP(16'hEB2A,4);
TASK_PP(16'hEB2B,4);
TASK_PP(16'hEB2C,4);
TASK_PP(16'hEB2D,4);
TASK_PP(16'hEB2E,4);
TASK_PP(16'hEB2F,4);
TASK_PP(16'hEB30,4);
TASK_PP(16'hEB31,4);
TASK_PP(16'hEB32,4);
TASK_PP(16'hEB33,4);
TASK_PP(16'hEB34,4);
TASK_PP(16'hEB35,4);
TASK_PP(16'hEB36,4);
TASK_PP(16'hEB37,4);
TASK_PP(16'hEB38,4);
TASK_PP(16'hEB39,4);
TASK_PP(16'hEB3A,4);
TASK_PP(16'hEB3B,4);
TASK_PP(16'hEB3C,4);
TASK_PP(16'hEB3D,4);
TASK_PP(16'hEB3E,4);
TASK_PP(16'hEB3F,4);
TASK_PP(16'hEB40,4);
TASK_PP(16'hEB41,4);
TASK_PP(16'hEB42,4);
TASK_PP(16'hEB43,4);
TASK_PP(16'hEB44,4);
TASK_PP(16'hEB45,4);
TASK_PP(16'hEB46,4);
TASK_PP(16'hEB47,4);
TASK_PP(16'hEB48,4);
TASK_PP(16'hEB49,4);
TASK_PP(16'hEB4A,4);
TASK_PP(16'hEB4B,4);
TASK_PP(16'hEB4C,4);
TASK_PP(16'hEB4D,4);
TASK_PP(16'hEB4E,4);
TASK_PP(16'hEB4F,4);
TASK_PP(16'hEB50,4);
TASK_PP(16'hEB51,4);
TASK_PP(16'hEB52,4);
TASK_PP(16'hEB53,4);
TASK_PP(16'hEB54,4);
TASK_PP(16'hEB55,4);
TASK_PP(16'hEB56,4);
TASK_PP(16'hEB57,4);
TASK_PP(16'hEB58,4);
TASK_PP(16'hEB59,4);
TASK_PP(16'hEB5A,4);
TASK_PP(16'hEB5B,4);
TASK_PP(16'hEB5C,4);
TASK_PP(16'hEB5D,4);
TASK_PP(16'hEB5E,4);
TASK_PP(16'hEB5F,4);
TASK_PP(16'hEB60,4);
TASK_PP(16'hEB61,4);
TASK_PP(16'hEB62,4);
TASK_PP(16'hEB63,4);
TASK_PP(16'hEB64,4);
TASK_PP(16'hEB65,4);
TASK_PP(16'hEB66,4);
TASK_PP(16'hEB67,4);
TASK_PP(16'hEB68,4);
TASK_PP(16'hEB69,4);
TASK_PP(16'hEB6A,4);
TASK_PP(16'hEB6B,4);
TASK_PP(16'hEB6C,4);
TASK_PP(16'hEB6D,4);
TASK_PP(16'hEB6E,4);
TASK_PP(16'hEB6F,4);
TASK_PP(16'hEB70,4);
TASK_PP(16'hEB71,4);
TASK_PP(16'hEB72,4);
TASK_PP(16'hEB73,4);
TASK_PP(16'hEB74,4);
TASK_PP(16'hEB75,4);
TASK_PP(16'hEB76,4);
TASK_PP(16'hEB77,4);
TASK_PP(16'hEB78,4);
TASK_PP(16'hEB79,4);
TASK_PP(16'hEB7A,4);
TASK_PP(16'hEB7B,4);
TASK_PP(16'hEB7C,4);
TASK_PP(16'hEB7D,4);
TASK_PP(16'hEB7E,4);
TASK_PP(16'hEB7F,4);
TASK_PP(16'hEB80,4);
TASK_PP(16'hEB81,4);
TASK_PP(16'hEB82,4);
TASK_PP(16'hEB83,4);
TASK_PP(16'hEB84,4);
TASK_PP(16'hEB85,4);
TASK_PP(16'hEB86,4);
TASK_PP(16'hEB87,4);
TASK_PP(16'hEB88,4);
TASK_PP(16'hEB89,4);
TASK_PP(16'hEB8A,4);
TASK_PP(16'hEB8B,4);
TASK_PP(16'hEB8C,4);
TASK_PP(16'hEB8D,4);
TASK_PP(16'hEB8E,4);
TASK_PP(16'hEB8F,4);
TASK_PP(16'hEB90,4);
TASK_PP(16'hEB91,4);
TASK_PP(16'hEB92,4);
TASK_PP(16'hEB93,4);
TASK_PP(16'hEB94,4);
TASK_PP(16'hEB95,4);
TASK_PP(16'hEB96,4);
TASK_PP(16'hEB97,4);
TASK_PP(16'hEB98,4);
TASK_PP(16'hEB99,4);
TASK_PP(16'hEB9A,4);
TASK_PP(16'hEB9B,4);
TASK_PP(16'hEB9C,4);
TASK_PP(16'hEB9D,4);
TASK_PP(16'hEB9E,4);
TASK_PP(16'hEB9F,4);
TASK_PP(16'hEBA0,4);
TASK_PP(16'hEBA1,4);
TASK_PP(16'hEBA2,4);
TASK_PP(16'hEBA3,4);
TASK_PP(16'hEBA4,4);
TASK_PP(16'hEBA5,4);
TASK_PP(16'hEBA6,4);
TASK_PP(16'hEBA7,4);
TASK_PP(16'hEBA8,4);
TASK_PP(16'hEBA9,4);
TASK_PP(16'hEBAA,4);
TASK_PP(16'hEBAB,4);
TASK_PP(16'hEBAC,4);
TASK_PP(16'hEBAD,4);
TASK_PP(16'hEBAE,4);
TASK_PP(16'hEBAF,4);
TASK_PP(16'hEBB0,4);
TASK_PP(16'hEBB1,4);
TASK_PP(16'hEBB2,4);
TASK_PP(16'hEBB3,4);
TASK_PP(16'hEBB4,4);
TASK_PP(16'hEBB5,4);
TASK_PP(16'hEBB6,4);
TASK_PP(16'hEBB7,4);
TASK_PP(16'hEBB8,4);
TASK_PP(16'hEBB9,4);
TASK_PP(16'hEBBA,4);
TASK_PP(16'hEBBB,4);
TASK_PP(16'hEBBC,4);
TASK_PP(16'hEBBD,4);
TASK_PP(16'hEBBE,4);
TASK_PP(16'hEBBF,4);
TASK_PP(16'hEBC0,4);
TASK_PP(16'hEBC1,4);
TASK_PP(16'hEBC2,4);
TASK_PP(16'hEBC3,4);
TASK_PP(16'hEBC4,4);
TASK_PP(16'hEBC5,4);
TASK_PP(16'hEBC6,4);
TASK_PP(16'hEBC7,4);
TASK_PP(16'hEBC8,4);
TASK_PP(16'hEBC9,4);
TASK_PP(16'hEBCA,4);
TASK_PP(16'hEBCB,4);
TASK_PP(16'hEBCC,4);
TASK_PP(16'hEBCD,4);
TASK_PP(16'hEBCE,4);
TASK_PP(16'hEBCF,4);
TASK_PP(16'hEBD0,4);
TASK_PP(16'hEBD1,4);
TASK_PP(16'hEBD2,4);
TASK_PP(16'hEBD3,4);
TASK_PP(16'hEBD4,4);
TASK_PP(16'hEBD5,4);
TASK_PP(16'hEBD6,4);
TASK_PP(16'hEBD7,4);
TASK_PP(16'hEBD8,4);
TASK_PP(16'hEBD9,4);
TASK_PP(16'hEBDA,4);
TASK_PP(16'hEBDB,4);
TASK_PP(16'hEBDC,4);
TASK_PP(16'hEBDD,4);
TASK_PP(16'hEBDE,4);
TASK_PP(16'hEBDF,4);
TASK_PP(16'hEBE0,4);
TASK_PP(16'hEBE1,4);
TASK_PP(16'hEBE2,4);
TASK_PP(16'hEBE3,4);
TASK_PP(16'hEBE4,4);
TASK_PP(16'hEBE5,4);
TASK_PP(16'hEBE6,4);
TASK_PP(16'hEBE7,4);
TASK_PP(16'hEBE8,4);
TASK_PP(16'hEBE9,4);
TASK_PP(16'hEBEA,4);
TASK_PP(16'hEBEB,4);
TASK_PP(16'hEBEC,4);
TASK_PP(16'hEBED,4);
TASK_PP(16'hEBEE,4);
TASK_PP(16'hEBEF,4);
TASK_PP(16'hEBF0,4);
TASK_PP(16'hEBF1,4);
TASK_PP(16'hEBF2,4);
TASK_PP(16'hEBF3,4);
TASK_PP(16'hEBF4,4);
TASK_PP(16'hEBF5,4);
TASK_PP(16'hEBF6,4);
TASK_PP(16'hEBF7,4);
TASK_PP(16'hEBF8,4);
TASK_PP(16'hEBF9,4);
TASK_PP(16'hEBFA,4);
TASK_PP(16'hEBFB,4);
TASK_PP(16'hEBFC,4);
TASK_PP(16'hEBFD,4);
TASK_PP(16'hEBFE,4);
TASK_PP(16'hEBFF,4);
TASK_PP(16'hEC00,4);
TASK_PP(16'hEC01,4);
TASK_PP(16'hEC02,4);
TASK_PP(16'hEC03,4);
TASK_PP(16'hEC04,4);
TASK_PP(16'hEC05,4);
TASK_PP(16'hEC06,4);
TASK_PP(16'hEC07,4);
TASK_PP(16'hEC08,4);
TASK_PP(16'hEC09,4);
TASK_PP(16'hEC0A,4);
TASK_PP(16'hEC0B,4);
TASK_PP(16'hEC0C,4);
TASK_PP(16'hEC0D,4);
TASK_PP(16'hEC0E,4);
TASK_PP(16'hEC0F,4);
TASK_PP(16'hEC10,4);
TASK_PP(16'hEC11,4);
TASK_PP(16'hEC12,4);
TASK_PP(16'hEC13,4);
TASK_PP(16'hEC14,4);
TASK_PP(16'hEC15,4);
TASK_PP(16'hEC16,4);
TASK_PP(16'hEC17,4);
TASK_PP(16'hEC18,4);
TASK_PP(16'hEC19,4);
TASK_PP(16'hEC1A,4);
TASK_PP(16'hEC1B,4);
TASK_PP(16'hEC1C,4);
TASK_PP(16'hEC1D,4);
TASK_PP(16'hEC1E,4);
TASK_PP(16'hEC1F,4);
TASK_PP(16'hEC20,4);
TASK_PP(16'hEC21,4);
TASK_PP(16'hEC22,4);
TASK_PP(16'hEC23,4);
TASK_PP(16'hEC24,4);
TASK_PP(16'hEC25,4);
TASK_PP(16'hEC26,4);
TASK_PP(16'hEC27,4);
TASK_PP(16'hEC28,4);
TASK_PP(16'hEC29,4);
TASK_PP(16'hEC2A,4);
TASK_PP(16'hEC2B,4);
TASK_PP(16'hEC2C,4);
TASK_PP(16'hEC2D,4);
TASK_PP(16'hEC2E,4);
TASK_PP(16'hEC2F,4);
TASK_PP(16'hEC30,4);
TASK_PP(16'hEC31,4);
TASK_PP(16'hEC32,4);
TASK_PP(16'hEC33,4);
TASK_PP(16'hEC34,4);
TASK_PP(16'hEC35,4);
TASK_PP(16'hEC36,4);
TASK_PP(16'hEC37,4);
TASK_PP(16'hEC38,4);
TASK_PP(16'hEC39,4);
TASK_PP(16'hEC3A,4);
TASK_PP(16'hEC3B,4);
TASK_PP(16'hEC3C,4);
TASK_PP(16'hEC3D,4);
TASK_PP(16'hEC3E,4);
TASK_PP(16'hEC3F,4);
TASK_PP(16'hEC40,4);
TASK_PP(16'hEC41,4);
TASK_PP(16'hEC42,4);
TASK_PP(16'hEC43,4);
TASK_PP(16'hEC44,4);
TASK_PP(16'hEC45,4);
TASK_PP(16'hEC46,4);
TASK_PP(16'hEC47,4);
TASK_PP(16'hEC48,4);
TASK_PP(16'hEC49,4);
TASK_PP(16'hEC4A,4);
TASK_PP(16'hEC4B,4);
TASK_PP(16'hEC4C,4);
TASK_PP(16'hEC4D,4);
TASK_PP(16'hEC4E,4);
TASK_PP(16'hEC4F,4);
TASK_PP(16'hEC50,4);
TASK_PP(16'hEC51,4);
TASK_PP(16'hEC52,4);
TASK_PP(16'hEC53,4);
TASK_PP(16'hEC54,4);
TASK_PP(16'hEC55,4);
TASK_PP(16'hEC56,4);
TASK_PP(16'hEC57,4);
TASK_PP(16'hEC58,4);
TASK_PP(16'hEC59,4);
TASK_PP(16'hEC5A,4);
TASK_PP(16'hEC5B,4);
TASK_PP(16'hEC5C,4);
TASK_PP(16'hEC5D,4);
TASK_PP(16'hEC5E,4);
TASK_PP(16'hEC5F,4);
TASK_PP(16'hEC60,4);
TASK_PP(16'hEC61,4);
TASK_PP(16'hEC62,4);
TASK_PP(16'hEC63,4);
TASK_PP(16'hEC64,4);
TASK_PP(16'hEC65,4);
TASK_PP(16'hEC66,4);
TASK_PP(16'hEC67,4);
TASK_PP(16'hEC68,4);
TASK_PP(16'hEC69,4);
TASK_PP(16'hEC6A,4);
TASK_PP(16'hEC6B,4);
TASK_PP(16'hEC6C,4);
TASK_PP(16'hEC6D,4);
TASK_PP(16'hEC6E,4);
TASK_PP(16'hEC6F,4);
TASK_PP(16'hEC70,4);
TASK_PP(16'hEC71,4);
TASK_PP(16'hEC72,4);
TASK_PP(16'hEC73,4);
TASK_PP(16'hEC74,4);
TASK_PP(16'hEC75,4);
TASK_PP(16'hEC76,4);
TASK_PP(16'hEC77,4);
TASK_PP(16'hEC78,4);
TASK_PP(16'hEC79,4);
TASK_PP(16'hEC7A,4);
TASK_PP(16'hEC7B,4);
TASK_PP(16'hEC7C,4);
TASK_PP(16'hEC7D,4);
TASK_PP(16'hEC7E,4);
TASK_PP(16'hEC7F,4);
TASK_PP(16'hEC80,4);
TASK_PP(16'hEC81,4);
TASK_PP(16'hEC82,4);
TASK_PP(16'hEC83,4);
TASK_PP(16'hEC84,4);
TASK_PP(16'hEC85,4);
TASK_PP(16'hEC86,4);
TASK_PP(16'hEC87,4);
TASK_PP(16'hEC88,4);
TASK_PP(16'hEC89,4);
TASK_PP(16'hEC8A,4);
TASK_PP(16'hEC8B,4);
TASK_PP(16'hEC8C,4);
TASK_PP(16'hEC8D,4);
TASK_PP(16'hEC8E,4);
TASK_PP(16'hEC8F,4);
TASK_PP(16'hEC90,4);
TASK_PP(16'hEC91,4);
TASK_PP(16'hEC92,4);
TASK_PP(16'hEC93,4);
TASK_PP(16'hEC94,4);
TASK_PP(16'hEC95,4);
TASK_PP(16'hEC96,4);
TASK_PP(16'hEC97,4);
TASK_PP(16'hEC98,4);
TASK_PP(16'hEC99,4);
TASK_PP(16'hEC9A,4);
TASK_PP(16'hEC9B,4);
TASK_PP(16'hEC9C,4);
TASK_PP(16'hEC9D,4);
TASK_PP(16'hEC9E,4);
TASK_PP(16'hEC9F,4);
TASK_PP(16'hECA0,4);
TASK_PP(16'hECA1,4);
TASK_PP(16'hECA2,4);
TASK_PP(16'hECA3,4);
TASK_PP(16'hECA4,4);
TASK_PP(16'hECA5,4);
TASK_PP(16'hECA6,4);
TASK_PP(16'hECA7,4);
TASK_PP(16'hECA8,4);
TASK_PP(16'hECA9,4);
TASK_PP(16'hECAA,4);
TASK_PP(16'hECAB,4);
TASK_PP(16'hECAC,4);
TASK_PP(16'hECAD,4);
TASK_PP(16'hECAE,4);
TASK_PP(16'hECAF,4);
TASK_PP(16'hECB0,4);
TASK_PP(16'hECB1,4);
TASK_PP(16'hECB2,4);
TASK_PP(16'hECB3,4);
TASK_PP(16'hECB4,4);
TASK_PP(16'hECB5,4);
TASK_PP(16'hECB6,4);
TASK_PP(16'hECB7,4);
TASK_PP(16'hECB8,4);
TASK_PP(16'hECB9,4);
TASK_PP(16'hECBA,4);
TASK_PP(16'hECBB,4);
TASK_PP(16'hECBC,4);
TASK_PP(16'hECBD,4);
TASK_PP(16'hECBE,4);
TASK_PP(16'hECBF,4);
TASK_PP(16'hECC0,4);
TASK_PP(16'hECC1,4);
TASK_PP(16'hECC2,4);
TASK_PP(16'hECC3,4);
TASK_PP(16'hECC4,4);
TASK_PP(16'hECC5,4);
TASK_PP(16'hECC6,4);
TASK_PP(16'hECC7,4);
TASK_PP(16'hECC8,4);
TASK_PP(16'hECC9,4);
TASK_PP(16'hECCA,4);
TASK_PP(16'hECCB,4);
TASK_PP(16'hECCC,4);
TASK_PP(16'hECCD,4);
TASK_PP(16'hECCE,4);
TASK_PP(16'hECCF,4);
TASK_PP(16'hECD0,4);
TASK_PP(16'hECD1,4);
TASK_PP(16'hECD2,4);
TASK_PP(16'hECD3,4);
TASK_PP(16'hECD4,4);
TASK_PP(16'hECD5,4);
TASK_PP(16'hECD6,4);
TASK_PP(16'hECD7,4);
TASK_PP(16'hECD8,4);
TASK_PP(16'hECD9,4);
TASK_PP(16'hECDA,4);
TASK_PP(16'hECDB,4);
TASK_PP(16'hECDC,4);
TASK_PP(16'hECDD,4);
TASK_PP(16'hECDE,4);
TASK_PP(16'hECDF,4);
TASK_PP(16'hECE0,4);
TASK_PP(16'hECE1,4);
TASK_PP(16'hECE2,4);
TASK_PP(16'hECE3,4);
TASK_PP(16'hECE4,4);
TASK_PP(16'hECE5,4);
TASK_PP(16'hECE6,4);
TASK_PP(16'hECE7,4);
TASK_PP(16'hECE8,4);
TASK_PP(16'hECE9,4);
TASK_PP(16'hECEA,4);
TASK_PP(16'hECEB,4);
TASK_PP(16'hECEC,4);
TASK_PP(16'hECED,4);
TASK_PP(16'hECEE,4);
TASK_PP(16'hECEF,4);
TASK_PP(16'hECF0,4);
TASK_PP(16'hECF1,4);
TASK_PP(16'hECF2,4);
TASK_PP(16'hECF3,4);
TASK_PP(16'hECF4,4);
TASK_PP(16'hECF5,4);
TASK_PP(16'hECF6,4);
TASK_PP(16'hECF7,4);
TASK_PP(16'hECF8,4);
TASK_PP(16'hECF9,4);
TASK_PP(16'hECFA,4);
TASK_PP(16'hECFB,4);
TASK_PP(16'hECFC,4);
TASK_PP(16'hECFD,4);
TASK_PP(16'hECFE,4);
TASK_PP(16'hECFF,4);
TASK_PP(16'hED00,4);
TASK_PP(16'hED01,4);
TASK_PP(16'hED02,4);
TASK_PP(16'hED03,4);
TASK_PP(16'hED04,4);
TASK_PP(16'hED05,4);
TASK_PP(16'hED06,4);
TASK_PP(16'hED07,4);
TASK_PP(16'hED08,4);
TASK_PP(16'hED09,4);
TASK_PP(16'hED0A,4);
TASK_PP(16'hED0B,4);
TASK_PP(16'hED0C,4);
TASK_PP(16'hED0D,4);
TASK_PP(16'hED0E,4);
TASK_PP(16'hED0F,4);
TASK_PP(16'hED10,4);
TASK_PP(16'hED11,4);
TASK_PP(16'hED12,4);
TASK_PP(16'hED13,4);
TASK_PP(16'hED14,4);
TASK_PP(16'hED15,4);
TASK_PP(16'hED16,4);
TASK_PP(16'hED17,4);
TASK_PP(16'hED18,4);
TASK_PP(16'hED19,4);
TASK_PP(16'hED1A,4);
TASK_PP(16'hED1B,4);
TASK_PP(16'hED1C,4);
TASK_PP(16'hED1D,4);
TASK_PP(16'hED1E,4);
TASK_PP(16'hED1F,4);
TASK_PP(16'hED20,4);
TASK_PP(16'hED21,4);
TASK_PP(16'hED22,4);
TASK_PP(16'hED23,4);
TASK_PP(16'hED24,4);
TASK_PP(16'hED25,4);
TASK_PP(16'hED26,4);
TASK_PP(16'hED27,4);
TASK_PP(16'hED28,4);
TASK_PP(16'hED29,4);
TASK_PP(16'hED2A,4);
TASK_PP(16'hED2B,4);
TASK_PP(16'hED2C,4);
TASK_PP(16'hED2D,4);
TASK_PP(16'hED2E,4);
TASK_PP(16'hED2F,4);
TASK_PP(16'hED30,4);
TASK_PP(16'hED31,4);
TASK_PP(16'hED32,4);
TASK_PP(16'hED33,4);
TASK_PP(16'hED34,4);
TASK_PP(16'hED35,4);
TASK_PP(16'hED36,4);
TASK_PP(16'hED37,4);
TASK_PP(16'hED38,4);
TASK_PP(16'hED39,4);
TASK_PP(16'hED3A,4);
TASK_PP(16'hED3B,4);
TASK_PP(16'hED3C,4);
TASK_PP(16'hED3D,4);
TASK_PP(16'hED3E,4);
TASK_PP(16'hED3F,4);
TASK_PP(16'hED40,4);
TASK_PP(16'hED41,4);
TASK_PP(16'hED42,4);
TASK_PP(16'hED43,4);
TASK_PP(16'hED44,4);
TASK_PP(16'hED45,4);
TASK_PP(16'hED46,4);
TASK_PP(16'hED47,4);
TASK_PP(16'hED48,4);
TASK_PP(16'hED49,4);
TASK_PP(16'hED4A,4);
TASK_PP(16'hED4B,4);
TASK_PP(16'hED4C,4);
TASK_PP(16'hED4D,4);
TASK_PP(16'hED4E,4);
TASK_PP(16'hED4F,4);
TASK_PP(16'hED50,4);
TASK_PP(16'hED51,4);
TASK_PP(16'hED52,4);
TASK_PP(16'hED53,4);
TASK_PP(16'hED54,4);
TASK_PP(16'hED55,4);
TASK_PP(16'hED56,4);
TASK_PP(16'hED57,4);
TASK_PP(16'hED58,4);
TASK_PP(16'hED59,4);
TASK_PP(16'hED5A,4);
TASK_PP(16'hED5B,4);
TASK_PP(16'hED5C,4);
TASK_PP(16'hED5D,4);
TASK_PP(16'hED5E,4);
TASK_PP(16'hED5F,4);
TASK_PP(16'hED60,4);
TASK_PP(16'hED61,4);
TASK_PP(16'hED62,4);
TASK_PP(16'hED63,4);
TASK_PP(16'hED64,4);
TASK_PP(16'hED65,4);
TASK_PP(16'hED66,4);
TASK_PP(16'hED67,4);
TASK_PP(16'hED68,4);
TASK_PP(16'hED69,4);
TASK_PP(16'hED6A,4);
TASK_PP(16'hED6B,4);
TASK_PP(16'hED6C,4);
TASK_PP(16'hED6D,4);
TASK_PP(16'hED6E,4);
TASK_PP(16'hED6F,4);
TASK_PP(16'hED70,4);
TASK_PP(16'hED71,4);
TASK_PP(16'hED72,4);
TASK_PP(16'hED73,4);
TASK_PP(16'hED74,4);
TASK_PP(16'hED75,4);
TASK_PP(16'hED76,4);
TASK_PP(16'hED77,4);
TASK_PP(16'hED78,4);
TASK_PP(16'hED79,4);
TASK_PP(16'hED7A,4);
TASK_PP(16'hED7B,4);
TASK_PP(16'hED7C,4);
TASK_PP(16'hED7D,4);
TASK_PP(16'hED7E,4);
TASK_PP(16'hED7F,4);
TASK_PP(16'hED80,4);
TASK_PP(16'hED81,4);
TASK_PP(16'hED82,4);
TASK_PP(16'hED83,4);
TASK_PP(16'hED84,4);
TASK_PP(16'hED85,4);
TASK_PP(16'hED86,4);
TASK_PP(16'hED87,4);
TASK_PP(16'hED88,4);
TASK_PP(16'hED89,4);
TASK_PP(16'hED8A,4);
TASK_PP(16'hED8B,4);
TASK_PP(16'hED8C,4);
TASK_PP(16'hED8D,4);
TASK_PP(16'hED8E,4);
TASK_PP(16'hED8F,4);
TASK_PP(16'hED90,4);
TASK_PP(16'hED91,4);
TASK_PP(16'hED92,4);
TASK_PP(16'hED93,4);
TASK_PP(16'hED94,4);
TASK_PP(16'hED95,4);
TASK_PP(16'hED96,4);
TASK_PP(16'hED97,4);
TASK_PP(16'hED98,4);
TASK_PP(16'hED99,4);
TASK_PP(16'hED9A,4);
TASK_PP(16'hED9B,4);
TASK_PP(16'hED9C,4);
TASK_PP(16'hED9D,4);
TASK_PP(16'hED9E,4);
TASK_PP(16'hED9F,4);
TASK_PP(16'hEDA0,4);
TASK_PP(16'hEDA1,4);
TASK_PP(16'hEDA2,4);
TASK_PP(16'hEDA3,4);
TASK_PP(16'hEDA4,4);
TASK_PP(16'hEDA5,4);
TASK_PP(16'hEDA6,4);
TASK_PP(16'hEDA7,4);
TASK_PP(16'hEDA8,4);
TASK_PP(16'hEDA9,4);
TASK_PP(16'hEDAA,4);
TASK_PP(16'hEDAB,4);
TASK_PP(16'hEDAC,4);
TASK_PP(16'hEDAD,4);
TASK_PP(16'hEDAE,4);
TASK_PP(16'hEDAF,4);
TASK_PP(16'hEDB0,4);
TASK_PP(16'hEDB1,4);
TASK_PP(16'hEDB2,4);
TASK_PP(16'hEDB3,4);
TASK_PP(16'hEDB4,4);
TASK_PP(16'hEDB5,4);
TASK_PP(16'hEDB6,4);
TASK_PP(16'hEDB7,4);
TASK_PP(16'hEDB8,4);
TASK_PP(16'hEDB9,4);
TASK_PP(16'hEDBA,4);
TASK_PP(16'hEDBB,4);
TASK_PP(16'hEDBC,4);
TASK_PP(16'hEDBD,4);
TASK_PP(16'hEDBE,4);
TASK_PP(16'hEDBF,4);
TASK_PP(16'hEDC0,4);
TASK_PP(16'hEDC1,4);
TASK_PP(16'hEDC2,4);
TASK_PP(16'hEDC3,4);
TASK_PP(16'hEDC4,4);
TASK_PP(16'hEDC5,4);
TASK_PP(16'hEDC6,4);
TASK_PP(16'hEDC7,4);
TASK_PP(16'hEDC8,4);
TASK_PP(16'hEDC9,4);
TASK_PP(16'hEDCA,4);
TASK_PP(16'hEDCB,4);
TASK_PP(16'hEDCC,4);
TASK_PP(16'hEDCD,4);
TASK_PP(16'hEDCE,4);
TASK_PP(16'hEDCF,4);
TASK_PP(16'hEDD0,4);
TASK_PP(16'hEDD1,4);
TASK_PP(16'hEDD2,4);
TASK_PP(16'hEDD3,4);
TASK_PP(16'hEDD4,4);
TASK_PP(16'hEDD5,4);
TASK_PP(16'hEDD6,4);
TASK_PP(16'hEDD7,4);
TASK_PP(16'hEDD8,4);
TASK_PP(16'hEDD9,4);
TASK_PP(16'hEDDA,4);
TASK_PP(16'hEDDB,4);
TASK_PP(16'hEDDC,4);
TASK_PP(16'hEDDD,4);
TASK_PP(16'hEDDE,4);
TASK_PP(16'hEDDF,4);
TASK_PP(16'hEDE0,4);
TASK_PP(16'hEDE1,4);
TASK_PP(16'hEDE2,4);
TASK_PP(16'hEDE3,4);
TASK_PP(16'hEDE4,4);
TASK_PP(16'hEDE5,4);
TASK_PP(16'hEDE6,4);
TASK_PP(16'hEDE7,4);
TASK_PP(16'hEDE8,4);
TASK_PP(16'hEDE9,4);
TASK_PP(16'hEDEA,4);
TASK_PP(16'hEDEB,4);
TASK_PP(16'hEDEC,4);
TASK_PP(16'hEDED,4);
TASK_PP(16'hEDEE,4);
TASK_PP(16'hEDEF,4);
TASK_PP(16'hEDF0,4);
TASK_PP(16'hEDF1,4);
TASK_PP(16'hEDF2,4);
TASK_PP(16'hEDF3,4);
TASK_PP(16'hEDF4,4);
TASK_PP(16'hEDF5,4);
TASK_PP(16'hEDF6,4);
TASK_PP(16'hEDF7,4);
TASK_PP(16'hEDF8,4);
TASK_PP(16'hEDF9,4);
TASK_PP(16'hEDFA,4);
TASK_PP(16'hEDFB,4);
TASK_PP(16'hEDFC,4);
TASK_PP(16'hEDFD,4);
TASK_PP(16'hEDFE,4);
TASK_PP(16'hEDFF,4);
TASK_PP(16'hEE00,4);
TASK_PP(16'hEE01,4);
TASK_PP(16'hEE02,4);
TASK_PP(16'hEE03,4);
TASK_PP(16'hEE04,4);
TASK_PP(16'hEE05,4);
TASK_PP(16'hEE06,4);
TASK_PP(16'hEE07,4);
TASK_PP(16'hEE08,4);
TASK_PP(16'hEE09,4);
TASK_PP(16'hEE0A,4);
TASK_PP(16'hEE0B,4);
TASK_PP(16'hEE0C,4);
TASK_PP(16'hEE0D,4);
TASK_PP(16'hEE0E,4);
TASK_PP(16'hEE0F,4);
TASK_PP(16'hEE10,4);
TASK_PP(16'hEE11,4);
TASK_PP(16'hEE12,4);
TASK_PP(16'hEE13,4);
TASK_PP(16'hEE14,4);
TASK_PP(16'hEE15,4);
TASK_PP(16'hEE16,4);
TASK_PP(16'hEE17,4);
TASK_PP(16'hEE18,4);
TASK_PP(16'hEE19,4);
TASK_PP(16'hEE1A,4);
TASK_PP(16'hEE1B,4);
TASK_PP(16'hEE1C,4);
TASK_PP(16'hEE1D,4);
TASK_PP(16'hEE1E,4);
TASK_PP(16'hEE1F,4);
TASK_PP(16'hEE20,4);
TASK_PP(16'hEE21,4);
TASK_PP(16'hEE22,4);
TASK_PP(16'hEE23,4);
TASK_PP(16'hEE24,4);
TASK_PP(16'hEE25,4);
TASK_PP(16'hEE26,4);
TASK_PP(16'hEE27,4);
TASK_PP(16'hEE28,4);
TASK_PP(16'hEE29,4);
TASK_PP(16'hEE2A,4);
TASK_PP(16'hEE2B,4);
TASK_PP(16'hEE2C,4);
TASK_PP(16'hEE2D,4);
TASK_PP(16'hEE2E,4);
TASK_PP(16'hEE2F,4);
TASK_PP(16'hEE30,4);
TASK_PP(16'hEE31,4);
TASK_PP(16'hEE32,4);
TASK_PP(16'hEE33,4);
TASK_PP(16'hEE34,4);
TASK_PP(16'hEE35,4);
TASK_PP(16'hEE36,4);
TASK_PP(16'hEE37,4);
TASK_PP(16'hEE38,4);
TASK_PP(16'hEE39,4);
TASK_PP(16'hEE3A,4);
TASK_PP(16'hEE3B,4);
TASK_PP(16'hEE3C,4);
TASK_PP(16'hEE3D,4);
TASK_PP(16'hEE3E,4);
TASK_PP(16'hEE3F,4);
TASK_PP(16'hEE40,4);
TASK_PP(16'hEE41,4);
TASK_PP(16'hEE42,4);
TASK_PP(16'hEE43,4);
TASK_PP(16'hEE44,4);
TASK_PP(16'hEE45,4);
TASK_PP(16'hEE46,4);
TASK_PP(16'hEE47,4);
TASK_PP(16'hEE48,4);
TASK_PP(16'hEE49,4);
TASK_PP(16'hEE4A,4);
TASK_PP(16'hEE4B,4);
TASK_PP(16'hEE4C,4);
TASK_PP(16'hEE4D,4);
TASK_PP(16'hEE4E,4);
TASK_PP(16'hEE4F,4);
TASK_PP(16'hEE50,4);
TASK_PP(16'hEE51,4);
TASK_PP(16'hEE52,4);
TASK_PP(16'hEE53,4);
TASK_PP(16'hEE54,4);
TASK_PP(16'hEE55,4);
TASK_PP(16'hEE56,4);
TASK_PP(16'hEE57,4);
TASK_PP(16'hEE58,4);
TASK_PP(16'hEE59,4);
TASK_PP(16'hEE5A,4);
TASK_PP(16'hEE5B,4);
TASK_PP(16'hEE5C,4);
TASK_PP(16'hEE5D,4);
TASK_PP(16'hEE5E,4);
TASK_PP(16'hEE5F,4);
TASK_PP(16'hEE60,4);
TASK_PP(16'hEE61,4);
TASK_PP(16'hEE62,4);
TASK_PP(16'hEE63,4);
TASK_PP(16'hEE64,4);
TASK_PP(16'hEE65,4);
TASK_PP(16'hEE66,4);
TASK_PP(16'hEE67,4);
TASK_PP(16'hEE68,4);
TASK_PP(16'hEE69,4);
TASK_PP(16'hEE6A,4);
TASK_PP(16'hEE6B,4);
TASK_PP(16'hEE6C,4);
TASK_PP(16'hEE6D,4);
TASK_PP(16'hEE6E,4);
TASK_PP(16'hEE6F,4);
TASK_PP(16'hEE70,4);
TASK_PP(16'hEE71,4);
TASK_PP(16'hEE72,4);
TASK_PP(16'hEE73,4);
TASK_PP(16'hEE74,4);
TASK_PP(16'hEE75,4);
TASK_PP(16'hEE76,4);
TASK_PP(16'hEE77,4);
TASK_PP(16'hEE78,4);
TASK_PP(16'hEE79,4);
TASK_PP(16'hEE7A,4);
TASK_PP(16'hEE7B,4);
TASK_PP(16'hEE7C,4);
TASK_PP(16'hEE7D,4);
TASK_PP(16'hEE7E,4);
TASK_PP(16'hEE7F,4);
TASK_PP(16'hEE80,4);
TASK_PP(16'hEE81,4);
TASK_PP(16'hEE82,4);
TASK_PP(16'hEE83,4);
TASK_PP(16'hEE84,4);
TASK_PP(16'hEE85,4);
TASK_PP(16'hEE86,4);
TASK_PP(16'hEE87,4);
TASK_PP(16'hEE88,4);
TASK_PP(16'hEE89,4);
TASK_PP(16'hEE8A,4);
TASK_PP(16'hEE8B,4);
TASK_PP(16'hEE8C,4);
TASK_PP(16'hEE8D,4);
TASK_PP(16'hEE8E,4);
TASK_PP(16'hEE8F,4);
TASK_PP(16'hEE90,4);
TASK_PP(16'hEE91,4);
TASK_PP(16'hEE92,4);
TASK_PP(16'hEE93,4);
TASK_PP(16'hEE94,4);
TASK_PP(16'hEE95,4);
TASK_PP(16'hEE96,4);
TASK_PP(16'hEE97,4);
TASK_PP(16'hEE98,4);
TASK_PP(16'hEE99,4);
TASK_PP(16'hEE9A,4);
TASK_PP(16'hEE9B,4);
TASK_PP(16'hEE9C,4);
TASK_PP(16'hEE9D,4);
TASK_PP(16'hEE9E,4);
TASK_PP(16'hEE9F,4);
TASK_PP(16'hEEA0,4);
TASK_PP(16'hEEA1,4);
TASK_PP(16'hEEA2,4);
TASK_PP(16'hEEA3,4);
TASK_PP(16'hEEA4,4);
TASK_PP(16'hEEA5,4);
TASK_PP(16'hEEA6,4);
TASK_PP(16'hEEA7,4);
TASK_PP(16'hEEA8,4);
TASK_PP(16'hEEA9,4);
TASK_PP(16'hEEAA,4);
TASK_PP(16'hEEAB,4);
TASK_PP(16'hEEAC,4);
TASK_PP(16'hEEAD,4);
TASK_PP(16'hEEAE,4);
TASK_PP(16'hEEAF,4);
TASK_PP(16'hEEB0,4);
TASK_PP(16'hEEB1,4);
TASK_PP(16'hEEB2,4);
TASK_PP(16'hEEB3,4);
TASK_PP(16'hEEB4,4);
TASK_PP(16'hEEB5,4);
TASK_PP(16'hEEB6,4);
TASK_PP(16'hEEB7,4);
TASK_PP(16'hEEB8,4);
TASK_PP(16'hEEB9,4);
TASK_PP(16'hEEBA,4);
TASK_PP(16'hEEBB,4);
TASK_PP(16'hEEBC,4);
TASK_PP(16'hEEBD,4);
TASK_PP(16'hEEBE,4);
TASK_PP(16'hEEBF,4);
TASK_PP(16'hEEC0,4);
TASK_PP(16'hEEC1,4);
TASK_PP(16'hEEC2,4);
TASK_PP(16'hEEC3,4);
TASK_PP(16'hEEC4,4);
TASK_PP(16'hEEC5,4);
TASK_PP(16'hEEC6,4);
TASK_PP(16'hEEC7,4);
TASK_PP(16'hEEC8,4);
TASK_PP(16'hEEC9,4);
TASK_PP(16'hEECA,4);
TASK_PP(16'hEECB,4);
TASK_PP(16'hEECC,4);
TASK_PP(16'hEECD,4);
TASK_PP(16'hEECE,4);
TASK_PP(16'hEECF,4);
TASK_PP(16'hEED0,4);
TASK_PP(16'hEED1,4);
TASK_PP(16'hEED2,4);
TASK_PP(16'hEED3,4);
TASK_PP(16'hEED4,4);
TASK_PP(16'hEED5,4);
TASK_PP(16'hEED6,4);
TASK_PP(16'hEED7,4);
TASK_PP(16'hEED8,4);
TASK_PP(16'hEED9,4);
TASK_PP(16'hEEDA,4);
TASK_PP(16'hEEDB,4);
TASK_PP(16'hEEDC,4);
TASK_PP(16'hEEDD,4);
TASK_PP(16'hEEDE,4);
TASK_PP(16'hEEDF,4);
TASK_PP(16'hEEE0,4);
TASK_PP(16'hEEE1,4);
TASK_PP(16'hEEE2,4);
TASK_PP(16'hEEE3,4);
TASK_PP(16'hEEE4,4);
TASK_PP(16'hEEE5,4);
TASK_PP(16'hEEE6,4);
TASK_PP(16'hEEE7,4);
TASK_PP(16'hEEE8,4);
TASK_PP(16'hEEE9,4);
TASK_PP(16'hEEEA,4);
TASK_PP(16'hEEEB,4);
TASK_PP(16'hEEEC,4);
TASK_PP(16'hEEED,4);
TASK_PP(16'hEEEE,4);
TASK_PP(16'hEEEF,4);
TASK_PP(16'hEEF0,4);
TASK_PP(16'hEEF1,4);
TASK_PP(16'hEEF2,4);
TASK_PP(16'hEEF3,4);
TASK_PP(16'hEEF4,4);
TASK_PP(16'hEEF5,4);
TASK_PP(16'hEEF6,4);
TASK_PP(16'hEEF7,4);
TASK_PP(16'hEEF8,4);
TASK_PP(16'hEEF9,4);
TASK_PP(16'hEEFA,4);
TASK_PP(16'hEEFB,4);
TASK_PP(16'hEEFC,4);
TASK_PP(16'hEEFD,4);
TASK_PP(16'hEEFE,4);
TASK_PP(16'hEEFF,4);
TASK_PP(16'hEF00,4);
TASK_PP(16'hEF01,4);
TASK_PP(16'hEF02,4);
TASK_PP(16'hEF03,4);
TASK_PP(16'hEF04,4);
TASK_PP(16'hEF05,4);
TASK_PP(16'hEF06,4);
TASK_PP(16'hEF07,4);
TASK_PP(16'hEF08,4);
TASK_PP(16'hEF09,4);
TASK_PP(16'hEF0A,4);
TASK_PP(16'hEF0B,4);
TASK_PP(16'hEF0C,4);
TASK_PP(16'hEF0D,4);
TASK_PP(16'hEF0E,4);
TASK_PP(16'hEF0F,4);
TASK_PP(16'hEF10,4);
TASK_PP(16'hEF11,4);
TASK_PP(16'hEF12,4);
TASK_PP(16'hEF13,4);
TASK_PP(16'hEF14,4);
TASK_PP(16'hEF15,4);
TASK_PP(16'hEF16,4);
TASK_PP(16'hEF17,4);
TASK_PP(16'hEF18,4);
TASK_PP(16'hEF19,4);
TASK_PP(16'hEF1A,4);
TASK_PP(16'hEF1B,4);
TASK_PP(16'hEF1C,4);
TASK_PP(16'hEF1D,4);
TASK_PP(16'hEF1E,4);
TASK_PP(16'hEF1F,4);
TASK_PP(16'hEF20,4);
TASK_PP(16'hEF21,4);
TASK_PP(16'hEF22,4);
TASK_PP(16'hEF23,4);
TASK_PP(16'hEF24,4);
TASK_PP(16'hEF25,4);
TASK_PP(16'hEF26,4);
TASK_PP(16'hEF27,4);
TASK_PP(16'hEF28,4);
TASK_PP(16'hEF29,4);
TASK_PP(16'hEF2A,4);
TASK_PP(16'hEF2B,4);
TASK_PP(16'hEF2C,4);
TASK_PP(16'hEF2D,4);
TASK_PP(16'hEF2E,4);
TASK_PP(16'hEF2F,4);
TASK_PP(16'hEF30,4);
TASK_PP(16'hEF31,4);
TASK_PP(16'hEF32,4);
TASK_PP(16'hEF33,4);
TASK_PP(16'hEF34,4);
TASK_PP(16'hEF35,4);
TASK_PP(16'hEF36,4);
TASK_PP(16'hEF37,4);
TASK_PP(16'hEF38,4);
TASK_PP(16'hEF39,4);
TASK_PP(16'hEF3A,4);
TASK_PP(16'hEF3B,4);
TASK_PP(16'hEF3C,4);
TASK_PP(16'hEF3D,4);
TASK_PP(16'hEF3E,4);
TASK_PP(16'hEF3F,4);
TASK_PP(16'hEF40,4);
TASK_PP(16'hEF41,4);
TASK_PP(16'hEF42,4);
TASK_PP(16'hEF43,4);
TASK_PP(16'hEF44,4);
TASK_PP(16'hEF45,4);
TASK_PP(16'hEF46,4);
TASK_PP(16'hEF47,4);
TASK_PP(16'hEF48,4);
TASK_PP(16'hEF49,4);
TASK_PP(16'hEF4A,4);
TASK_PP(16'hEF4B,4);
TASK_PP(16'hEF4C,4);
TASK_PP(16'hEF4D,4);
TASK_PP(16'hEF4E,4);
TASK_PP(16'hEF4F,4);
TASK_PP(16'hEF50,4);
TASK_PP(16'hEF51,4);
TASK_PP(16'hEF52,4);
TASK_PP(16'hEF53,4);
TASK_PP(16'hEF54,4);
TASK_PP(16'hEF55,4);
TASK_PP(16'hEF56,4);
TASK_PP(16'hEF57,4);
TASK_PP(16'hEF58,4);
TASK_PP(16'hEF59,4);
TASK_PP(16'hEF5A,4);
TASK_PP(16'hEF5B,4);
TASK_PP(16'hEF5C,4);
TASK_PP(16'hEF5D,4);
TASK_PP(16'hEF5E,4);
TASK_PP(16'hEF5F,4);
TASK_PP(16'hEF60,4);
TASK_PP(16'hEF61,4);
TASK_PP(16'hEF62,4);
TASK_PP(16'hEF63,4);
TASK_PP(16'hEF64,4);
TASK_PP(16'hEF65,4);
TASK_PP(16'hEF66,4);
TASK_PP(16'hEF67,4);
TASK_PP(16'hEF68,4);
TASK_PP(16'hEF69,4);
TASK_PP(16'hEF6A,4);
TASK_PP(16'hEF6B,4);
TASK_PP(16'hEF6C,4);
TASK_PP(16'hEF6D,4);
TASK_PP(16'hEF6E,4);
TASK_PP(16'hEF6F,4);
TASK_PP(16'hEF70,4);
TASK_PP(16'hEF71,4);
TASK_PP(16'hEF72,4);
TASK_PP(16'hEF73,4);
TASK_PP(16'hEF74,4);
TASK_PP(16'hEF75,4);
TASK_PP(16'hEF76,4);
TASK_PP(16'hEF77,4);
TASK_PP(16'hEF78,4);
TASK_PP(16'hEF79,4);
TASK_PP(16'hEF7A,4);
TASK_PP(16'hEF7B,4);
TASK_PP(16'hEF7C,4);
TASK_PP(16'hEF7D,4);
TASK_PP(16'hEF7E,4);
TASK_PP(16'hEF7F,4);
TASK_PP(16'hEF80,4);
TASK_PP(16'hEF81,4);
TASK_PP(16'hEF82,4);
TASK_PP(16'hEF83,4);
TASK_PP(16'hEF84,4);
TASK_PP(16'hEF85,4);
TASK_PP(16'hEF86,4);
TASK_PP(16'hEF87,4);
TASK_PP(16'hEF88,4);
TASK_PP(16'hEF89,4);
TASK_PP(16'hEF8A,4);
TASK_PP(16'hEF8B,4);
TASK_PP(16'hEF8C,4);
TASK_PP(16'hEF8D,4);
TASK_PP(16'hEF8E,4);
TASK_PP(16'hEF8F,4);
TASK_PP(16'hEF90,4);
TASK_PP(16'hEF91,4);
TASK_PP(16'hEF92,4);
TASK_PP(16'hEF93,4);
TASK_PP(16'hEF94,4);
TASK_PP(16'hEF95,4);
TASK_PP(16'hEF96,4);
TASK_PP(16'hEF97,4);
TASK_PP(16'hEF98,4);
TASK_PP(16'hEF99,4);
TASK_PP(16'hEF9A,4);
TASK_PP(16'hEF9B,4);
TASK_PP(16'hEF9C,4);
TASK_PP(16'hEF9D,4);
TASK_PP(16'hEF9E,4);
TASK_PP(16'hEF9F,4);
TASK_PP(16'hEFA0,4);
TASK_PP(16'hEFA1,4);
TASK_PP(16'hEFA2,4);
TASK_PP(16'hEFA3,4);
TASK_PP(16'hEFA4,4);
TASK_PP(16'hEFA5,4);
TASK_PP(16'hEFA6,4);
TASK_PP(16'hEFA7,4);
TASK_PP(16'hEFA8,4);
TASK_PP(16'hEFA9,4);
TASK_PP(16'hEFAA,4);
TASK_PP(16'hEFAB,4);
TASK_PP(16'hEFAC,4);
TASK_PP(16'hEFAD,4);
TASK_PP(16'hEFAE,4);
TASK_PP(16'hEFAF,4);
TASK_PP(16'hEFB0,4);
TASK_PP(16'hEFB1,4);
TASK_PP(16'hEFB2,4);
TASK_PP(16'hEFB3,4);
TASK_PP(16'hEFB4,4);
TASK_PP(16'hEFB5,4);
TASK_PP(16'hEFB6,4);
TASK_PP(16'hEFB7,4);
TASK_PP(16'hEFB8,4);
TASK_PP(16'hEFB9,4);
TASK_PP(16'hEFBA,4);
TASK_PP(16'hEFBB,4);
TASK_PP(16'hEFBC,4);
TASK_PP(16'hEFBD,4);
TASK_PP(16'hEFBE,4);
TASK_PP(16'hEFBF,4);
TASK_PP(16'hEFC0,4);
TASK_PP(16'hEFC1,4);
TASK_PP(16'hEFC2,4);
TASK_PP(16'hEFC3,4);
TASK_PP(16'hEFC4,4);
TASK_PP(16'hEFC5,4);
TASK_PP(16'hEFC6,4);
TASK_PP(16'hEFC7,4);
TASK_PP(16'hEFC8,4);
TASK_PP(16'hEFC9,4);
TASK_PP(16'hEFCA,4);
TASK_PP(16'hEFCB,4);
TASK_PP(16'hEFCC,4);
TASK_PP(16'hEFCD,4);
TASK_PP(16'hEFCE,4);
TASK_PP(16'hEFCF,4);
TASK_PP(16'hEFD0,4);
TASK_PP(16'hEFD1,4);
TASK_PP(16'hEFD2,4);
TASK_PP(16'hEFD3,4);
TASK_PP(16'hEFD4,4);
TASK_PP(16'hEFD5,4);
TASK_PP(16'hEFD6,4);
TASK_PP(16'hEFD7,4);
TASK_PP(16'hEFD8,4);
TASK_PP(16'hEFD9,4);
TASK_PP(16'hEFDA,4);
TASK_PP(16'hEFDB,4);
TASK_PP(16'hEFDC,4);
TASK_PP(16'hEFDD,4);
TASK_PP(16'hEFDE,4);
TASK_PP(16'hEFDF,4);
TASK_PP(16'hEFE0,4);
TASK_PP(16'hEFE1,4);
TASK_PP(16'hEFE2,4);
TASK_PP(16'hEFE3,4);
TASK_PP(16'hEFE4,4);
TASK_PP(16'hEFE5,4);
TASK_PP(16'hEFE6,4);
TASK_PP(16'hEFE7,4);
TASK_PP(16'hEFE8,4);
TASK_PP(16'hEFE9,4);
TASK_PP(16'hEFEA,4);
TASK_PP(16'hEFEB,4);
TASK_PP(16'hEFEC,4);
TASK_PP(16'hEFED,4);
TASK_PP(16'hEFEE,4);
TASK_PP(16'hEFEF,4);
TASK_PP(16'hEFF0,4);
TASK_PP(16'hEFF1,4);
TASK_PP(16'hEFF2,4);
TASK_PP(16'hEFF3,4);
TASK_PP(16'hEFF4,4);
TASK_PP(16'hEFF5,4);
TASK_PP(16'hEFF6,4);
TASK_PP(16'hEFF7,4);
TASK_PP(16'hEFF8,4);
TASK_PP(16'hEFF9,4);
TASK_PP(16'hEFFA,4);
TASK_PP(16'hEFFB,4);
TASK_PP(16'hEFFC,4);
TASK_PP(16'hEFFD,4);
TASK_PP(16'hEFFE,4);
TASK_PP(16'hEFFF,4);
TASK_PP(16'hF000,4);
TASK_PP(16'hF001,4);
TASK_PP(16'hF002,4);
TASK_PP(16'hF003,4);
TASK_PP(16'hF004,4);
TASK_PP(16'hF005,4);
TASK_PP(16'hF006,4);
TASK_PP(16'hF007,4);
TASK_PP(16'hF008,4);
TASK_PP(16'hF009,4);
TASK_PP(16'hF00A,4);
TASK_PP(16'hF00B,4);
TASK_PP(16'hF00C,4);
TASK_PP(16'hF00D,4);
TASK_PP(16'hF00E,4);
TASK_PP(16'hF00F,4);
TASK_PP(16'hF010,4);
TASK_PP(16'hF011,4);
TASK_PP(16'hF012,4);
TASK_PP(16'hF013,4);
TASK_PP(16'hF014,4);
TASK_PP(16'hF015,4);
TASK_PP(16'hF016,4);
TASK_PP(16'hF017,4);
TASK_PP(16'hF018,4);
TASK_PP(16'hF019,4);
TASK_PP(16'hF01A,4);
TASK_PP(16'hF01B,4);
TASK_PP(16'hF01C,4);
TASK_PP(16'hF01D,4);
TASK_PP(16'hF01E,4);
TASK_PP(16'hF01F,4);
TASK_PP(16'hF020,4);
TASK_PP(16'hF021,4);
TASK_PP(16'hF022,4);
TASK_PP(16'hF023,4);
TASK_PP(16'hF024,4);
TASK_PP(16'hF025,4);
TASK_PP(16'hF026,4);
TASK_PP(16'hF027,4);
TASK_PP(16'hF028,4);
TASK_PP(16'hF029,4);
TASK_PP(16'hF02A,4);
TASK_PP(16'hF02B,4);
TASK_PP(16'hF02C,4);
TASK_PP(16'hF02D,4);
TASK_PP(16'hF02E,4);
TASK_PP(16'hF02F,4);
TASK_PP(16'hF030,4);
TASK_PP(16'hF031,4);
TASK_PP(16'hF032,4);
TASK_PP(16'hF033,4);
TASK_PP(16'hF034,4);
TASK_PP(16'hF035,4);
TASK_PP(16'hF036,4);
TASK_PP(16'hF037,4);
TASK_PP(16'hF038,4);
TASK_PP(16'hF039,4);
TASK_PP(16'hF03A,4);
TASK_PP(16'hF03B,4);
TASK_PP(16'hF03C,4);
TASK_PP(16'hF03D,4);
TASK_PP(16'hF03E,4);
TASK_PP(16'hF03F,4);
TASK_PP(16'hF040,4);
TASK_PP(16'hF041,4);
TASK_PP(16'hF042,4);
TASK_PP(16'hF043,4);
TASK_PP(16'hF044,4);
TASK_PP(16'hF045,4);
TASK_PP(16'hF046,4);
TASK_PP(16'hF047,4);
TASK_PP(16'hF048,4);
TASK_PP(16'hF049,4);
TASK_PP(16'hF04A,4);
TASK_PP(16'hF04B,4);
TASK_PP(16'hF04C,4);
TASK_PP(16'hF04D,4);
TASK_PP(16'hF04E,4);
TASK_PP(16'hF04F,4);
TASK_PP(16'hF050,4);
TASK_PP(16'hF051,4);
TASK_PP(16'hF052,4);
TASK_PP(16'hF053,4);
TASK_PP(16'hF054,4);
TASK_PP(16'hF055,4);
TASK_PP(16'hF056,4);
TASK_PP(16'hF057,4);
TASK_PP(16'hF058,4);
TASK_PP(16'hF059,4);
TASK_PP(16'hF05A,4);
TASK_PP(16'hF05B,4);
TASK_PP(16'hF05C,4);
TASK_PP(16'hF05D,4);
TASK_PP(16'hF05E,4);
TASK_PP(16'hF05F,4);
TASK_PP(16'hF060,4);
TASK_PP(16'hF061,4);
TASK_PP(16'hF062,4);
TASK_PP(16'hF063,4);
TASK_PP(16'hF064,4);
TASK_PP(16'hF065,4);
TASK_PP(16'hF066,4);
TASK_PP(16'hF067,4);
TASK_PP(16'hF068,4);
TASK_PP(16'hF069,4);
TASK_PP(16'hF06A,4);
TASK_PP(16'hF06B,4);
TASK_PP(16'hF06C,4);
TASK_PP(16'hF06D,4);
TASK_PP(16'hF06E,4);
TASK_PP(16'hF06F,4);
TASK_PP(16'hF070,4);
TASK_PP(16'hF071,4);
TASK_PP(16'hF072,4);
TASK_PP(16'hF073,4);
TASK_PP(16'hF074,4);
TASK_PP(16'hF075,4);
TASK_PP(16'hF076,4);
TASK_PP(16'hF077,4);
TASK_PP(16'hF078,4);
TASK_PP(16'hF079,4);
TASK_PP(16'hF07A,4);
TASK_PP(16'hF07B,4);
TASK_PP(16'hF07C,4);
TASK_PP(16'hF07D,4);
TASK_PP(16'hF07E,4);
TASK_PP(16'hF07F,4);
TASK_PP(16'hF080,4);
TASK_PP(16'hF081,4);
TASK_PP(16'hF082,4);
TASK_PP(16'hF083,4);
TASK_PP(16'hF084,4);
TASK_PP(16'hF085,4);
TASK_PP(16'hF086,4);
TASK_PP(16'hF087,4);
TASK_PP(16'hF088,4);
TASK_PP(16'hF089,4);
TASK_PP(16'hF08A,4);
TASK_PP(16'hF08B,4);
TASK_PP(16'hF08C,4);
TASK_PP(16'hF08D,4);
TASK_PP(16'hF08E,4);
TASK_PP(16'hF08F,4);
TASK_PP(16'hF090,4);
TASK_PP(16'hF091,4);
TASK_PP(16'hF092,4);
TASK_PP(16'hF093,4);
TASK_PP(16'hF094,4);
TASK_PP(16'hF095,4);
TASK_PP(16'hF096,4);
TASK_PP(16'hF097,4);
TASK_PP(16'hF098,4);
TASK_PP(16'hF099,4);
TASK_PP(16'hF09A,4);
TASK_PP(16'hF09B,4);
TASK_PP(16'hF09C,4);
TASK_PP(16'hF09D,4);
TASK_PP(16'hF09E,4);
TASK_PP(16'hF09F,4);
TASK_PP(16'hF0A0,4);
TASK_PP(16'hF0A1,4);
TASK_PP(16'hF0A2,4);
TASK_PP(16'hF0A3,4);
TASK_PP(16'hF0A4,4);
TASK_PP(16'hF0A5,4);
TASK_PP(16'hF0A6,4);
TASK_PP(16'hF0A7,4);
TASK_PP(16'hF0A8,4);
TASK_PP(16'hF0A9,4);
TASK_PP(16'hF0AA,4);
TASK_PP(16'hF0AB,4);
TASK_PP(16'hF0AC,4);
TASK_PP(16'hF0AD,4);
TASK_PP(16'hF0AE,4);
TASK_PP(16'hF0AF,4);
TASK_PP(16'hF0B0,4);
TASK_PP(16'hF0B1,4);
TASK_PP(16'hF0B2,4);
TASK_PP(16'hF0B3,4);
TASK_PP(16'hF0B4,4);
TASK_PP(16'hF0B5,4);
TASK_PP(16'hF0B6,4);
TASK_PP(16'hF0B7,4);
TASK_PP(16'hF0B8,4);
TASK_PP(16'hF0B9,4);
TASK_PP(16'hF0BA,4);
TASK_PP(16'hF0BB,4);
TASK_PP(16'hF0BC,4);
TASK_PP(16'hF0BD,4);
TASK_PP(16'hF0BE,4);
TASK_PP(16'hF0BF,4);
TASK_PP(16'hF0C0,4);
TASK_PP(16'hF0C1,4);
TASK_PP(16'hF0C2,4);
TASK_PP(16'hF0C3,4);
TASK_PP(16'hF0C4,4);
TASK_PP(16'hF0C5,4);
TASK_PP(16'hF0C6,4);
TASK_PP(16'hF0C7,4);
TASK_PP(16'hF0C8,4);
TASK_PP(16'hF0C9,4);
TASK_PP(16'hF0CA,4);
TASK_PP(16'hF0CB,4);
TASK_PP(16'hF0CC,4);
TASK_PP(16'hF0CD,4);
TASK_PP(16'hF0CE,4);
TASK_PP(16'hF0CF,4);
TASK_PP(16'hF0D0,4);
TASK_PP(16'hF0D1,4);
TASK_PP(16'hF0D2,4);
TASK_PP(16'hF0D3,4);
TASK_PP(16'hF0D4,4);
TASK_PP(16'hF0D5,4);
TASK_PP(16'hF0D6,4);
TASK_PP(16'hF0D7,4);
TASK_PP(16'hF0D8,4);
TASK_PP(16'hF0D9,4);
TASK_PP(16'hF0DA,4);
TASK_PP(16'hF0DB,4);
TASK_PP(16'hF0DC,4);
TASK_PP(16'hF0DD,4);
TASK_PP(16'hF0DE,4);
TASK_PP(16'hF0DF,4);
TASK_PP(16'hF0E0,4);
TASK_PP(16'hF0E1,4);
TASK_PP(16'hF0E2,4);
TASK_PP(16'hF0E3,4);
TASK_PP(16'hF0E4,4);
TASK_PP(16'hF0E5,4);
TASK_PP(16'hF0E6,4);
TASK_PP(16'hF0E7,4);
TASK_PP(16'hF0E8,4);
TASK_PP(16'hF0E9,4);
TASK_PP(16'hF0EA,4);
TASK_PP(16'hF0EB,4);
TASK_PP(16'hF0EC,4);
TASK_PP(16'hF0ED,4);
TASK_PP(16'hF0EE,4);
TASK_PP(16'hF0EF,4);
TASK_PP(16'hF0F0,4);
TASK_PP(16'hF0F1,4);
TASK_PP(16'hF0F2,4);
TASK_PP(16'hF0F3,4);
TASK_PP(16'hF0F4,4);
TASK_PP(16'hF0F5,4);
TASK_PP(16'hF0F6,4);
TASK_PP(16'hF0F7,4);
TASK_PP(16'hF0F8,4);
TASK_PP(16'hF0F9,4);
TASK_PP(16'hF0FA,4);
TASK_PP(16'hF0FB,4);
TASK_PP(16'hF0FC,4);
TASK_PP(16'hF0FD,4);
TASK_PP(16'hF0FE,4);
TASK_PP(16'hF0FF,4);
TASK_PP(16'hF100,4);
TASK_PP(16'hF101,4);
TASK_PP(16'hF102,4);
TASK_PP(16'hF103,4);
TASK_PP(16'hF104,4);
TASK_PP(16'hF105,4);
TASK_PP(16'hF106,4);
TASK_PP(16'hF107,4);
TASK_PP(16'hF108,4);
TASK_PP(16'hF109,4);
TASK_PP(16'hF10A,4);
TASK_PP(16'hF10B,4);
TASK_PP(16'hF10C,4);
TASK_PP(16'hF10D,4);
TASK_PP(16'hF10E,4);
TASK_PP(16'hF10F,4);
TASK_PP(16'hF110,4);
TASK_PP(16'hF111,4);
TASK_PP(16'hF112,4);
TASK_PP(16'hF113,4);
TASK_PP(16'hF114,4);
TASK_PP(16'hF115,4);
TASK_PP(16'hF116,4);
TASK_PP(16'hF117,4);
TASK_PP(16'hF118,4);
TASK_PP(16'hF119,4);
TASK_PP(16'hF11A,4);
TASK_PP(16'hF11B,4);
TASK_PP(16'hF11C,4);
TASK_PP(16'hF11D,4);
TASK_PP(16'hF11E,4);
TASK_PP(16'hF11F,4);
TASK_PP(16'hF120,4);
TASK_PP(16'hF121,4);
TASK_PP(16'hF122,4);
TASK_PP(16'hF123,4);
TASK_PP(16'hF124,4);
TASK_PP(16'hF125,4);
TASK_PP(16'hF126,4);
TASK_PP(16'hF127,4);
TASK_PP(16'hF128,4);
TASK_PP(16'hF129,4);
TASK_PP(16'hF12A,4);
TASK_PP(16'hF12B,4);
TASK_PP(16'hF12C,4);
TASK_PP(16'hF12D,4);
TASK_PP(16'hF12E,4);
TASK_PP(16'hF12F,4);
TASK_PP(16'hF130,4);
TASK_PP(16'hF131,4);
TASK_PP(16'hF132,4);
TASK_PP(16'hF133,4);
TASK_PP(16'hF134,4);
TASK_PP(16'hF135,4);
TASK_PP(16'hF136,4);
TASK_PP(16'hF137,4);
TASK_PP(16'hF138,4);
TASK_PP(16'hF139,4);
TASK_PP(16'hF13A,4);
TASK_PP(16'hF13B,4);
TASK_PP(16'hF13C,4);
TASK_PP(16'hF13D,4);
TASK_PP(16'hF13E,4);
TASK_PP(16'hF13F,4);
TASK_PP(16'hF140,4);
TASK_PP(16'hF141,4);
TASK_PP(16'hF142,4);
TASK_PP(16'hF143,4);
TASK_PP(16'hF144,4);
TASK_PP(16'hF145,4);
TASK_PP(16'hF146,4);
TASK_PP(16'hF147,4);
TASK_PP(16'hF148,4);
TASK_PP(16'hF149,4);
TASK_PP(16'hF14A,4);
TASK_PP(16'hF14B,4);
TASK_PP(16'hF14C,4);
TASK_PP(16'hF14D,4);
TASK_PP(16'hF14E,4);
TASK_PP(16'hF14F,4);
TASK_PP(16'hF150,4);
TASK_PP(16'hF151,4);
TASK_PP(16'hF152,4);
TASK_PP(16'hF153,4);
TASK_PP(16'hF154,4);
TASK_PP(16'hF155,4);
TASK_PP(16'hF156,4);
TASK_PP(16'hF157,4);
TASK_PP(16'hF158,4);
TASK_PP(16'hF159,4);
TASK_PP(16'hF15A,4);
TASK_PP(16'hF15B,4);
TASK_PP(16'hF15C,4);
TASK_PP(16'hF15D,4);
TASK_PP(16'hF15E,4);
TASK_PP(16'hF15F,4);
TASK_PP(16'hF160,4);
TASK_PP(16'hF161,4);
TASK_PP(16'hF162,4);
TASK_PP(16'hF163,4);
TASK_PP(16'hF164,4);
TASK_PP(16'hF165,4);
TASK_PP(16'hF166,4);
TASK_PP(16'hF167,4);
TASK_PP(16'hF168,4);
TASK_PP(16'hF169,4);
TASK_PP(16'hF16A,4);
TASK_PP(16'hF16B,4);
TASK_PP(16'hF16C,4);
TASK_PP(16'hF16D,4);
TASK_PP(16'hF16E,4);
TASK_PP(16'hF16F,4);
TASK_PP(16'hF170,4);
TASK_PP(16'hF171,4);
TASK_PP(16'hF172,4);
TASK_PP(16'hF173,4);
TASK_PP(16'hF174,4);
TASK_PP(16'hF175,4);
TASK_PP(16'hF176,4);
TASK_PP(16'hF177,4);
TASK_PP(16'hF178,4);
TASK_PP(16'hF179,4);
TASK_PP(16'hF17A,4);
TASK_PP(16'hF17B,4);
TASK_PP(16'hF17C,4);
TASK_PP(16'hF17D,4);
TASK_PP(16'hF17E,4);
TASK_PP(16'hF17F,4);
TASK_PP(16'hF180,4);
TASK_PP(16'hF181,4);
TASK_PP(16'hF182,4);
TASK_PP(16'hF183,4);
TASK_PP(16'hF184,4);
TASK_PP(16'hF185,4);
TASK_PP(16'hF186,4);
TASK_PP(16'hF187,4);
TASK_PP(16'hF188,4);
TASK_PP(16'hF189,4);
TASK_PP(16'hF18A,4);
TASK_PP(16'hF18B,4);
TASK_PP(16'hF18C,4);
TASK_PP(16'hF18D,4);
TASK_PP(16'hF18E,4);
TASK_PP(16'hF18F,4);
TASK_PP(16'hF190,4);
TASK_PP(16'hF191,4);
TASK_PP(16'hF192,4);
TASK_PP(16'hF193,4);
TASK_PP(16'hF194,4);
TASK_PP(16'hF195,4);
TASK_PP(16'hF196,4);
TASK_PP(16'hF197,4);
TASK_PP(16'hF198,4);
TASK_PP(16'hF199,4);
TASK_PP(16'hF19A,4);
TASK_PP(16'hF19B,4);
TASK_PP(16'hF19C,4);
TASK_PP(16'hF19D,4);
TASK_PP(16'hF19E,4);
TASK_PP(16'hF19F,4);
TASK_PP(16'hF1A0,4);
TASK_PP(16'hF1A1,4);
TASK_PP(16'hF1A2,4);
TASK_PP(16'hF1A3,4);
TASK_PP(16'hF1A4,4);
TASK_PP(16'hF1A5,4);
TASK_PP(16'hF1A6,4);
TASK_PP(16'hF1A7,4);
TASK_PP(16'hF1A8,4);
TASK_PP(16'hF1A9,4);
TASK_PP(16'hF1AA,4);
TASK_PP(16'hF1AB,4);
TASK_PP(16'hF1AC,4);
TASK_PP(16'hF1AD,4);
TASK_PP(16'hF1AE,4);
TASK_PP(16'hF1AF,4);
TASK_PP(16'hF1B0,4);
TASK_PP(16'hF1B1,4);
TASK_PP(16'hF1B2,4);
TASK_PP(16'hF1B3,4);
TASK_PP(16'hF1B4,4);
TASK_PP(16'hF1B5,4);
TASK_PP(16'hF1B6,4);
TASK_PP(16'hF1B7,4);
TASK_PP(16'hF1B8,4);
TASK_PP(16'hF1B9,4);
TASK_PP(16'hF1BA,4);
TASK_PP(16'hF1BB,4);
TASK_PP(16'hF1BC,4);
TASK_PP(16'hF1BD,4);
TASK_PP(16'hF1BE,4);
TASK_PP(16'hF1BF,4);
TASK_PP(16'hF1C0,4);
TASK_PP(16'hF1C1,4);
TASK_PP(16'hF1C2,4);
TASK_PP(16'hF1C3,4);
TASK_PP(16'hF1C4,4);
TASK_PP(16'hF1C5,4);
TASK_PP(16'hF1C6,4);
TASK_PP(16'hF1C7,4);
TASK_PP(16'hF1C8,4);
TASK_PP(16'hF1C9,4);
TASK_PP(16'hF1CA,4);
TASK_PP(16'hF1CB,4);
TASK_PP(16'hF1CC,4);
TASK_PP(16'hF1CD,4);
TASK_PP(16'hF1CE,4);
TASK_PP(16'hF1CF,4);
TASK_PP(16'hF1D0,4);
TASK_PP(16'hF1D1,4);
TASK_PP(16'hF1D2,4);
TASK_PP(16'hF1D3,4);
TASK_PP(16'hF1D4,4);
TASK_PP(16'hF1D5,4);
TASK_PP(16'hF1D6,4);
TASK_PP(16'hF1D7,4);
TASK_PP(16'hF1D8,4);
TASK_PP(16'hF1D9,4);
TASK_PP(16'hF1DA,4);
TASK_PP(16'hF1DB,4);
TASK_PP(16'hF1DC,4);
TASK_PP(16'hF1DD,4);
TASK_PP(16'hF1DE,4);
TASK_PP(16'hF1DF,4);
TASK_PP(16'hF1E0,4);
TASK_PP(16'hF1E1,4);
TASK_PP(16'hF1E2,4);
TASK_PP(16'hF1E3,4);
TASK_PP(16'hF1E4,4);
TASK_PP(16'hF1E5,4);
TASK_PP(16'hF1E6,4);
TASK_PP(16'hF1E7,4);
TASK_PP(16'hF1E8,4);
TASK_PP(16'hF1E9,4);
TASK_PP(16'hF1EA,4);
TASK_PP(16'hF1EB,4);
TASK_PP(16'hF1EC,4);
TASK_PP(16'hF1ED,4);
TASK_PP(16'hF1EE,4);
TASK_PP(16'hF1EF,4);
TASK_PP(16'hF1F0,4);
TASK_PP(16'hF1F1,4);
TASK_PP(16'hF1F2,4);
TASK_PP(16'hF1F3,4);
TASK_PP(16'hF1F4,4);
TASK_PP(16'hF1F5,4);
TASK_PP(16'hF1F6,4);
TASK_PP(16'hF1F7,4);
TASK_PP(16'hF1F8,4);
TASK_PP(16'hF1F9,4);
TASK_PP(16'hF1FA,4);
TASK_PP(16'hF1FB,4);
TASK_PP(16'hF1FC,4);
TASK_PP(16'hF1FD,4);
TASK_PP(16'hF1FE,4);
TASK_PP(16'hF1FF,4);
TASK_PP(16'hF200,4);
TASK_PP(16'hF201,4);
TASK_PP(16'hF202,4);
TASK_PP(16'hF203,4);
TASK_PP(16'hF204,4);
TASK_PP(16'hF205,4);
TASK_PP(16'hF206,4);
TASK_PP(16'hF207,4);
TASK_PP(16'hF208,4);
TASK_PP(16'hF209,4);
TASK_PP(16'hF20A,4);
TASK_PP(16'hF20B,4);
TASK_PP(16'hF20C,4);
TASK_PP(16'hF20D,4);
TASK_PP(16'hF20E,4);
TASK_PP(16'hF20F,4);
TASK_PP(16'hF210,4);
TASK_PP(16'hF211,4);
TASK_PP(16'hF212,4);
TASK_PP(16'hF213,4);
TASK_PP(16'hF214,4);
TASK_PP(16'hF215,4);
TASK_PP(16'hF216,4);
TASK_PP(16'hF217,4);
TASK_PP(16'hF218,4);
TASK_PP(16'hF219,4);
TASK_PP(16'hF21A,4);
TASK_PP(16'hF21B,4);
TASK_PP(16'hF21C,4);
TASK_PP(16'hF21D,4);
TASK_PP(16'hF21E,4);
TASK_PP(16'hF21F,4);
TASK_PP(16'hF220,4);
TASK_PP(16'hF221,4);
TASK_PP(16'hF222,4);
TASK_PP(16'hF223,4);
TASK_PP(16'hF224,4);
TASK_PP(16'hF225,4);
TASK_PP(16'hF226,4);
TASK_PP(16'hF227,4);
TASK_PP(16'hF228,4);
TASK_PP(16'hF229,4);
TASK_PP(16'hF22A,4);
TASK_PP(16'hF22B,4);
TASK_PP(16'hF22C,4);
TASK_PP(16'hF22D,4);
TASK_PP(16'hF22E,4);
TASK_PP(16'hF22F,4);
TASK_PP(16'hF230,4);
TASK_PP(16'hF231,4);
TASK_PP(16'hF232,4);
TASK_PP(16'hF233,4);
TASK_PP(16'hF234,4);
TASK_PP(16'hF235,4);
TASK_PP(16'hF236,4);
TASK_PP(16'hF237,4);
TASK_PP(16'hF238,4);
TASK_PP(16'hF239,4);
TASK_PP(16'hF23A,4);
TASK_PP(16'hF23B,4);
TASK_PP(16'hF23C,4);
TASK_PP(16'hF23D,4);
TASK_PP(16'hF23E,4);
TASK_PP(16'hF23F,4);
TASK_PP(16'hF240,4);
TASK_PP(16'hF241,4);
TASK_PP(16'hF242,4);
TASK_PP(16'hF243,4);
TASK_PP(16'hF244,4);
TASK_PP(16'hF245,4);
TASK_PP(16'hF246,4);
TASK_PP(16'hF247,4);
TASK_PP(16'hF248,4);
TASK_PP(16'hF249,4);
TASK_PP(16'hF24A,4);
TASK_PP(16'hF24B,4);
TASK_PP(16'hF24C,4);
TASK_PP(16'hF24D,4);
TASK_PP(16'hF24E,4);
TASK_PP(16'hF24F,4);
TASK_PP(16'hF250,4);
TASK_PP(16'hF251,4);
TASK_PP(16'hF252,4);
TASK_PP(16'hF253,4);
TASK_PP(16'hF254,4);
TASK_PP(16'hF255,4);
TASK_PP(16'hF256,4);
TASK_PP(16'hF257,4);
TASK_PP(16'hF258,4);
TASK_PP(16'hF259,4);
TASK_PP(16'hF25A,4);
TASK_PP(16'hF25B,4);
TASK_PP(16'hF25C,4);
TASK_PP(16'hF25D,4);
TASK_PP(16'hF25E,4);
TASK_PP(16'hF25F,4);
TASK_PP(16'hF260,4);
TASK_PP(16'hF261,4);
TASK_PP(16'hF262,4);
TASK_PP(16'hF263,4);
TASK_PP(16'hF264,4);
TASK_PP(16'hF265,4);
TASK_PP(16'hF266,4);
TASK_PP(16'hF267,4);
TASK_PP(16'hF268,4);
TASK_PP(16'hF269,4);
TASK_PP(16'hF26A,4);
TASK_PP(16'hF26B,4);
TASK_PP(16'hF26C,4);
TASK_PP(16'hF26D,4);
TASK_PP(16'hF26E,4);
TASK_PP(16'hF26F,4);
TASK_PP(16'hF270,4);
TASK_PP(16'hF271,4);
TASK_PP(16'hF272,4);
TASK_PP(16'hF273,4);
TASK_PP(16'hF274,4);
TASK_PP(16'hF275,4);
TASK_PP(16'hF276,4);
TASK_PP(16'hF277,4);
TASK_PP(16'hF278,4);
TASK_PP(16'hF279,4);
TASK_PP(16'hF27A,4);
TASK_PP(16'hF27B,4);
TASK_PP(16'hF27C,4);
TASK_PP(16'hF27D,4);
TASK_PP(16'hF27E,4);
TASK_PP(16'hF27F,4);
TASK_PP(16'hF280,4);
TASK_PP(16'hF281,4);
TASK_PP(16'hF282,4);
TASK_PP(16'hF283,4);
TASK_PP(16'hF284,4);
TASK_PP(16'hF285,4);
TASK_PP(16'hF286,4);
TASK_PP(16'hF287,4);
TASK_PP(16'hF288,4);
TASK_PP(16'hF289,4);
TASK_PP(16'hF28A,4);
TASK_PP(16'hF28B,4);
TASK_PP(16'hF28C,4);
TASK_PP(16'hF28D,4);
TASK_PP(16'hF28E,4);
TASK_PP(16'hF28F,4);
TASK_PP(16'hF290,4);
TASK_PP(16'hF291,4);
TASK_PP(16'hF292,4);
TASK_PP(16'hF293,4);
TASK_PP(16'hF294,4);
TASK_PP(16'hF295,4);
TASK_PP(16'hF296,4);
TASK_PP(16'hF297,4);
TASK_PP(16'hF298,4);
TASK_PP(16'hF299,4);
TASK_PP(16'hF29A,4);
TASK_PP(16'hF29B,4);
TASK_PP(16'hF29C,4);
TASK_PP(16'hF29D,4);
TASK_PP(16'hF29E,4);
TASK_PP(16'hF29F,4);
TASK_PP(16'hF2A0,4);
TASK_PP(16'hF2A1,4);
TASK_PP(16'hF2A2,4);
TASK_PP(16'hF2A3,4);
TASK_PP(16'hF2A4,4);
TASK_PP(16'hF2A5,4);
TASK_PP(16'hF2A6,4);
TASK_PP(16'hF2A7,4);
TASK_PP(16'hF2A8,4);
TASK_PP(16'hF2A9,4);
TASK_PP(16'hF2AA,4);
TASK_PP(16'hF2AB,4);
TASK_PP(16'hF2AC,4);
TASK_PP(16'hF2AD,4);
TASK_PP(16'hF2AE,4);
TASK_PP(16'hF2AF,4);
TASK_PP(16'hF2B0,4);
TASK_PP(16'hF2B1,4);
TASK_PP(16'hF2B2,4);
TASK_PP(16'hF2B3,4);
TASK_PP(16'hF2B4,4);
TASK_PP(16'hF2B5,4);
TASK_PP(16'hF2B6,4);
TASK_PP(16'hF2B7,4);
TASK_PP(16'hF2B8,4);
TASK_PP(16'hF2B9,4);
TASK_PP(16'hF2BA,4);
TASK_PP(16'hF2BB,4);
TASK_PP(16'hF2BC,4);
TASK_PP(16'hF2BD,4);
TASK_PP(16'hF2BE,4);
TASK_PP(16'hF2BF,4);
TASK_PP(16'hF2C0,4);
TASK_PP(16'hF2C1,4);
TASK_PP(16'hF2C2,4);
TASK_PP(16'hF2C3,4);
TASK_PP(16'hF2C4,4);
TASK_PP(16'hF2C5,4);
TASK_PP(16'hF2C6,4);
TASK_PP(16'hF2C7,4);
TASK_PP(16'hF2C8,4);
TASK_PP(16'hF2C9,4);
TASK_PP(16'hF2CA,4);
TASK_PP(16'hF2CB,4);
TASK_PP(16'hF2CC,4);
TASK_PP(16'hF2CD,4);
TASK_PP(16'hF2CE,4);
TASK_PP(16'hF2CF,4);
TASK_PP(16'hF2D0,4);
TASK_PP(16'hF2D1,4);
TASK_PP(16'hF2D2,4);
TASK_PP(16'hF2D3,4);
TASK_PP(16'hF2D4,4);
TASK_PP(16'hF2D5,4);
TASK_PP(16'hF2D6,4);
TASK_PP(16'hF2D7,4);
TASK_PP(16'hF2D8,4);
TASK_PP(16'hF2D9,4);
TASK_PP(16'hF2DA,4);
TASK_PP(16'hF2DB,4);
TASK_PP(16'hF2DC,4);
TASK_PP(16'hF2DD,4);
TASK_PP(16'hF2DE,4);
TASK_PP(16'hF2DF,4);
TASK_PP(16'hF2E0,4);
TASK_PP(16'hF2E1,4);
TASK_PP(16'hF2E2,4);
TASK_PP(16'hF2E3,4);
TASK_PP(16'hF2E4,4);
TASK_PP(16'hF2E5,4);
TASK_PP(16'hF2E6,4);
TASK_PP(16'hF2E7,4);
TASK_PP(16'hF2E8,4);
TASK_PP(16'hF2E9,4);
TASK_PP(16'hF2EA,4);
TASK_PP(16'hF2EB,4);
TASK_PP(16'hF2EC,4);
TASK_PP(16'hF2ED,4);
TASK_PP(16'hF2EE,4);
TASK_PP(16'hF2EF,4);
TASK_PP(16'hF2F0,4);
TASK_PP(16'hF2F1,4);
TASK_PP(16'hF2F2,4);
TASK_PP(16'hF2F3,4);
TASK_PP(16'hF2F4,4);
TASK_PP(16'hF2F5,4);
TASK_PP(16'hF2F6,4);
TASK_PP(16'hF2F7,4);
TASK_PP(16'hF2F8,4);
TASK_PP(16'hF2F9,4);
TASK_PP(16'hF2FA,4);
TASK_PP(16'hF2FB,4);
TASK_PP(16'hF2FC,4);
TASK_PP(16'hF2FD,4);
TASK_PP(16'hF2FE,4);
TASK_PP(16'hF2FF,4);
TASK_PP(16'hF300,4);
TASK_PP(16'hF301,4);
TASK_PP(16'hF302,4);
TASK_PP(16'hF303,4);
TASK_PP(16'hF304,4);
TASK_PP(16'hF305,4);
TASK_PP(16'hF306,4);
TASK_PP(16'hF307,4);
TASK_PP(16'hF308,4);
TASK_PP(16'hF309,4);
TASK_PP(16'hF30A,4);
TASK_PP(16'hF30B,4);
TASK_PP(16'hF30C,4);
TASK_PP(16'hF30D,4);
TASK_PP(16'hF30E,4);
TASK_PP(16'hF30F,4);
TASK_PP(16'hF310,4);
TASK_PP(16'hF311,4);
TASK_PP(16'hF312,4);
TASK_PP(16'hF313,4);
TASK_PP(16'hF314,4);
TASK_PP(16'hF315,4);
TASK_PP(16'hF316,4);
TASK_PP(16'hF317,4);
TASK_PP(16'hF318,4);
TASK_PP(16'hF319,4);
TASK_PP(16'hF31A,4);
TASK_PP(16'hF31B,4);
TASK_PP(16'hF31C,4);
TASK_PP(16'hF31D,4);
TASK_PP(16'hF31E,4);
TASK_PP(16'hF31F,4);
TASK_PP(16'hF320,4);
TASK_PP(16'hF321,4);
TASK_PP(16'hF322,4);
TASK_PP(16'hF323,4);
TASK_PP(16'hF324,4);
TASK_PP(16'hF325,4);
TASK_PP(16'hF326,4);
TASK_PP(16'hF327,4);
TASK_PP(16'hF328,4);
TASK_PP(16'hF329,4);
TASK_PP(16'hF32A,4);
TASK_PP(16'hF32B,4);
TASK_PP(16'hF32C,4);
TASK_PP(16'hF32D,4);
TASK_PP(16'hF32E,4);
TASK_PP(16'hF32F,4);
TASK_PP(16'hF330,4);
TASK_PP(16'hF331,4);
TASK_PP(16'hF332,4);
TASK_PP(16'hF333,4);
TASK_PP(16'hF334,4);
TASK_PP(16'hF335,4);
TASK_PP(16'hF336,4);
TASK_PP(16'hF337,4);
TASK_PP(16'hF338,4);
TASK_PP(16'hF339,4);
TASK_PP(16'hF33A,4);
TASK_PP(16'hF33B,4);
TASK_PP(16'hF33C,4);
TASK_PP(16'hF33D,4);
TASK_PP(16'hF33E,4);
TASK_PP(16'hF33F,4);
TASK_PP(16'hF340,4);
TASK_PP(16'hF341,4);
TASK_PP(16'hF342,4);
TASK_PP(16'hF343,4);
TASK_PP(16'hF344,4);
TASK_PP(16'hF345,4);
TASK_PP(16'hF346,4);
TASK_PP(16'hF347,4);
TASK_PP(16'hF348,4);
TASK_PP(16'hF349,4);
TASK_PP(16'hF34A,4);
TASK_PP(16'hF34B,4);
TASK_PP(16'hF34C,4);
TASK_PP(16'hF34D,4);
TASK_PP(16'hF34E,4);
TASK_PP(16'hF34F,4);
TASK_PP(16'hF350,4);
TASK_PP(16'hF351,4);
TASK_PP(16'hF352,4);
TASK_PP(16'hF353,4);
TASK_PP(16'hF354,4);
TASK_PP(16'hF355,4);
TASK_PP(16'hF356,4);
TASK_PP(16'hF357,4);
TASK_PP(16'hF358,4);
TASK_PP(16'hF359,4);
TASK_PP(16'hF35A,4);
TASK_PP(16'hF35B,4);
TASK_PP(16'hF35C,4);
TASK_PP(16'hF35D,4);
TASK_PP(16'hF35E,4);
TASK_PP(16'hF35F,4);
TASK_PP(16'hF360,4);
TASK_PP(16'hF361,4);
TASK_PP(16'hF362,4);
TASK_PP(16'hF363,4);
TASK_PP(16'hF364,4);
TASK_PP(16'hF365,4);
TASK_PP(16'hF366,4);
TASK_PP(16'hF367,4);
TASK_PP(16'hF368,4);
TASK_PP(16'hF369,4);
TASK_PP(16'hF36A,4);
TASK_PP(16'hF36B,4);
TASK_PP(16'hF36C,4);
TASK_PP(16'hF36D,4);
TASK_PP(16'hF36E,4);
TASK_PP(16'hF36F,4);
TASK_PP(16'hF370,4);
TASK_PP(16'hF371,4);
TASK_PP(16'hF372,4);
TASK_PP(16'hF373,4);
TASK_PP(16'hF374,4);
TASK_PP(16'hF375,4);
TASK_PP(16'hF376,4);
TASK_PP(16'hF377,4);
TASK_PP(16'hF378,4);
TASK_PP(16'hF379,4);
TASK_PP(16'hF37A,4);
TASK_PP(16'hF37B,4);
TASK_PP(16'hF37C,4);
TASK_PP(16'hF37D,4);
TASK_PP(16'hF37E,4);
TASK_PP(16'hF37F,4);
TASK_PP(16'hF380,4);
TASK_PP(16'hF381,4);
TASK_PP(16'hF382,4);
TASK_PP(16'hF383,4);
TASK_PP(16'hF384,4);
TASK_PP(16'hF385,4);
TASK_PP(16'hF386,4);
TASK_PP(16'hF387,4);
TASK_PP(16'hF388,4);
TASK_PP(16'hF389,4);
TASK_PP(16'hF38A,4);
TASK_PP(16'hF38B,4);
TASK_PP(16'hF38C,4);
TASK_PP(16'hF38D,4);
TASK_PP(16'hF38E,4);
TASK_PP(16'hF38F,4);
TASK_PP(16'hF390,4);
TASK_PP(16'hF391,4);
TASK_PP(16'hF392,4);
TASK_PP(16'hF393,4);
TASK_PP(16'hF394,4);
TASK_PP(16'hF395,4);
TASK_PP(16'hF396,4);
TASK_PP(16'hF397,4);
TASK_PP(16'hF398,4);
TASK_PP(16'hF399,4);
TASK_PP(16'hF39A,4);
TASK_PP(16'hF39B,4);
TASK_PP(16'hF39C,4);
TASK_PP(16'hF39D,4);
TASK_PP(16'hF39E,4);
TASK_PP(16'hF39F,4);
TASK_PP(16'hF3A0,4);
TASK_PP(16'hF3A1,4);
TASK_PP(16'hF3A2,4);
TASK_PP(16'hF3A3,4);
TASK_PP(16'hF3A4,4);
TASK_PP(16'hF3A5,4);
TASK_PP(16'hF3A6,4);
TASK_PP(16'hF3A7,4);
TASK_PP(16'hF3A8,4);
TASK_PP(16'hF3A9,4);
TASK_PP(16'hF3AA,4);
TASK_PP(16'hF3AB,4);
TASK_PP(16'hF3AC,4);
TASK_PP(16'hF3AD,4);
TASK_PP(16'hF3AE,4);
TASK_PP(16'hF3AF,4);
TASK_PP(16'hF3B0,4);
TASK_PP(16'hF3B1,4);
TASK_PP(16'hF3B2,4);
TASK_PP(16'hF3B3,4);
TASK_PP(16'hF3B4,4);
TASK_PP(16'hF3B5,4);
TASK_PP(16'hF3B6,4);
TASK_PP(16'hF3B7,4);
TASK_PP(16'hF3B8,4);
TASK_PP(16'hF3B9,4);
TASK_PP(16'hF3BA,4);
TASK_PP(16'hF3BB,4);
TASK_PP(16'hF3BC,4);
TASK_PP(16'hF3BD,4);
TASK_PP(16'hF3BE,4);
TASK_PP(16'hF3BF,4);
TASK_PP(16'hF3C0,4);
TASK_PP(16'hF3C1,4);
TASK_PP(16'hF3C2,4);
TASK_PP(16'hF3C3,4);
TASK_PP(16'hF3C4,4);
TASK_PP(16'hF3C5,4);
TASK_PP(16'hF3C6,4);
TASK_PP(16'hF3C7,4);
TASK_PP(16'hF3C8,4);
TASK_PP(16'hF3C9,4);
TASK_PP(16'hF3CA,4);
TASK_PP(16'hF3CB,4);
TASK_PP(16'hF3CC,4);
TASK_PP(16'hF3CD,4);
TASK_PP(16'hF3CE,4);
TASK_PP(16'hF3CF,4);
TASK_PP(16'hF3D0,4);
TASK_PP(16'hF3D1,4);
TASK_PP(16'hF3D2,4);
TASK_PP(16'hF3D3,4);
TASK_PP(16'hF3D4,4);
TASK_PP(16'hF3D5,4);
TASK_PP(16'hF3D6,4);
TASK_PP(16'hF3D7,4);
TASK_PP(16'hF3D8,4);
TASK_PP(16'hF3D9,4);
TASK_PP(16'hF3DA,4);
TASK_PP(16'hF3DB,4);
TASK_PP(16'hF3DC,4);
TASK_PP(16'hF3DD,4);
TASK_PP(16'hF3DE,4);
TASK_PP(16'hF3DF,4);
TASK_PP(16'hF3E0,4);
TASK_PP(16'hF3E1,4);
TASK_PP(16'hF3E2,4);
TASK_PP(16'hF3E3,4);
TASK_PP(16'hF3E4,4);
TASK_PP(16'hF3E5,4);
TASK_PP(16'hF3E6,4);
TASK_PP(16'hF3E7,4);
TASK_PP(16'hF3E8,4);
TASK_PP(16'hF3E9,4);
TASK_PP(16'hF3EA,4);
TASK_PP(16'hF3EB,4);
TASK_PP(16'hF3EC,4);
TASK_PP(16'hF3ED,4);
TASK_PP(16'hF3EE,4);
TASK_PP(16'hF3EF,4);
TASK_PP(16'hF3F0,4);
TASK_PP(16'hF3F1,4);
TASK_PP(16'hF3F2,4);
TASK_PP(16'hF3F3,4);
TASK_PP(16'hF3F4,4);
TASK_PP(16'hF3F5,4);
TASK_PP(16'hF3F6,4);
TASK_PP(16'hF3F7,4);
TASK_PP(16'hF3F8,4);
TASK_PP(16'hF3F9,4);
TASK_PP(16'hF3FA,4);
TASK_PP(16'hF3FB,4);
TASK_PP(16'hF3FC,4);
TASK_PP(16'hF3FD,4);
TASK_PP(16'hF3FE,4);
TASK_PP(16'hF3FF,4);
TASK_PP(16'hF400,4);
TASK_PP(16'hF401,4);
TASK_PP(16'hF402,4);
TASK_PP(16'hF403,4);
TASK_PP(16'hF404,4);
TASK_PP(16'hF405,4);
TASK_PP(16'hF406,4);
TASK_PP(16'hF407,4);
TASK_PP(16'hF408,4);
TASK_PP(16'hF409,4);
TASK_PP(16'hF40A,4);
TASK_PP(16'hF40B,4);
TASK_PP(16'hF40C,4);
TASK_PP(16'hF40D,4);
TASK_PP(16'hF40E,4);
TASK_PP(16'hF40F,4);
TASK_PP(16'hF410,4);
TASK_PP(16'hF411,4);
TASK_PP(16'hF412,4);
TASK_PP(16'hF413,4);
TASK_PP(16'hF414,4);
TASK_PP(16'hF415,4);
TASK_PP(16'hF416,4);
TASK_PP(16'hF417,4);
TASK_PP(16'hF418,4);
TASK_PP(16'hF419,4);
TASK_PP(16'hF41A,4);
TASK_PP(16'hF41B,4);
TASK_PP(16'hF41C,4);
TASK_PP(16'hF41D,4);
TASK_PP(16'hF41E,4);
TASK_PP(16'hF41F,4);
TASK_PP(16'hF420,4);
TASK_PP(16'hF421,4);
TASK_PP(16'hF422,4);
TASK_PP(16'hF423,4);
TASK_PP(16'hF424,4);
TASK_PP(16'hF425,4);
TASK_PP(16'hF426,4);
TASK_PP(16'hF427,4);
TASK_PP(16'hF428,4);
TASK_PP(16'hF429,4);
TASK_PP(16'hF42A,4);
TASK_PP(16'hF42B,4);
TASK_PP(16'hF42C,4);
TASK_PP(16'hF42D,4);
TASK_PP(16'hF42E,4);
TASK_PP(16'hF42F,4);
TASK_PP(16'hF430,4);
TASK_PP(16'hF431,4);
TASK_PP(16'hF432,4);
TASK_PP(16'hF433,4);
TASK_PP(16'hF434,4);
TASK_PP(16'hF435,4);
TASK_PP(16'hF436,4);
TASK_PP(16'hF437,4);
TASK_PP(16'hF438,4);
TASK_PP(16'hF439,4);
TASK_PP(16'hF43A,4);
TASK_PP(16'hF43B,4);
TASK_PP(16'hF43C,4);
TASK_PP(16'hF43D,4);
TASK_PP(16'hF43E,4);
TASK_PP(16'hF43F,4);
TASK_PP(16'hF440,4);
TASK_PP(16'hF441,4);
TASK_PP(16'hF442,4);
TASK_PP(16'hF443,4);
TASK_PP(16'hF444,4);
TASK_PP(16'hF445,4);
TASK_PP(16'hF446,4);
TASK_PP(16'hF447,4);
TASK_PP(16'hF448,4);
TASK_PP(16'hF449,4);
TASK_PP(16'hF44A,4);
TASK_PP(16'hF44B,4);
TASK_PP(16'hF44C,4);
TASK_PP(16'hF44D,4);
TASK_PP(16'hF44E,4);
TASK_PP(16'hF44F,4);
TASK_PP(16'hF450,4);
TASK_PP(16'hF451,4);
TASK_PP(16'hF452,4);
TASK_PP(16'hF453,4);
TASK_PP(16'hF454,4);
TASK_PP(16'hF455,4);
TASK_PP(16'hF456,4);
TASK_PP(16'hF457,4);
TASK_PP(16'hF458,4);
TASK_PP(16'hF459,4);
TASK_PP(16'hF45A,4);
TASK_PP(16'hF45B,4);
TASK_PP(16'hF45C,4);
TASK_PP(16'hF45D,4);
TASK_PP(16'hF45E,4);
TASK_PP(16'hF45F,4);
TASK_PP(16'hF460,4);
TASK_PP(16'hF461,4);
TASK_PP(16'hF462,4);
TASK_PP(16'hF463,4);
TASK_PP(16'hF464,4);
TASK_PP(16'hF465,4);
TASK_PP(16'hF466,4);
TASK_PP(16'hF467,4);
TASK_PP(16'hF468,4);
TASK_PP(16'hF469,4);
TASK_PP(16'hF46A,4);
TASK_PP(16'hF46B,4);
TASK_PP(16'hF46C,4);
TASK_PP(16'hF46D,4);
TASK_PP(16'hF46E,4);
TASK_PP(16'hF46F,4);
TASK_PP(16'hF470,4);
TASK_PP(16'hF471,4);
TASK_PP(16'hF472,4);
TASK_PP(16'hF473,4);
TASK_PP(16'hF474,4);
TASK_PP(16'hF475,4);
TASK_PP(16'hF476,4);
TASK_PP(16'hF477,4);
TASK_PP(16'hF478,4);
TASK_PP(16'hF479,4);
TASK_PP(16'hF47A,4);
TASK_PP(16'hF47B,4);
TASK_PP(16'hF47C,4);
TASK_PP(16'hF47D,4);
TASK_PP(16'hF47E,4);
TASK_PP(16'hF47F,4);
TASK_PP(16'hF480,4);
TASK_PP(16'hF481,4);
TASK_PP(16'hF482,4);
TASK_PP(16'hF483,4);
TASK_PP(16'hF484,4);
TASK_PP(16'hF485,4);
TASK_PP(16'hF486,4);
TASK_PP(16'hF487,4);
TASK_PP(16'hF488,4);
TASK_PP(16'hF489,4);
TASK_PP(16'hF48A,4);
TASK_PP(16'hF48B,4);
TASK_PP(16'hF48C,4);
TASK_PP(16'hF48D,4);
TASK_PP(16'hF48E,4);
TASK_PP(16'hF48F,4);
TASK_PP(16'hF490,4);
TASK_PP(16'hF491,4);
TASK_PP(16'hF492,4);
TASK_PP(16'hF493,4);
TASK_PP(16'hF494,4);
TASK_PP(16'hF495,4);
TASK_PP(16'hF496,4);
TASK_PP(16'hF497,4);
TASK_PP(16'hF498,4);
TASK_PP(16'hF499,4);
TASK_PP(16'hF49A,4);
TASK_PP(16'hF49B,4);
TASK_PP(16'hF49C,4);
TASK_PP(16'hF49D,4);
TASK_PP(16'hF49E,4);
TASK_PP(16'hF49F,4);
TASK_PP(16'hF4A0,4);
TASK_PP(16'hF4A1,4);
TASK_PP(16'hF4A2,4);
TASK_PP(16'hF4A3,4);
TASK_PP(16'hF4A4,4);
TASK_PP(16'hF4A5,4);
TASK_PP(16'hF4A6,4);
TASK_PP(16'hF4A7,4);
TASK_PP(16'hF4A8,4);
TASK_PP(16'hF4A9,4);
TASK_PP(16'hF4AA,4);
TASK_PP(16'hF4AB,4);
TASK_PP(16'hF4AC,4);
TASK_PP(16'hF4AD,4);
TASK_PP(16'hF4AE,4);
TASK_PP(16'hF4AF,4);
TASK_PP(16'hF4B0,4);
TASK_PP(16'hF4B1,4);
TASK_PP(16'hF4B2,4);
TASK_PP(16'hF4B3,4);
TASK_PP(16'hF4B4,4);
TASK_PP(16'hF4B5,4);
TASK_PP(16'hF4B6,4);
TASK_PP(16'hF4B7,4);
TASK_PP(16'hF4B8,4);
TASK_PP(16'hF4B9,4);
TASK_PP(16'hF4BA,4);
TASK_PP(16'hF4BB,4);
TASK_PP(16'hF4BC,4);
TASK_PP(16'hF4BD,4);
TASK_PP(16'hF4BE,4);
TASK_PP(16'hF4BF,4);
TASK_PP(16'hF4C0,4);
TASK_PP(16'hF4C1,4);
TASK_PP(16'hF4C2,4);
TASK_PP(16'hF4C3,4);
TASK_PP(16'hF4C4,4);
TASK_PP(16'hF4C5,4);
TASK_PP(16'hF4C6,4);
TASK_PP(16'hF4C7,4);
TASK_PP(16'hF4C8,4);
TASK_PP(16'hF4C9,4);
TASK_PP(16'hF4CA,4);
TASK_PP(16'hF4CB,4);
TASK_PP(16'hF4CC,4);
TASK_PP(16'hF4CD,4);
TASK_PP(16'hF4CE,4);
TASK_PP(16'hF4CF,4);
TASK_PP(16'hF4D0,4);
TASK_PP(16'hF4D1,4);
TASK_PP(16'hF4D2,4);
TASK_PP(16'hF4D3,4);
TASK_PP(16'hF4D4,4);
TASK_PP(16'hF4D5,4);
TASK_PP(16'hF4D6,4);
TASK_PP(16'hF4D7,4);
TASK_PP(16'hF4D8,4);
TASK_PP(16'hF4D9,4);
TASK_PP(16'hF4DA,4);
TASK_PP(16'hF4DB,4);
TASK_PP(16'hF4DC,4);
TASK_PP(16'hF4DD,4);
TASK_PP(16'hF4DE,4);
TASK_PP(16'hF4DF,4);
TASK_PP(16'hF4E0,4);
TASK_PP(16'hF4E1,4);
TASK_PP(16'hF4E2,4);
TASK_PP(16'hF4E3,4);
TASK_PP(16'hF4E4,4);
TASK_PP(16'hF4E5,4);
TASK_PP(16'hF4E6,4);
TASK_PP(16'hF4E7,4);
TASK_PP(16'hF4E8,4);
TASK_PP(16'hF4E9,4);
TASK_PP(16'hF4EA,4);
TASK_PP(16'hF4EB,4);
TASK_PP(16'hF4EC,4);
TASK_PP(16'hF4ED,4);
TASK_PP(16'hF4EE,4);
TASK_PP(16'hF4EF,4);
TASK_PP(16'hF4F0,4);
TASK_PP(16'hF4F1,4);
TASK_PP(16'hF4F2,4);
TASK_PP(16'hF4F3,4);
TASK_PP(16'hF4F4,4);
TASK_PP(16'hF4F5,4);
TASK_PP(16'hF4F6,4);
TASK_PP(16'hF4F7,4);
TASK_PP(16'hF4F8,4);
TASK_PP(16'hF4F9,4);
TASK_PP(16'hF4FA,4);
TASK_PP(16'hF4FB,4);
TASK_PP(16'hF4FC,4);
TASK_PP(16'hF4FD,4);
TASK_PP(16'hF4FE,4);
TASK_PP(16'hF4FF,4);
TASK_PP(16'hF500,4);
TASK_PP(16'hF501,4);
TASK_PP(16'hF502,4);
TASK_PP(16'hF503,4);
TASK_PP(16'hF504,4);
TASK_PP(16'hF505,4);
TASK_PP(16'hF506,4);
TASK_PP(16'hF507,4);
TASK_PP(16'hF508,4);
TASK_PP(16'hF509,4);
TASK_PP(16'hF50A,4);
TASK_PP(16'hF50B,4);
TASK_PP(16'hF50C,4);
TASK_PP(16'hF50D,4);
TASK_PP(16'hF50E,4);
TASK_PP(16'hF50F,4);
TASK_PP(16'hF510,4);
TASK_PP(16'hF511,4);
TASK_PP(16'hF512,4);
TASK_PP(16'hF513,4);
TASK_PP(16'hF514,4);
TASK_PP(16'hF515,4);
TASK_PP(16'hF516,4);
TASK_PP(16'hF517,4);
TASK_PP(16'hF518,4);
TASK_PP(16'hF519,4);
TASK_PP(16'hF51A,4);
TASK_PP(16'hF51B,4);
TASK_PP(16'hF51C,4);
TASK_PP(16'hF51D,4);
TASK_PP(16'hF51E,4);
TASK_PP(16'hF51F,4);
TASK_PP(16'hF520,4);
TASK_PP(16'hF521,4);
TASK_PP(16'hF522,4);
TASK_PP(16'hF523,4);
TASK_PP(16'hF524,4);
TASK_PP(16'hF525,4);
TASK_PP(16'hF526,4);
TASK_PP(16'hF527,4);
TASK_PP(16'hF528,4);
TASK_PP(16'hF529,4);
TASK_PP(16'hF52A,4);
TASK_PP(16'hF52B,4);
TASK_PP(16'hF52C,4);
TASK_PP(16'hF52D,4);
TASK_PP(16'hF52E,4);
TASK_PP(16'hF52F,4);
TASK_PP(16'hF530,4);
TASK_PP(16'hF531,4);
TASK_PP(16'hF532,4);
TASK_PP(16'hF533,4);
TASK_PP(16'hF534,4);
TASK_PP(16'hF535,4);
TASK_PP(16'hF536,4);
TASK_PP(16'hF537,4);
TASK_PP(16'hF538,4);
TASK_PP(16'hF539,4);
TASK_PP(16'hF53A,4);
TASK_PP(16'hF53B,4);
TASK_PP(16'hF53C,4);
TASK_PP(16'hF53D,4);
TASK_PP(16'hF53E,4);
TASK_PP(16'hF53F,4);
TASK_PP(16'hF540,4);
TASK_PP(16'hF541,4);
TASK_PP(16'hF542,4);
TASK_PP(16'hF543,4);
TASK_PP(16'hF544,4);
TASK_PP(16'hF545,4);
TASK_PP(16'hF546,4);
TASK_PP(16'hF547,4);
TASK_PP(16'hF548,4);
TASK_PP(16'hF549,4);
TASK_PP(16'hF54A,4);
TASK_PP(16'hF54B,4);
TASK_PP(16'hF54C,4);
TASK_PP(16'hF54D,4);
TASK_PP(16'hF54E,4);
TASK_PP(16'hF54F,4);
TASK_PP(16'hF550,4);
TASK_PP(16'hF551,4);
TASK_PP(16'hF552,4);
TASK_PP(16'hF553,4);
TASK_PP(16'hF554,4);
TASK_PP(16'hF555,4);
TASK_PP(16'hF556,4);
TASK_PP(16'hF557,4);
TASK_PP(16'hF558,4);
TASK_PP(16'hF559,4);
TASK_PP(16'hF55A,4);
TASK_PP(16'hF55B,4);
TASK_PP(16'hF55C,4);
TASK_PP(16'hF55D,4);
TASK_PP(16'hF55E,4);
TASK_PP(16'hF55F,4);
TASK_PP(16'hF560,4);
TASK_PP(16'hF561,4);
TASK_PP(16'hF562,4);
TASK_PP(16'hF563,4);
TASK_PP(16'hF564,4);
TASK_PP(16'hF565,4);
TASK_PP(16'hF566,4);
TASK_PP(16'hF567,4);
TASK_PP(16'hF568,4);
TASK_PP(16'hF569,4);
TASK_PP(16'hF56A,4);
TASK_PP(16'hF56B,4);
TASK_PP(16'hF56C,4);
TASK_PP(16'hF56D,4);
TASK_PP(16'hF56E,4);
TASK_PP(16'hF56F,4);
TASK_PP(16'hF570,4);
TASK_PP(16'hF571,4);
TASK_PP(16'hF572,4);
TASK_PP(16'hF573,4);
TASK_PP(16'hF574,4);
TASK_PP(16'hF575,4);
TASK_PP(16'hF576,4);
TASK_PP(16'hF577,4);
TASK_PP(16'hF578,4);
TASK_PP(16'hF579,4);
TASK_PP(16'hF57A,4);
TASK_PP(16'hF57B,4);
TASK_PP(16'hF57C,4);
TASK_PP(16'hF57D,4);
TASK_PP(16'hF57E,4);
TASK_PP(16'hF57F,4);
TASK_PP(16'hF580,4);
TASK_PP(16'hF581,4);
TASK_PP(16'hF582,4);
TASK_PP(16'hF583,4);
TASK_PP(16'hF584,4);
TASK_PP(16'hF585,4);
TASK_PP(16'hF586,4);
TASK_PP(16'hF587,4);
TASK_PP(16'hF588,4);
TASK_PP(16'hF589,4);
TASK_PP(16'hF58A,4);
TASK_PP(16'hF58B,4);
TASK_PP(16'hF58C,4);
TASK_PP(16'hF58D,4);
TASK_PP(16'hF58E,4);
TASK_PP(16'hF58F,4);
TASK_PP(16'hF590,4);
TASK_PP(16'hF591,4);
TASK_PP(16'hF592,4);
TASK_PP(16'hF593,4);
TASK_PP(16'hF594,4);
TASK_PP(16'hF595,4);
TASK_PP(16'hF596,4);
TASK_PP(16'hF597,4);
TASK_PP(16'hF598,4);
TASK_PP(16'hF599,4);
TASK_PP(16'hF59A,4);
TASK_PP(16'hF59B,4);
TASK_PP(16'hF59C,4);
TASK_PP(16'hF59D,4);
TASK_PP(16'hF59E,4);
TASK_PP(16'hF59F,4);
TASK_PP(16'hF5A0,4);
TASK_PP(16'hF5A1,4);
TASK_PP(16'hF5A2,4);
TASK_PP(16'hF5A3,4);
TASK_PP(16'hF5A4,4);
TASK_PP(16'hF5A5,4);
TASK_PP(16'hF5A6,4);
TASK_PP(16'hF5A7,4);
TASK_PP(16'hF5A8,4);
TASK_PP(16'hF5A9,4);
TASK_PP(16'hF5AA,4);
TASK_PP(16'hF5AB,4);
TASK_PP(16'hF5AC,4);
TASK_PP(16'hF5AD,4);
TASK_PP(16'hF5AE,4);
TASK_PP(16'hF5AF,4);
TASK_PP(16'hF5B0,4);
TASK_PP(16'hF5B1,4);
TASK_PP(16'hF5B2,4);
TASK_PP(16'hF5B3,4);
TASK_PP(16'hF5B4,4);
TASK_PP(16'hF5B5,4);
TASK_PP(16'hF5B6,4);
TASK_PP(16'hF5B7,4);
TASK_PP(16'hF5B8,4);
TASK_PP(16'hF5B9,4);
TASK_PP(16'hF5BA,4);
TASK_PP(16'hF5BB,4);
TASK_PP(16'hF5BC,4);
TASK_PP(16'hF5BD,4);
TASK_PP(16'hF5BE,4);
TASK_PP(16'hF5BF,4);
TASK_PP(16'hF5C0,4);
TASK_PP(16'hF5C1,4);
TASK_PP(16'hF5C2,4);
TASK_PP(16'hF5C3,4);
TASK_PP(16'hF5C4,4);
TASK_PP(16'hF5C5,4);
TASK_PP(16'hF5C6,4);
TASK_PP(16'hF5C7,4);
TASK_PP(16'hF5C8,4);
TASK_PP(16'hF5C9,4);
TASK_PP(16'hF5CA,4);
TASK_PP(16'hF5CB,4);
TASK_PP(16'hF5CC,4);
TASK_PP(16'hF5CD,4);
TASK_PP(16'hF5CE,4);
TASK_PP(16'hF5CF,4);
TASK_PP(16'hF5D0,4);
TASK_PP(16'hF5D1,4);
TASK_PP(16'hF5D2,4);
TASK_PP(16'hF5D3,4);
TASK_PP(16'hF5D4,4);
TASK_PP(16'hF5D5,4);
TASK_PP(16'hF5D6,4);
TASK_PP(16'hF5D7,4);
TASK_PP(16'hF5D8,4);
TASK_PP(16'hF5D9,4);
TASK_PP(16'hF5DA,4);
TASK_PP(16'hF5DB,4);
TASK_PP(16'hF5DC,4);
TASK_PP(16'hF5DD,4);
TASK_PP(16'hF5DE,4);
TASK_PP(16'hF5DF,4);
TASK_PP(16'hF5E0,4);
TASK_PP(16'hF5E1,4);
TASK_PP(16'hF5E2,4);
TASK_PP(16'hF5E3,4);
TASK_PP(16'hF5E4,4);
TASK_PP(16'hF5E5,4);
TASK_PP(16'hF5E6,4);
TASK_PP(16'hF5E7,4);
TASK_PP(16'hF5E8,4);
TASK_PP(16'hF5E9,4);
TASK_PP(16'hF5EA,4);
TASK_PP(16'hF5EB,4);
TASK_PP(16'hF5EC,4);
TASK_PP(16'hF5ED,4);
TASK_PP(16'hF5EE,4);
TASK_PP(16'hF5EF,4);
TASK_PP(16'hF5F0,4);
TASK_PP(16'hF5F1,4);
TASK_PP(16'hF5F2,4);
TASK_PP(16'hF5F3,4);
TASK_PP(16'hF5F4,4);
TASK_PP(16'hF5F5,4);
TASK_PP(16'hF5F6,4);
TASK_PP(16'hF5F7,4);
TASK_PP(16'hF5F8,4);
TASK_PP(16'hF5F9,4);
TASK_PP(16'hF5FA,4);
TASK_PP(16'hF5FB,4);
TASK_PP(16'hF5FC,4);
TASK_PP(16'hF5FD,4);
TASK_PP(16'hF5FE,4);
TASK_PP(16'hF5FF,4);
TASK_PP(16'hF600,4);
TASK_PP(16'hF601,4);
TASK_PP(16'hF602,4);
TASK_PP(16'hF603,4);
TASK_PP(16'hF604,4);
TASK_PP(16'hF605,4);
TASK_PP(16'hF606,4);
TASK_PP(16'hF607,4);
TASK_PP(16'hF608,4);
TASK_PP(16'hF609,4);
TASK_PP(16'hF60A,4);
TASK_PP(16'hF60B,4);
TASK_PP(16'hF60C,4);
TASK_PP(16'hF60D,4);
TASK_PP(16'hF60E,4);
TASK_PP(16'hF60F,4);
TASK_PP(16'hF610,4);
TASK_PP(16'hF611,4);
TASK_PP(16'hF612,4);
TASK_PP(16'hF613,4);
TASK_PP(16'hF614,4);
TASK_PP(16'hF615,4);
TASK_PP(16'hF616,4);
TASK_PP(16'hF617,4);
TASK_PP(16'hF618,4);
TASK_PP(16'hF619,4);
TASK_PP(16'hF61A,4);
TASK_PP(16'hF61B,4);
TASK_PP(16'hF61C,4);
TASK_PP(16'hF61D,4);
TASK_PP(16'hF61E,4);
TASK_PP(16'hF61F,4);
TASK_PP(16'hF620,4);
TASK_PP(16'hF621,4);
TASK_PP(16'hF622,4);
TASK_PP(16'hF623,4);
TASK_PP(16'hF624,4);
TASK_PP(16'hF625,4);
TASK_PP(16'hF626,4);
TASK_PP(16'hF627,4);
TASK_PP(16'hF628,4);
TASK_PP(16'hF629,4);
TASK_PP(16'hF62A,4);
TASK_PP(16'hF62B,4);
TASK_PP(16'hF62C,4);
TASK_PP(16'hF62D,4);
TASK_PP(16'hF62E,4);
TASK_PP(16'hF62F,4);
TASK_PP(16'hF630,4);
TASK_PP(16'hF631,4);
TASK_PP(16'hF632,4);
TASK_PP(16'hF633,4);
TASK_PP(16'hF634,4);
TASK_PP(16'hF635,4);
TASK_PP(16'hF636,4);
TASK_PP(16'hF637,4);
TASK_PP(16'hF638,4);
TASK_PP(16'hF639,4);
TASK_PP(16'hF63A,4);
TASK_PP(16'hF63B,4);
TASK_PP(16'hF63C,4);
TASK_PP(16'hF63D,4);
TASK_PP(16'hF63E,4);
TASK_PP(16'hF63F,4);
TASK_PP(16'hF640,4);
TASK_PP(16'hF641,4);
TASK_PP(16'hF642,4);
TASK_PP(16'hF643,4);
TASK_PP(16'hF644,4);
TASK_PP(16'hF645,4);
TASK_PP(16'hF646,4);
TASK_PP(16'hF647,4);
TASK_PP(16'hF648,4);
TASK_PP(16'hF649,4);
TASK_PP(16'hF64A,4);
TASK_PP(16'hF64B,4);
TASK_PP(16'hF64C,4);
TASK_PP(16'hF64D,4);
TASK_PP(16'hF64E,4);
TASK_PP(16'hF64F,4);
TASK_PP(16'hF650,4);
TASK_PP(16'hF651,4);
TASK_PP(16'hF652,4);
TASK_PP(16'hF653,4);
TASK_PP(16'hF654,4);
TASK_PP(16'hF655,4);
TASK_PP(16'hF656,4);
TASK_PP(16'hF657,4);
TASK_PP(16'hF658,4);
TASK_PP(16'hF659,4);
TASK_PP(16'hF65A,4);
TASK_PP(16'hF65B,4);
TASK_PP(16'hF65C,4);
TASK_PP(16'hF65D,4);
TASK_PP(16'hF65E,4);
TASK_PP(16'hF65F,4);
TASK_PP(16'hF660,4);
TASK_PP(16'hF661,4);
TASK_PP(16'hF662,4);
TASK_PP(16'hF663,4);
TASK_PP(16'hF664,4);
TASK_PP(16'hF665,4);
TASK_PP(16'hF666,4);
TASK_PP(16'hF667,4);
TASK_PP(16'hF668,4);
TASK_PP(16'hF669,4);
TASK_PP(16'hF66A,4);
TASK_PP(16'hF66B,4);
TASK_PP(16'hF66C,4);
TASK_PP(16'hF66D,4);
TASK_PP(16'hF66E,4);
TASK_PP(16'hF66F,4);
TASK_PP(16'hF670,4);
TASK_PP(16'hF671,4);
TASK_PP(16'hF672,4);
TASK_PP(16'hF673,4);
TASK_PP(16'hF674,4);
TASK_PP(16'hF675,4);
TASK_PP(16'hF676,4);
TASK_PP(16'hF677,4);
TASK_PP(16'hF678,4);
TASK_PP(16'hF679,4);
TASK_PP(16'hF67A,4);
TASK_PP(16'hF67B,4);
TASK_PP(16'hF67C,4);
TASK_PP(16'hF67D,4);
TASK_PP(16'hF67E,4);
TASK_PP(16'hF67F,4);
TASK_PP(16'hF680,4);
TASK_PP(16'hF681,4);
TASK_PP(16'hF682,4);
TASK_PP(16'hF683,4);
TASK_PP(16'hF684,4);
TASK_PP(16'hF685,4);
TASK_PP(16'hF686,4);
TASK_PP(16'hF687,4);
TASK_PP(16'hF688,4);
TASK_PP(16'hF689,4);
TASK_PP(16'hF68A,4);
TASK_PP(16'hF68B,4);
TASK_PP(16'hF68C,4);
TASK_PP(16'hF68D,4);
TASK_PP(16'hF68E,4);
TASK_PP(16'hF68F,4);
TASK_PP(16'hF690,4);
TASK_PP(16'hF691,4);
TASK_PP(16'hF692,4);
TASK_PP(16'hF693,4);
TASK_PP(16'hF694,4);
TASK_PP(16'hF695,4);
TASK_PP(16'hF696,4);
TASK_PP(16'hF697,4);
TASK_PP(16'hF698,4);
TASK_PP(16'hF699,4);
TASK_PP(16'hF69A,4);
TASK_PP(16'hF69B,4);
TASK_PP(16'hF69C,4);
TASK_PP(16'hF69D,4);
TASK_PP(16'hF69E,4);
TASK_PP(16'hF69F,4);
TASK_PP(16'hF6A0,4);
TASK_PP(16'hF6A1,4);
TASK_PP(16'hF6A2,4);
TASK_PP(16'hF6A3,4);
TASK_PP(16'hF6A4,4);
TASK_PP(16'hF6A5,4);
TASK_PP(16'hF6A6,4);
TASK_PP(16'hF6A7,4);
TASK_PP(16'hF6A8,4);
TASK_PP(16'hF6A9,4);
TASK_PP(16'hF6AA,4);
TASK_PP(16'hF6AB,4);
TASK_PP(16'hF6AC,4);
TASK_PP(16'hF6AD,4);
TASK_PP(16'hF6AE,4);
TASK_PP(16'hF6AF,4);
TASK_PP(16'hF6B0,4);
TASK_PP(16'hF6B1,4);
TASK_PP(16'hF6B2,4);
TASK_PP(16'hF6B3,4);
TASK_PP(16'hF6B4,4);
TASK_PP(16'hF6B5,4);
TASK_PP(16'hF6B6,4);
TASK_PP(16'hF6B7,4);
TASK_PP(16'hF6B8,4);
TASK_PP(16'hF6B9,4);
TASK_PP(16'hF6BA,4);
TASK_PP(16'hF6BB,4);
TASK_PP(16'hF6BC,4);
TASK_PP(16'hF6BD,4);
TASK_PP(16'hF6BE,4);
TASK_PP(16'hF6BF,4);
TASK_PP(16'hF6C0,4);
TASK_PP(16'hF6C1,4);
TASK_PP(16'hF6C2,4);
TASK_PP(16'hF6C3,4);
TASK_PP(16'hF6C4,4);
TASK_PP(16'hF6C5,4);
TASK_PP(16'hF6C6,4);
TASK_PP(16'hF6C7,4);
TASK_PP(16'hF6C8,4);
TASK_PP(16'hF6C9,4);
TASK_PP(16'hF6CA,4);
TASK_PP(16'hF6CB,4);
TASK_PP(16'hF6CC,4);
TASK_PP(16'hF6CD,4);
TASK_PP(16'hF6CE,4);
TASK_PP(16'hF6CF,4);
TASK_PP(16'hF6D0,4);
TASK_PP(16'hF6D1,4);
TASK_PP(16'hF6D2,4);
TASK_PP(16'hF6D3,4);
TASK_PP(16'hF6D4,4);
TASK_PP(16'hF6D5,4);
TASK_PP(16'hF6D6,4);
TASK_PP(16'hF6D7,4);
TASK_PP(16'hF6D8,4);
TASK_PP(16'hF6D9,4);
TASK_PP(16'hF6DA,4);
TASK_PP(16'hF6DB,4);
TASK_PP(16'hF6DC,4);
TASK_PP(16'hF6DD,4);
TASK_PP(16'hF6DE,4);
TASK_PP(16'hF6DF,4);
TASK_PP(16'hF6E0,4);
TASK_PP(16'hF6E1,4);
TASK_PP(16'hF6E2,4);
TASK_PP(16'hF6E3,4);
TASK_PP(16'hF6E4,4);
TASK_PP(16'hF6E5,4);
TASK_PP(16'hF6E6,4);
TASK_PP(16'hF6E7,4);
TASK_PP(16'hF6E8,4);
TASK_PP(16'hF6E9,4);
TASK_PP(16'hF6EA,4);
TASK_PP(16'hF6EB,4);
TASK_PP(16'hF6EC,4);
TASK_PP(16'hF6ED,4);
TASK_PP(16'hF6EE,4);
TASK_PP(16'hF6EF,4);
TASK_PP(16'hF6F0,4);
TASK_PP(16'hF6F1,4);
TASK_PP(16'hF6F2,4);
TASK_PP(16'hF6F3,4);
TASK_PP(16'hF6F4,4);
TASK_PP(16'hF6F5,4);
TASK_PP(16'hF6F6,4);
TASK_PP(16'hF6F7,4);
TASK_PP(16'hF6F8,4);
TASK_PP(16'hF6F9,4);
TASK_PP(16'hF6FA,4);
TASK_PP(16'hF6FB,4);
TASK_PP(16'hF6FC,4);
TASK_PP(16'hF6FD,4);
TASK_PP(16'hF6FE,4);
TASK_PP(16'hF6FF,4);
TASK_PP(16'hF700,4);
TASK_PP(16'hF701,4);
TASK_PP(16'hF702,4);
TASK_PP(16'hF703,4);
TASK_PP(16'hF704,4);
TASK_PP(16'hF705,4);
TASK_PP(16'hF706,4);
TASK_PP(16'hF707,4);
TASK_PP(16'hF708,4);
TASK_PP(16'hF709,4);
TASK_PP(16'hF70A,4);
TASK_PP(16'hF70B,4);
TASK_PP(16'hF70C,4);
TASK_PP(16'hF70D,4);
TASK_PP(16'hF70E,4);
TASK_PP(16'hF70F,4);
TASK_PP(16'hF710,4);
TASK_PP(16'hF711,4);
TASK_PP(16'hF712,4);
TASK_PP(16'hF713,4);
TASK_PP(16'hF714,4);
TASK_PP(16'hF715,4);
TASK_PP(16'hF716,4);
TASK_PP(16'hF717,4);
TASK_PP(16'hF718,4);
TASK_PP(16'hF719,4);
TASK_PP(16'hF71A,4);
TASK_PP(16'hF71B,4);
TASK_PP(16'hF71C,4);
TASK_PP(16'hF71D,4);
TASK_PP(16'hF71E,4);
TASK_PP(16'hF71F,4);
TASK_PP(16'hF720,4);
TASK_PP(16'hF721,4);
TASK_PP(16'hF722,4);
TASK_PP(16'hF723,4);
TASK_PP(16'hF724,4);
TASK_PP(16'hF725,4);
TASK_PP(16'hF726,4);
TASK_PP(16'hF727,4);
TASK_PP(16'hF728,4);
TASK_PP(16'hF729,4);
TASK_PP(16'hF72A,4);
TASK_PP(16'hF72B,4);
TASK_PP(16'hF72C,4);
TASK_PP(16'hF72D,4);
TASK_PP(16'hF72E,4);
TASK_PP(16'hF72F,4);
TASK_PP(16'hF730,4);
TASK_PP(16'hF731,4);
TASK_PP(16'hF732,4);
TASK_PP(16'hF733,4);
TASK_PP(16'hF734,4);
TASK_PP(16'hF735,4);
TASK_PP(16'hF736,4);
TASK_PP(16'hF737,4);
TASK_PP(16'hF738,4);
TASK_PP(16'hF739,4);
TASK_PP(16'hF73A,4);
TASK_PP(16'hF73B,4);
TASK_PP(16'hF73C,4);
TASK_PP(16'hF73D,4);
TASK_PP(16'hF73E,4);
TASK_PP(16'hF73F,4);
TASK_PP(16'hF740,4);
TASK_PP(16'hF741,4);
TASK_PP(16'hF742,4);
TASK_PP(16'hF743,4);
TASK_PP(16'hF744,4);
TASK_PP(16'hF745,4);
TASK_PP(16'hF746,4);
TASK_PP(16'hF747,4);
TASK_PP(16'hF748,4);
TASK_PP(16'hF749,4);
TASK_PP(16'hF74A,4);
TASK_PP(16'hF74B,4);
TASK_PP(16'hF74C,4);
TASK_PP(16'hF74D,4);
TASK_PP(16'hF74E,4);
TASK_PP(16'hF74F,4);
TASK_PP(16'hF750,4);
TASK_PP(16'hF751,4);
TASK_PP(16'hF752,4);
TASK_PP(16'hF753,4);
TASK_PP(16'hF754,4);
TASK_PP(16'hF755,4);
TASK_PP(16'hF756,4);
TASK_PP(16'hF757,4);
TASK_PP(16'hF758,4);
TASK_PP(16'hF759,4);
TASK_PP(16'hF75A,4);
TASK_PP(16'hF75B,4);
TASK_PP(16'hF75C,4);
TASK_PP(16'hF75D,4);
TASK_PP(16'hF75E,4);
TASK_PP(16'hF75F,4);
TASK_PP(16'hF760,4);
TASK_PP(16'hF761,4);
TASK_PP(16'hF762,4);
TASK_PP(16'hF763,4);
TASK_PP(16'hF764,4);
TASK_PP(16'hF765,4);
TASK_PP(16'hF766,4);
TASK_PP(16'hF767,4);
TASK_PP(16'hF768,4);
TASK_PP(16'hF769,4);
TASK_PP(16'hF76A,4);
TASK_PP(16'hF76B,4);
TASK_PP(16'hF76C,4);
TASK_PP(16'hF76D,4);
TASK_PP(16'hF76E,4);
TASK_PP(16'hF76F,4);
TASK_PP(16'hF770,4);
TASK_PP(16'hF771,4);
TASK_PP(16'hF772,4);
TASK_PP(16'hF773,4);
TASK_PP(16'hF774,4);
TASK_PP(16'hF775,4);
TASK_PP(16'hF776,4);
TASK_PP(16'hF777,4);
TASK_PP(16'hF778,4);
TASK_PP(16'hF779,4);
TASK_PP(16'hF77A,4);
TASK_PP(16'hF77B,4);
TASK_PP(16'hF77C,4);
TASK_PP(16'hF77D,4);
TASK_PP(16'hF77E,4);
TASK_PP(16'hF77F,4);
TASK_PP(16'hF780,4);
TASK_PP(16'hF781,4);
TASK_PP(16'hF782,4);
TASK_PP(16'hF783,4);
TASK_PP(16'hF784,4);
TASK_PP(16'hF785,4);
TASK_PP(16'hF786,4);
TASK_PP(16'hF787,4);
TASK_PP(16'hF788,4);
TASK_PP(16'hF789,4);
TASK_PP(16'hF78A,4);
TASK_PP(16'hF78B,4);
TASK_PP(16'hF78C,4);
TASK_PP(16'hF78D,4);
TASK_PP(16'hF78E,4);
TASK_PP(16'hF78F,4);
TASK_PP(16'hF790,4);
TASK_PP(16'hF791,4);
TASK_PP(16'hF792,4);
TASK_PP(16'hF793,4);
TASK_PP(16'hF794,4);
TASK_PP(16'hF795,4);
TASK_PP(16'hF796,4);
TASK_PP(16'hF797,4);
TASK_PP(16'hF798,4);
TASK_PP(16'hF799,4);
TASK_PP(16'hF79A,4);
TASK_PP(16'hF79B,4);
TASK_PP(16'hF79C,4);
TASK_PP(16'hF79D,4);
TASK_PP(16'hF79E,4);
TASK_PP(16'hF79F,4);
TASK_PP(16'hF7A0,4);
TASK_PP(16'hF7A1,4);
TASK_PP(16'hF7A2,4);
TASK_PP(16'hF7A3,4);
TASK_PP(16'hF7A4,4);
TASK_PP(16'hF7A5,4);
TASK_PP(16'hF7A6,4);
TASK_PP(16'hF7A7,4);
TASK_PP(16'hF7A8,4);
TASK_PP(16'hF7A9,4);
TASK_PP(16'hF7AA,4);
TASK_PP(16'hF7AB,4);
TASK_PP(16'hF7AC,4);
TASK_PP(16'hF7AD,4);
TASK_PP(16'hF7AE,4);
TASK_PP(16'hF7AF,4);
TASK_PP(16'hF7B0,4);
TASK_PP(16'hF7B1,4);
TASK_PP(16'hF7B2,4);
TASK_PP(16'hF7B3,4);
TASK_PP(16'hF7B4,4);
TASK_PP(16'hF7B5,4);
TASK_PP(16'hF7B6,4);
TASK_PP(16'hF7B7,4);
TASK_PP(16'hF7B8,4);
TASK_PP(16'hF7B9,4);
TASK_PP(16'hF7BA,4);
TASK_PP(16'hF7BB,4);
TASK_PP(16'hF7BC,4);
TASK_PP(16'hF7BD,4);
TASK_PP(16'hF7BE,4);
TASK_PP(16'hF7BF,4);
TASK_PP(16'hF7C0,4);
TASK_PP(16'hF7C1,4);
TASK_PP(16'hF7C2,4);
TASK_PP(16'hF7C3,4);
TASK_PP(16'hF7C4,4);
TASK_PP(16'hF7C5,4);
TASK_PP(16'hF7C6,4);
TASK_PP(16'hF7C7,4);
TASK_PP(16'hF7C8,4);
TASK_PP(16'hF7C9,4);
TASK_PP(16'hF7CA,4);
TASK_PP(16'hF7CB,4);
TASK_PP(16'hF7CC,4);
TASK_PP(16'hF7CD,4);
TASK_PP(16'hF7CE,4);
TASK_PP(16'hF7CF,4);
TASK_PP(16'hF7D0,4);
TASK_PP(16'hF7D1,4);
TASK_PP(16'hF7D2,4);
TASK_PP(16'hF7D3,4);
TASK_PP(16'hF7D4,4);
TASK_PP(16'hF7D5,4);
TASK_PP(16'hF7D6,4);
TASK_PP(16'hF7D7,4);
TASK_PP(16'hF7D8,4);
TASK_PP(16'hF7D9,4);
TASK_PP(16'hF7DA,4);
TASK_PP(16'hF7DB,4);
TASK_PP(16'hF7DC,4);
TASK_PP(16'hF7DD,4);
TASK_PP(16'hF7DE,4);
TASK_PP(16'hF7DF,4);
TASK_PP(16'hF7E0,4);
TASK_PP(16'hF7E1,4);
TASK_PP(16'hF7E2,4);
TASK_PP(16'hF7E3,4);
TASK_PP(16'hF7E4,4);
TASK_PP(16'hF7E5,4);
TASK_PP(16'hF7E6,4);
TASK_PP(16'hF7E7,4);
TASK_PP(16'hF7E8,4);
TASK_PP(16'hF7E9,4);
TASK_PP(16'hF7EA,4);
TASK_PP(16'hF7EB,4);
TASK_PP(16'hF7EC,4);
TASK_PP(16'hF7ED,4);
TASK_PP(16'hF7EE,4);
TASK_PP(16'hF7EF,4);
TASK_PP(16'hF7F0,4);
TASK_PP(16'hF7F1,4);
TASK_PP(16'hF7F2,4);
TASK_PP(16'hF7F3,4);
TASK_PP(16'hF7F4,4);
TASK_PP(16'hF7F5,4);
TASK_PP(16'hF7F6,4);
TASK_PP(16'hF7F7,4);
TASK_PP(16'hF7F8,4);
TASK_PP(16'hF7F9,4);
TASK_PP(16'hF7FA,4);
TASK_PP(16'hF7FB,4);
TASK_PP(16'hF7FC,4);
TASK_PP(16'hF7FD,4);
TASK_PP(16'hF7FE,4);
TASK_PP(16'hF7FF,4);
TASK_PP(16'hF800,4);
TASK_PP(16'hF801,4);
TASK_PP(16'hF802,4);
TASK_PP(16'hF803,4);
TASK_PP(16'hF804,4);
TASK_PP(16'hF805,4);
TASK_PP(16'hF806,4);
TASK_PP(16'hF807,4);
TASK_PP(16'hF808,4);
TASK_PP(16'hF809,4);
TASK_PP(16'hF80A,4);
TASK_PP(16'hF80B,4);
TASK_PP(16'hF80C,4);
TASK_PP(16'hF80D,4);
TASK_PP(16'hF80E,4);
TASK_PP(16'hF80F,4);
TASK_PP(16'hF810,4);
TASK_PP(16'hF811,4);
TASK_PP(16'hF812,4);
TASK_PP(16'hF813,4);
TASK_PP(16'hF814,4);
TASK_PP(16'hF815,4);
TASK_PP(16'hF816,4);
TASK_PP(16'hF817,4);
TASK_PP(16'hF818,4);
TASK_PP(16'hF819,4);
TASK_PP(16'hF81A,4);
TASK_PP(16'hF81B,4);
TASK_PP(16'hF81C,4);
TASK_PP(16'hF81D,4);
TASK_PP(16'hF81E,4);
TASK_PP(16'hF81F,4);
TASK_PP(16'hF820,4);
TASK_PP(16'hF821,4);
TASK_PP(16'hF822,4);
TASK_PP(16'hF823,4);
TASK_PP(16'hF824,4);
TASK_PP(16'hF825,4);
TASK_PP(16'hF826,4);
TASK_PP(16'hF827,4);
TASK_PP(16'hF828,4);
TASK_PP(16'hF829,4);
TASK_PP(16'hF82A,4);
TASK_PP(16'hF82B,4);
TASK_PP(16'hF82C,4);
TASK_PP(16'hF82D,4);
TASK_PP(16'hF82E,4);
TASK_PP(16'hF82F,4);
TASK_PP(16'hF830,4);
TASK_PP(16'hF831,4);
TASK_PP(16'hF832,4);
TASK_PP(16'hF833,4);
TASK_PP(16'hF834,4);
TASK_PP(16'hF835,4);
TASK_PP(16'hF836,4);
TASK_PP(16'hF837,4);
TASK_PP(16'hF838,4);
TASK_PP(16'hF839,4);
TASK_PP(16'hF83A,4);
TASK_PP(16'hF83B,4);
TASK_PP(16'hF83C,4);
TASK_PP(16'hF83D,4);
TASK_PP(16'hF83E,4);
TASK_PP(16'hF83F,4);
TASK_PP(16'hF840,4);
TASK_PP(16'hF841,4);
TASK_PP(16'hF842,4);
TASK_PP(16'hF843,4);
TASK_PP(16'hF844,4);
TASK_PP(16'hF845,4);
TASK_PP(16'hF846,4);
TASK_PP(16'hF847,4);
TASK_PP(16'hF848,4);
TASK_PP(16'hF849,4);
TASK_PP(16'hF84A,4);
TASK_PP(16'hF84B,4);
TASK_PP(16'hF84C,4);
TASK_PP(16'hF84D,4);
TASK_PP(16'hF84E,4);
TASK_PP(16'hF84F,4);
TASK_PP(16'hF850,4);
TASK_PP(16'hF851,4);
TASK_PP(16'hF852,4);
TASK_PP(16'hF853,4);
TASK_PP(16'hF854,4);
TASK_PP(16'hF855,4);
TASK_PP(16'hF856,4);
TASK_PP(16'hF857,4);
TASK_PP(16'hF858,4);
TASK_PP(16'hF859,4);
TASK_PP(16'hF85A,4);
TASK_PP(16'hF85B,4);
TASK_PP(16'hF85C,4);
TASK_PP(16'hF85D,4);
TASK_PP(16'hF85E,4);
TASK_PP(16'hF85F,4);
TASK_PP(16'hF860,4);
TASK_PP(16'hF861,4);
TASK_PP(16'hF862,4);
TASK_PP(16'hF863,4);
TASK_PP(16'hF864,4);
TASK_PP(16'hF865,4);
TASK_PP(16'hF866,4);
TASK_PP(16'hF867,4);
TASK_PP(16'hF868,4);
TASK_PP(16'hF869,4);
TASK_PP(16'hF86A,4);
TASK_PP(16'hF86B,4);
TASK_PP(16'hF86C,4);
TASK_PP(16'hF86D,4);
TASK_PP(16'hF86E,4);
TASK_PP(16'hF86F,4);
TASK_PP(16'hF870,4);
TASK_PP(16'hF871,4);
TASK_PP(16'hF872,4);
TASK_PP(16'hF873,4);
TASK_PP(16'hF874,4);
TASK_PP(16'hF875,4);
TASK_PP(16'hF876,4);
TASK_PP(16'hF877,4);
TASK_PP(16'hF878,4);
TASK_PP(16'hF879,4);
TASK_PP(16'hF87A,4);
TASK_PP(16'hF87B,4);
TASK_PP(16'hF87C,4);
TASK_PP(16'hF87D,4);
TASK_PP(16'hF87E,4);
TASK_PP(16'hF87F,4);
TASK_PP(16'hF880,4);
TASK_PP(16'hF881,4);
TASK_PP(16'hF882,4);
TASK_PP(16'hF883,4);
TASK_PP(16'hF884,4);
TASK_PP(16'hF885,4);
TASK_PP(16'hF886,4);
TASK_PP(16'hF887,4);
TASK_PP(16'hF888,4);
TASK_PP(16'hF889,4);
TASK_PP(16'hF88A,4);
TASK_PP(16'hF88B,4);
TASK_PP(16'hF88C,4);
TASK_PP(16'hF88D,4);
TASK_PP(16'hF88E,4);
TASK_PP(16'hF88F,4);
TASK_PP(16'hF890,4);
TASK_PP(16'hF891,4);
TASK_PP(16'hF892,4);
TASK_PP(16'hF893,4);
TASK_PP(16'hF894,4);
TASK_PP(16'hF895,4);
TASK_PP(16'hF896,4);
TASK_PP(16'hF897,4);
TASK_PP(16'hF898,4);
TASK_PP(16'hF899,4);
TASK_PP(16'hF89A,4);
TASK_PP(16'hF89B,4);
TASK_PP(16'hF89C,4);
TASK_PP(16'hF89D,4);
TASK_PP(16'hF89E,4);
TASK_PP(16'hF89F,4);
TASK_PP(16'hF8A0,4);
TASK_PP(16'hF8A1,4);
TASK_PP(16'hF8A2,4);
TASK_PP(16'hF8A3,4);
TASK_PP(16'hF8A4,4);
TASK_PP(16'hF8A5,4);
TASK_PP(16'hF8A6,4);
TASK_PP(16'hF8A7,4);
TASK_PP(16'hF8A8,4);
TASK_PP(16'hF8A9,4);
TASK_PP(16'hF8AA,4);
TASK_PP(16'hF8AB,4);
TASK_PP(16'hF8AC,4);
TASK_PP(16'hF8AD,4);
TASK_PP(16'hF8AE,4);
TASK_PP(16'hF8AF,4);
TASK_PP(16'hF8B0,4);
TASK_PP(16'hF8B1,4);
TASK_PP(16'hF8B2,4);
TASK_PP(16'hF8B3,4);
TASK_PP(16'hF8B4,4);
TASK_PP(16'hF8B5,4);
TASK_PP(16'hF8B6,4);
TASK_PP(16'hF8B7,4);
TASK_PP(16'hF8B8,4);
TASK_PP(16'hF8B9,4);
TASK_PP(16'hF8BA,4);
TASK_PP(16'hF8BB,4);
TASK_PP(16'hF8BC,4);
TASK_PP(16'hF8BD,4);
TASK_PP(16'hF8BE,4);
TASK_PP(16'hF8BF,4);
TASK_PP(16'hF8C0,4);
TASK_PP(16'hF8C1,4);
TASK_PP(16'hF8C2,4);
TASK_PP(16'hF8C3,4);
TASK_PP(16'hF8C4,4);
TASK_PP(16'hF8C5,4);
TASK_PP(16'hF8C6,4);
TASK_PP(16'hF8C7,4);
TASK_PP(16'hF8C8,4);
TASK_PP(16'hF8C9,4);
TASK_PP(16'hF8CA,4);
TASK_PP(16'hF8CB,4);
TASK_PP(16'hF8CC,4);
TASK_PP(16'hF8CD,4);
TASK_PP(16'hF8CE,4);
TASK_PP(16'hF8CF,4);
TASK_PP(16'hF8D0,4);
TASK_PP(16'hF8D1,4);
TASK_PP(16'hF8D2,4);
TASK_PP(16'hF8D3,4);
TASK_PP(16'hF8D4,4);
TASK_PP(16'hF8D5,4);
TASK_PP(16'hF8D6,4);
TASK_PP(16'hF8D7,4);
TASK_PP(16'hF8D8,4);
TASK_PP(16'hF8D9,4);
TASK_PP(16'hF8DA,4);
TASK_PP(16'hF8DB,4);
TASK_PP(16'hF8DC,4);
TASK_PP(16'hF8DD,4);
TASK_PP(16'hF8DE,4);
TASK_PP(16'hF8DF,4);
TASK_PP(16'hF8E0,4);
TASK_PP(16'hF8E1,4);
TASK_PP(16'hF8E2,4);
TASK_PP(16'hF8E3,4);
TASK_PP(16'hF8E4,4);
TASK_PP(16'hF8E5,4);
TASK_PP(16'hF8E6,4);
TASK_PP(16'hF8E7,4);
TASK_PP(16'hF8E8,4);
TASK_PP(16'hF8E9,4);
TASK_PP(16'hF8EA,4);
TASK_PP(16'hF8EB,4);
TASK_PP(16'hF8EC,4);
TASK_PP(16'hF8ED,4);
TASK_PP(16'hF8EE,4);
TASK_PP(16'hF8EF,4);
TASK_PP(16'hF8F0,4);
TASK_PP(16'hF8F1,4);
TASK_PP(16'hF8F2,4);
TASK_PP(16'hF8F3,4);
TASK_PP(16'hF8F4,4);
TASK_PP(16'hF8F5,4);
TASK_PP(16'hF8F6,4);
TASK_PP(16'hF8F7,4);
TASK_PP(16'hF8F8,4);
TASK_PP(16'hF8F9,4);
TASK_PP(16'hF8FA,4);
TASK_PP(16'hF8FB,4);
TASK_PP(16'hF8FC,4);
TASK_PP(16'hF8FD,4);
TASK_PP(16'hF8FE,4);
TASK_PP(16'hF8FF,4);
TASK_PP(16'hF900,4);
TASK_PP(16'hF901,4);
TASK_PP(16'hF902,4);
TASK_PP(16'hF903,4);
TASK_PP(16'hF904,4);
TASK_PP(16'hF905,4);
TASK_PP(16'hF906,4);
TASK_PP(16'hF907,4);
TASK_PP(16'hF908,4);
TASK_PP(16'hF909,4);
TASK_PP(16'hF90A,4);
TASK_PP(16'hF90B,4);
TASK_PP(16'hF90C,4);
TASK_PP(16'hF90D,4);
TASK_PP(16'hF90E,4);
TASK_PP(16'hF90F,4);
TASK_PP(16'hF910,4);
TASK_PP(16'hF911,4);
TASK_PP(16'hF912,4);
TASK_PP(16'hF913,4);
TASK_PP(16'hF914,4);
TASK_PP(16'hF915,4);
TASK_PP(16'hF916,4);
TASK_PP(16'hF917,4);
TASK_PP(16'hF918,4);
TASK_PP(16'hF919,4);
TASK_PP(16'hF91A,4);
TASK_PP(16'hF91B,4);
TASK_PP(16'hF91C,4);
TASK_PP(16'hF91D,4);
TASK_PP(16'hF91E,4);
TASK_PP(16'hF91F,4);
TASK_PP(16'hF920,4);
TASK_PP(16'hF921,4);
TASK_PP(16'hF922,4);
TASK_PP(16'hF923,4);
TASK_PP(16'hF924,4);
TASK_PP(16'hF925,4);
TASK_PP(16'hF926,4);
TASK_PP(16'hF927,4);
TASK_PP(16'hF928,4);
TASK_PP(16'hF929,4);
TASK_PP(16'hF92A,4);
TASK_PP(16'hF92B,4);
TASK_PP(16'hF92C,4);
TASK_PP(16'hF92D,4);
TASK_PP(16'hF92E,4);
TASK_PP(16'hF92F,4);
TASK_PP(16'hF930,4);
TASK_PP(16'hF931,4);
TASK_PP(16'hF932,4);
TASK_PP(16'hF933,4);
TASK_PP(16'hF934,4);
TASK_PP(16'hF935,4);
TASK_PP(16'hF936,4);
TASK_PP(16'hF937,4);
TASK_PP(16'hF938,4);
TASK_PP(16'hF939,4);
TASK_PP(16'hF93A,4);
TASK_PP(16'hF93B,4);
TASK_PP(16'hF93C,4);
TASK_PP(16'hF93D,4);
TASK_PP(16'hF93E,4);
TASK_PP(16'hF93F,4);
TASK_PP(16'hF940,4);
TASK_PP(16'hF941,4);
TASK_PP(16'hF942,4);
TASK_PP(16'hF943,4);
TASK_PP(16'hF944,4);
TASK_PP(16'hF945,4);
TASK_PP(16'hF946,4);
TASK_PP(16'hF947,4);
TASK_PP(16'hF948,4);
TASK_PP(16'hF949,4);
TASK_PP(16'hF94A,4);
TASK_PP(16'hF94B,4);
TASK_PP(16'hF94C,4);
TASK_PP(16'hF94D,4);
TASK_PP(16'hF94E,4);
TASK_PP(16'hF94F,4);
TASK_PP(16'hF950,4);
TASK_PP(16'hF951,4);
TASK_PP(16'hF952,4);
TASK_PP(16'hF953,4);
TASK_PP(16'hF954,4);
TASK_PP(16'hF955,4);
TASK_PP(16'hF956,4);
TASK_PP(16'hF957,4);
TASK_PP(16'hF958,4);
TASK_PP(16'hF959,4);
TASK_PP(16'hF95A,4);
TASK_PP(16'hF95B,4);
TASK_PP(16'hF95C,4);
TASK_PP(16'hF95D,4);
TASK_PP(16'hF95E,4);
TASK_PP(16'hF95F,4);
TASK_PP(16'hF960,4);
TASK_PP(16'hF961,4);
TASK_PP(16'hF962,4);
TASK_PP(16'hF963,4);
TASK_PP(16'hF964,4);
TASK_PP(16'hF965,4);
TASK_PP(16'hF966,4);
TASK_PP(16'hF967,4);
TASK_PP(16'hF968,4);
TASK_PP(16'hF969,4);
TASK_PP(16'hF96A,4);
TASK_PP(16'hF96B,4);
TASK_PP(16'hF96C,4);
TASK_PP(16'hF96D,4);
TASK_PP(16'hF96E,4);
TASK_PP(16'hF96F,4);
TASK_PP(16'hF970,4);
TASK_PP(16'hF971,4);
TASK_PP(16'hF972,4);
TASK_PP(16'hF973,4);
TASK_PP(16'hF974,4);
TASK_PP(16'hF975,4);
TASK_PP(16'hF976,4);
TASK_PP(16'hF977,4);
TASK_PP(16'hF978,4);
TASK_PP(16'hF979,4);
TASK_PP(16'hF97A,4);
TASK_PP(16'hF97B,4);
TASK_PP(16'hF97C,4);
TASK_PP(16'hF97D,4);
TASK_PP(16'hF97E,4);
TASK_PP(16'hF97F,4);
TASK_PP(16'hF980,4);
TASK_PP(16'hF981,4);
TASK_PP(16'hF982,4);
TASK_PP(16'hF983,4);
TASK_PP(16'hF984,4);
TASK_PP(16'hF985,4);
TASK_PP(16'hF986,4);
TASK_PP(16'hF987,4);
TASK_PP(16'hF988,4);
TASK_PP(16'hF989,4);
TASK_PP(16'hF98A,4);
TASK_PP(16'hF98B,4);
TASK_PP(16'hF98C,4);
TASK_PP(16'hF98D,4);
TASK_PP(16'hF98E,4);
TASK_PP(16'hF98F,4);
TASK_PP(16'hF990,4);
TASK_PP(16'hF991,4);
TASK_PP(16'hF992,4);
TASK_PP(16'hF993,4);
TASK_PP(16'hF994,4);
TASK_PP(16'hF995,4);
TASK_PP(16'hF996,4);
TASK_PP(16'hF997,4);
TASK_PP(16'hF998,4);
TASK_PP(16'hF999,4);
TASK_PP(16'hF99A,4);
TASK_PP(16'hF99B,4);
TASK_PP(16'hF99C,4);
TASK_PP(16'hF99D,4);
TASK_PP(16'hF99E,4);
TASK_PP(16'hF99F,4);
TASK_PP(16'hF9A0,4);
TASK_PP(16'hF9A1,4);
TASK_PP(16'hF9A2,4);
TASK_PP(16'hF9A3,4);
TASK_PP(16'hF9A4,4);
TASK_PP(16'hF9A5,4);
TASK_PP(16'hF9A6,4);
TASK_PP(16'hF9A7,4);
TASK_PP(16'hF9A8,4);
TASK_PP(16'hF9A9,4);
TASK_PP(16'hF9AA,4);
TASK_PP(16'hF9AB,4);
TASK_PP(16'hF9AC,4);
TASK_PP(16'hF9AD,4);
TASK_PP(16'hF9AE,4);
TASK_PP(16'hF9AF,4);
TASK_PP(16'hF9B0,4);
TASK_PP(16'hF9B1,4);
TASK_PP(16'hF9B2,4);
TASK_PP(16'hF9B3,4);
TASK_PP(16'hF9B4,4);
TASK_PP(16'hF9B5,4);
TASK_PP(16'hF9B6,4);
TASK_PP(16'hF9B7,4);
TASK_PP(16'hF9B8,4);
TASK_PP(16'hF9B9,4);
TASK_PP(16'hF9BA,4);
TASK_PP(16'hF9BB,4);
TASK_PP(16'hF9BC,4);
TASK_PP(16'hF9BD,4);
TASK_PP(16'hF9BE,4);
TASK_PP(16'hF9BF,4);
TASK_PP(16'hF9C0,4);
TASK_PP(16'hF9C1,4);
TASK_PP(16'hF9C2,4);
TASK_PP(16'hF9C3,4);
TASK_PP(16'hF9C4,4);
TASK_PP(16'hF9C5,4);
TASK_PP(16'hF9C6,4);
TASK_PP(16'hF9C7,4);
TASK_PP(16'hF9C8,4);
TASK_PP(16'hF9C9,4);
TASK_PP(16'hF9CA,4);
TASK_PP(16'hF9CB,4);
TASK_PP(16'hF9CC,4);
TASK_PP(16'hF9CD,4);
TASK_PP(16'hF9CE,4);
TASK_PP(16'hF9CF,4);
TASK_PP(16'hF9D0,4);
TASK_PP(16'hF9D1,4);
TASK_PP(16'hF9D2,4);
TASK_PP(16'hF9D3,4);
TASK_PP(16'hF9D4,4);
TASK_PP(16'hF9D5,4);
TASK_PP(16'hF9D6,4);
TASK_PP(16'hF9D7,4);
TASK_PP(16'hF9D8,4);
TASK_PP(16'hF9D9,4);
TASK_PP(16'hF9DA,4);
TASK_PP(16'hF9DB,4);
TASK_PP(16'hF9DC,4);
TASK_PP(16'hF9DD,4);
TASK_PP(16'hF9DE,4);
TASK_PP(16'hF9DF,4);
TASK_PP(16'hF9E0,4);
TASK_PP(16'hF9E1,4);
TASK_PP(16'hF9E2,4);
TASK_PP(16'hF9E3,4);
TASK_PP(16'hF9E4,4);
TASK_PP(16'hF9E5,4);
TASK_PP(16'hF9E6,4);
TASK_PP(16'hF9E7,4);
TASK_PP(16'hF9E8,4);
TASK_PP(16'hF9E9,4);
TASK_PP(16'hF9EA,4);
TASK_PP(16'hF9EB,4);
TASK_PP(16'hF9EC,4);
TASK_PP(16'hF9ED,4);
TASK_PP(16'hF9EE,4);
TASK_PP(16'hF9EF,4);
TASK_PP(16'hF9F0,4);
TASK_PP(16'hF9F1,4);
TASK_PP(16'hF9F2,4);
TASK_PP(16'hF9F3,4);
TASK_PP(16'hF9F4,4);
TASK_PP(16'hF9F5,4);
TASK_PP(16'hF9F6,4);
TASK_PP(16'hF9F7,4);
TASK_PP(16'hF9F8,4);
TASK_PP(16'hF9F9,4);
TASK_PP(16'hF9FA,4);
TASK_PP(16'hF9FB,4);
TASK_PP(16'hF9FC,4);
TASK_PP(16'hF9FD,4);
TASK_PP(16'hF9FE,4);
TASK_PP(16'hF9FF,4);
TASK_PP(16'hFA00,4);
TASK_PP(16'hFA01,4);
TASK_PP(16'hFA02,4);
TASK_PP(16'hFA03,4);
TASK_PP(16'hFA04,4);
TASK_PP(16'hFA05,4);
TASK_PP(16'hFA06,4);
TASK_PP(16'hFA07,4);
TASK_PP(16'hFA08,4);
TASK_PP(16'hFA09,4);
TASK_PP(16'hFA0A,4);
TASK_PP(16'hFA0B,4);
TASK_PP(16'hFA0C,4);
TASK_PP(16'hFA0D,4);
TASK_PP(16'hFA0E,4);
TASK_PP(16'hFA0F,4);
TASK_PP(16'hFA10,4);
TASK_PP(16'hFA11,4);
TASK_PP(16'hFA12,4);
TASK_PP(16'hFA13,4);
TASK_PP(16'hFA14,4);
TASK_PP(16'hFA15,4);
TASK_PP(16'hFA16,4);
TASK_PP(16'hFA17,4);
TASK_PP(16'hFA18,4);
TASK_PP(16'hFA19,4);
TASK_PP(16'hFA1A,4);
TASK_PP(16'hFA1B,4);
TASK_PP(16'hFA1C,4);
TASK_PP(16'hFA1D,4);
TASK_PP(16'hFA1E,4);
TASK_PP(16'hFA1F,4);
TASK_PP(16'hFA20,4);
TASK_PP(16'hFA21,4);
TASK_PP(16'hFA22,4);
TASK_PP(16'hFA23,4);
TASK_PP(16'hFA24,4);
TASK_PP(16'hFA25,4);
TASK_PP(16'hFA26,4);
TASK_PP(16'hFA27,4);
TASK_PP(16'hFA28,4);
TASK_PP(16'hFA29,4);
TASK_PP(16'hFA2A,4);
TASK_PP(16'hFA2B,4);
TASK_PP(16'hFA2C,4);
TASK_PP(16'hFA2D,4);
TASK_PP(16'hFA2E,4);
TASK_PP(16'hFA2F,4);
TASK_PP(16'hFA30,4);
TASK_PP(16'hFA31,4);
TASK_PP(16'hFA32,4);
TASK_PP(16'hFA33,4);
TASK_PP(16'hFA34,4);
TASK_PP(16'hFA35,4);
TASK_PP(16'hFA36,4);
TASK_PP(16'hFA37,4);
TASK_PP(16'hFA38,4);
TASK_PP(16'hFA39,4);
TASK_PP(16'hFA3A,4);
TASK_PP(16'hFA3B,4);
TASK_PP(16'hFA3C,4);
TASK_PP(16'hFA3D,4);
TASK_PP(16'hFA3E,4);
TASK_PP(16'hFA3F,4);
TASK_PP(16'hFA40,4);
TASK_PP(16'hFA41,4);
TASK_PP(16'hFA42,4);
TASK_PP(16'hFA43,4);
TASK_PP(16'hFA44,4);
TASK_PP(16'hFA45,4);
TASK_PP(16'hFA46,4);
TASK_PP(16'hFA47,4);
TASK_PP(16'hFA48,4);
TASK_PP(16'hFA49,4);
TASK_PP(16'hFA4A,4);
TASK_PP(16'hFA4B,4);
TASK_PP(16'hFA4C,4);
TASK_PP(16'hFA4D,4);
TASK_PP(16'hFA4E,4);
TASK_PP(16'hFA4F,4);
TASK_PP(16'hFA50,4);
TASK_PP(16'hFA51,4);
TASK_PP(16'hFA52,4);
TASK_PP(16'hFA53,4);
TASK_PP(16'hFA54,4);
TASK_PP(16'hFA55,4);
TASK_PP(16'hFA56,4);
TASK_PP(16'hFA57,4);
TASK_PP(16'hFA58,4);
TASK_PP(16'hFA59,4);
TASK_PP(16'hFA5A,4);
TASK_PP(16'hFA5B,4);
TASK_PP(16'hFA5C,4);
TASK_PP(16'hFA5D,4);
TASK_PP(16'hFA5E,4);
TASK_PP(16'hFA5F,4);
TASK_PP(16'hFA60,4);
TASK_PP(16'hFA61,4);
TASK_PP(16'hFA62,4);
TASK_PP(16'hFA63,4);
TASK_PP(16'hFA64,4);
TASK_PP(16'hFA65,4);
TASK_PP(16'hFA66,4);
TASK_PP(16'hFA67,4);
TASK_PP(16'hFA68,4);
TASK_PP(16'hFA69,4);
TASK_PP(16'hFA6A,4);
TASK_PP(16'hFA6B,4);
TASK_PP(16'hFA6C,4);
TASK_PP(16'hFA6D,4);
TASK_PP(16'hFA6E,4);
TASK_PP(16'hFA6F,4);
TASK_PP(16'hFA70,4);
TASK_PP(16'hFA71,4);
TASK_PP(16'hFA72,4);
TASK_PP(16'hFA73,4);
TASK_PP(16'hFA74,4);
TASK_PP(16'hFA75,4);
TASK_PP(16'hFA76,4);
TASK_PP(16'hFA77,4);
TASK_PP(16'hFA78,4);
TASK_PP(16'hFA79,4);
TASK_PP(16'hFA7A,4);
TASK_PP(16'hFA7B,4);
TASK_PP(16'hFA7C,4);
TASK_PP(16'hFA7D,4);
TASK_PP(16'hFA7E,4);
TASK_PP(16'hFA7F,4);
TASK_PP(16'hFA80,4);
TASK_PP(16'hFA81,4);
TASK_PP(16'hFA82,4);
TASK_PP(16'hFA83,4);
TASK_PP(16'hFA84,4);
TASK_PP(16'hFA85,4);
TASK_PP(16'hFA86,4);
TASK_PP(16'hFA87,4);
TASK_PP(16'hFA88,4);
TASK_PP(16'hFA89,4);
TASK_PP(16'hFA8A,4);
TASK_PP(16'hFA8B,4);
TASK_PP(16'hFA8C,4);
TASK_PP(16'hFA8D,4);
TASK_PP(16'hFA8E,4);
TASK_PP(16'hFA8F,4);
TASK_PP(16'hFA90,4);
TASK_PP(16'hFA91,4);
TASK_PP(16'hFA92,4);
TASK_PP(16'hFA93,4);
TASK_PP(16'hFA94,4);
TASK_PP(16'hFA95,4);
TASK_PP(16'hFA96,4);
TASK_PP(16'hFA97,4);
TASK_PP(16'hFA98,4);
TASK_PP(16'hFA99,4);
TASK_PP(16'hFA9A,4);
TASK_PP(16'hFA9B,4);
TASK_PP(16'hFA9C,4);
TASK_PP(16'hFA9D,4);
TASK_PP(16'hFA9E,4);
TASK_PP(16'hFA9F,4);
TASK_PP(16'hFAA0,4);
TASK_PP(16'hFAA1,4);
TASK_PP(16'hFAA2,4);
TASK_PP(16'hFAA3,4);
TASK_PP(16'hFAA4,4);
TASK_PP(16'hFAA5,4);
TASK_PP(16'hFAA6,4);
TASK_PP(16'hFAA7,4);
TASK_PP(16'hFAA8,4);
TASK_PP(16'hFAA9,4);
TASK_PP(16'hFAAA,4);
TASK_PP(16'hFAAB,4);
TASK_PP(16'hFAAC,4);
TASK_PP(16'hFAAD,4);
TASK_PP(16'hFAAE,4);
TASK_PP(16'hFAAF,4);
TASK_PP(16'hFAB0,4);
TASK_PP(16'hFAB1,4);
TASK_PP(16'hFAB2,4);
TASK_PP(16'hFAB3,4);
TASK_PP(16'hFAB4,4);
TASK_PP(16'hFAB5,4);
TASK_PP(16'hFAB6,4);
TASK_PP(16'hFAB7,4);
TASK_PP(16'hFAB8,4);
TASK_PP(16'hFAB9,4);
TASK_PP(16'hFABA,4);
TASK_PP(16'hFABB,4);
TASK_PP(16'hFABC,4);
TASK_PP(16'hFABD,4);
TASK_PP(16'hFABE,4);
TASK_PP(16'hFABF,4);
TASK_PP(16'hFAC0,4);
TASK_PP(16'hFAC1,4);
TASK_PP(16'hFAC2,4);
TASK_PP(16'hFAC3,4);
TASK_PP(16'hFAC4,4);
TASK_PP(16'hFAC5,4);
TASK_PP(16'hFAC6,4);
TASK_PP(16'hFAC7,4);
TASK_PP(16'hFAC8,4);
TASK_PP(16'hFAC9,4);
TASK_PP(16'hFACA,4);
TASK_PP(16'hFACB,4);
TASK_PP(16'hFACC,4);
TASK_PP(16'hFACD,4);
TASK_PP(16'hFACE,4);
TASK_PP(16'hFACF,4);
TASK_PP(16'hFAD0,4);
TASK_PP(16'hFAD1,4);
TASK_PP(16'hFAD2,4);
TASK_PP(16'hFAD3,4);
TASK_PP(16'hFAD4,4);
TASK_PP(16'hFAD5,4);
TASK_PP(16'hFAD6,4);
TASK_PP(16'hFAD7,4);
TASK_PP(16'hFAD8,4);
TASK_PP(16'hFAD9,4);
TASK_PP(16'hFADA,4);
TASK_PP(16'hFADB,4);
TASK_PP(16'hFADC,4);
TASK_PP(16'hFADD,4);
TASK_PP(16'hFADE,4);
TASK_PP(16'hFADF,4);
TASK_PP(16'hFAE0,4);
TASK_PP(16'hFAE1,4);
TASK_PP(16'hFAE2,4);
TASK_PP(16'hFAE3,4);
TASK_PP(16'hFAE4,4);
TASK_PP(16'hFAE5,4);
TASK_PP(16'hFAE6,4);
TASK_PP(16'hFAE7,4);
TASK_PP(16'hFAE8,4);
TASK_PP(16'hFAE9,4);
TASK_PP(16'hFAEA,4);
TASK_PP(16'hFAEB,4);
TASK_PP(16'hFAEC,4);
TASK_PP(16'hFAED,4);
TASK_PP(16'hFAEE,4);
TASK_PP(16'hFAEF,4);
TASK_PP(16'hFAF0,4);
TASK_PP(16'hFAF1,4);
TASK_PP(16'hFAF2,4);
TASK_PP(16'hFAF3,4);
TASK_PP(16'hFAF4,4);
TASK_PP(16'hFAF5,4);
TASK_PP(16'hFAF6,4);
TASK_PP(16'hFAF7,4);
TASK_PP(16'hFAF8,4);
TASK_PP(16'hFAF9,4);
TASK_PP(16'hFAFA,4);
TASK_PP(16'hFAFB,4);
TASK_PP(16'hFAFC,4);
TASK_PP(16'hFAFD,4);
TASK_PP(16'hFAFE,4);
TASK_PP(16'hFAFF,4);
TASK_PP(16'hFB00,4);
TASK_PP(16'hFB01,4);
TASK_PP(16'hFB02,4);
TASK_PP(16'hFB03,4);
TASK_PP(16'hFB04,4);
TASK_PP(16'hFB05,4);
TASK_PP(16'hFB06,4);
TASK_PP(16'hFB07,4);
TASK_PP(16'hFB08,4);
TASK_PP(16'hFB09,4);
TASK_PP(16'hFB0A,4);
TASK_PP(16'hFB0B,4);
TASK_PP(16'hFB0C,4);
TASK_PP(16'hFB0D,4);
TASK_PP(16'hFB0E,4);
TASK_PP(16'hFB0F,4);
TASK_PP(16'hFB10,4);
TASK_PP(16'hFB11,4);
TASK_PP(16'hFB12,4);
TASK_PP(16'hFB13,4);
TASK_PP(16'hFB14,4);
TASK_PP(16'hFB15,4);
TASK_PP(16'hFB16,4);
TASK_PP(16'hFB17,4);
TASK_PP(16'hFB18,4);
TASK_PP(16'hFB19,4);
TASK_PP(16'hFB1A,4);
TASK_PP(16'hFB1B,4);
TASK_PP(16'hFB1C,4);
TASK_PP(16'hFB1D,4);
TASK_PP(16'hFB1E,4);
TASK_PP(16'hFB1F,4);
TASK_PP(16'hFB20,4);
TASK_PP(16'hFB21,4);
TASK_PP(16'hFB22,4);
TASK_PP(16'hFB23,4);
TASK_PP(16'hFB24,4);
TASK_PP(16'hFB25,4);
TASK_PP(16'hFB26,4);
TASK_PP(16'hFB27,4);
TASK_PP(16'hFB28,4);
TASK_PP(16'hFB29,4);
TASK_PP(16'hFB2A,4);
TASK_PP(16'hFB2B,4);
TASK_PP(16'hFB2C,4);
TASK_PP(16'hFB2D,4);
TASK_PP(16'hFB2E,4);
TASK_PP(16'hFB2F,4);
TASK_PP(16'hFB30,4);
TASK_PP(16'hFB31,4);
TASK_PP(16'hFB32,4);
TASK_PP(16'hFB33,4);
TASK_PP(16'hFB34,4);
TASK_PP(16'hFB35,4);
TASK_PP(16'hFB36,4);
TASK_PP(16'hFB37,4);
TASK_PP(16'hFB38,4);
TASK_PP(16'hFB39,4);
TASK_PP(16'hFB3A,4);
TASK_PP(16'hFB3B,4);
TASK_PP(16'hFB3C,4);
TASK_PP(16'hFB3D,4);
TASK_PP(16'hFB3E,4);
TASK_PP(16'hFB3F,4);
TASK_PP(16'hFB40,4);
TASK_PP(16'hFB41,4);
TASK_PP(16'hFB42,4);
TASK_PP(16'hFB43,4);
TASK_PP(16'hFB44,4);
TASK_PP(16'hFB45,4);
TASK_PP(16'hFB46,4);
TASK_PP(16'hFB47,4);
TASK_PP(16'hFB48,4);
TASK_PP(16'hFB49,4);
TASK_PP(16'hFB4A,4);
TASK_PP(16'hFB4B,4);
TASK_PP(16'hFB4C,4);
TASK_PP(16'hFB4D,4);
TASK_PP(16'hFB4E,4);
TASK_PP(16'hFB4F,4);
TASK_PP(16'hFB50,4);
TASK_PP(16'hFB51,4);
TASK_PP(16'hFB52,4);
TASK_PP(16'hFB53,4);
TASK_PP(16'hFB54,4);
TASK_PP(16'hFB55,4);
TASK_PP(16'hFB56,4);
TASK_PP(16'hFB57,4);
TASK_PP(16'hFB58,4);
TASK_PP(16'hFB59,4);
TASK_PP(16'hFB5A,4);
TASK_PP(16'hFB5B,4);
TASK_PP(16'hFB5C,4);
TASK_PP(16'hFB5D,4);
TASK_PP(16'hFB5E,4);
TASK_PP(16'hFB5F,4);
TASK_PP(16'hFB60,4);
TASK_PP(16'hFB61,4);
TASK_PP(16'hFB62,4);
TASK_PP(16'hFB63,4);
TASK_PP(16'hFB64,4);
TASK_PP(16'hFB65,4);
TASK_PP(16'hFB66,4);
TASK_PP(16'hFB67,4);
TASK_PP(16'hFB68,4);
TASK_PP(16'hFB69,4);
TASK_PP(16'hFB6A,4);
TASK_PP(16'hFB6B,4);
TASK_PP(16'hFB6C,4);
TASK_PP(16'hFB6D,4);
TASK_PP(16'hFB6E,4);
TASK_PP(16'hFB6F,4);
TASK_PP(16'hFB70,4);
TASK_PP(16'hFB71,4);
TASK_PP(16'hFB72,4);
TASK_PP(16'hFB73,4);
TASK_PP(16'hFB74,4);
TASK_PP(16'hFB75,4);
TASK_PP(16'hFB76,4);
TASK_PP(16'hFB77,4);
TASK_PP(16'hFB78,4);
TASK_PP(16'hFB79,4);
TASK_PP(16'hFB7A,4);
TASK_PP(16'hFB7B,4);
TASK_PP(16'hFB7C,4);
TASK_PP(16'hFB7D,4);
TASK_PP(16'hFB7E,4);
TASK_PP(16'hFB7F,4);
TASK_PP(16'hFB80,4);
TASK_PP(16'hFB81,4);
TASK_PP(16'hFB82,4);
TASK_PP(16'hFB83,4);
TASK_PP(16'hFB84,4);
TASK_PP(16'hFB85,4);
TASK_PP(16'hFB86,4);
TASK_PP(16'hFB87,4);
TASK_PP(16'hFB88,4);
TASK_PP(16'hFB89,4);
TASK_PP(16'hFB8A,4);
TASK_PP(16'hFB8B,4);
TASK_PP(16'hFB8C,4);
TASK_PP(16'hFB8D,4);
TASK_PP(16'hFB8E,4);
TASK_PP(16'hFB8F,4);
TASK_PP(16'hFB90,4);
TASK_PP(16'hFB91,4);
TASK_PP(16'hFB92,4);
TASK_PP(16'hFB93,4);
TASK_PP(16'hFB94,4);
TASK_PP(16'hFB95,4);
TASK_PP(16'hFB96,4);
TASK_PP(16'hFB97,4);
TASK_PP(16'hFB98,4);
TASK_PP(16'hFB99,4);
TASK_PP(16'hFB9A,4);
TASK_PP(16'hFB9B,4);
TASK_PP(16'hFB9C,4);
TASK_PP(16'hFB9D,4);
TASK_PP(16'hFB9E,4);
TASK_PP(16'hFB9F,4);
TASK_PP(16'hFBA0,4);
TASK_PP(16'hFBA1,4);
TASK_PP(16'hFBA2,4);
TASK_PP(16'hFBA3,4);
TASK_PP(16'hFBA4,4);
TASK_PP(16'hFBA5,4);
TASK_PP(16'hFBA6,4);
TASK_PP(16'hFBA7,4);
TASK_PP(16'hFBA8,4);
TASK_PP(16'hFBA9,4);
TASK_PP(16'hFBAA,4);
TASK_PP(16'hFBAB,4);
TASK_PP(16'hFBAC,4);
TASK_PP(16'hFBAD,4);
TASK_PP(16'hFBAE,4);
TASK_PP(16'hFBAF,4);
TASK_PP(16'hFBB0,4);
TASK_PP(16'hFBB1,4);
TASK_PP(16'hFBB2,4);
TASK_PP(16'hFBB3,4);
TASK_PP(16'hFBB4,4);
TASK_PP(16'hFBB5,4);
TASK_PP(16'hFBB6,4);
TASK_PP(16'hFBB7,4);
TASK_PP(16'hFBB8,4);
TASK_PP(16'hFBB9,4);
TASK_PP(16'hFBBA,4);
TASK_PP(16'hFBBB,4);
TASK_PP(16'hFBBC,4);
TASK_PP(16'hFBBD,4);
TASK_PP(16'hFBBE,4);
TASK_PP(16'hFBBF,4);
TASK_PP(16'hFBC0,4);
TASK_PP(16'hFBC1,4);
TASK_PP(16'hFBC2,4);
TASK_PP(16'hFBC3,4);
TASK_PP(16'hFBC4,4);
TASK_PP(16'hFBC5,4);
TASK_PP(16'hFBC6,4);
TASK_PP(16'hFBC7,4);
TASK_PP(16'hFBC8,4);
TASK_PP(16'hFBC9,4);
TASK_PP(16'hFBCA,4);
TASK_PP(16'hFBCB,4);
TASK_PP(16'hFBCC,4);
TASK_PP(16'hFBCD,4);
TASK_PP(16'hFBCE,4);
TASK_PP(16'hFBCF,4);
TASK_PP(16'hFBD0,4);
TASK_PP(16'hFBD1,4);
TASK_PP(16'hFBD2,4);
TASK_PP(16'hFBD3,4);
TASK_PP(16'hFBD4,4);
TASK_PP(16'hFBD5,4);
TASK_PP(16'hFBD6,4);
TASK_PP(16'hFBD7,4);
TASK_PP(16'hFBD8,4);
TASK_PP(16'hFBD9,4);
TASK_PP(16'hFBDA,4);
TASK_PP(16'hFBDB,4);
TASK_PP(16'hFBDC,4);
TASK_PP(16'hFBDD,4);
TASK_PP(16'hFBDE,4);
TASK_PP(16'hFBDF,4);
TASK_PP(16'hFBE0,4);
TASK_PP(16'hFBE1,4);
TASK_PP(16'hFBE2,4);
TASK_PP(16'hFBE3,4);
TASK_PP(16'hFBE4,4);
TASK_PP(16'hFBE5,4);
TASK_PP(16'hFBE6,4);
TASK_PP(16'hFBE7,4);
TASK_PP(16'hFBE8,4);
TASK_PP(16'hFBE9,4);
TASK_PP(16'hFBEA,4);
TASK_PP(16'hFBEB,4);
TASK_PP(16'hFBEC,4);
TASK_PP(16'hFBED,4);
TASK_PP(16'hFBEE,4);
TASK_PP(16'hFBEF,4);
TASK_PP(16'hFBF0,4);
TASK_PP(16'hFBF1,4);
TASK_PP(16'hFBF2,4);
TASK_PP(16'hFBF3,4);
TASK_PP(16'hFBF4,4);
TASK_PP(16'hFBF5,4);
TASK_PP(16'hFBF6,4);
TASK_PP(16'hFBF7,4);
TASK_PP(16'hFBF8,4);
TASK_PP(16'hFBF9,4);
TASK_PP(16'hFBFA,4);
TASK_PP(16'hFBFB,4);
TASK_PP(16'hFBFC,4);
TASK_PP(16'hFBFD,4);
TASK_PP(16'hFBFE,4);
TASK_PP(16'hFBFF,4);
TASK_PP(16'hFC00,4);
TASK_PP(16'hFC01,4);
TASK_PP(16'hFC02,4);
TASK_PP(16'hFC03,4);
TASK_PP(16'hFC04,4);
TASK_PP(16'hFC05,4);
TASK_PP(16'hFC06,4);
TASK_PP(16'hFC07,4);
TASK_PP(16'hFC08,4);
TASK_PP(16'hFC09,4);
TASK_PP(16'hFC0A,4);
TASK_PP(16'hFC0B,4);
TASK_PP(16'hFC0C,4);
TASK_PP(16'hFC0D,4);
TASK_PP(16'hFC0E,4);
TASK_PP(16'hFC0F,4);
TASK_PP(16'hFC10,4);
TASK_PP(16'hFC11,4);
TASK_PP(16'hFC12,4);
TASK_PP(16'hFC13,4);
TASK_PP(16'hFC14,4);
TASK_PP(16'hFC15,4);
TASK_PP(16'hFC16,4);
TASK_PP(16'hFC17,4);
TASK_PP(16'hFC18,4);
TASK_PP(16'hFC19,4);
TASK_PP(16'hFC1A,4);
TASK_PP(16'hFC1B,4);
TASK_PP(16'hFC1C,4);
TASK_PP(16'hFC1D,4);
TASK_PP(16'hFC1E,4);
TASK_PP(16'hFC1F,4);
TASK_PP(16'hFC20,4);
TASK_PP(16'hFC21,4);
TASK_PP(16'hFC22,4);
TASK_PP(16'hFC23,4);
TASK_PP(16'hFC24,4);
TASK_PP(16'hFC25,4);
TASK_PP(16'hFC26,4);
TASK_PP(16'hFC27,4);
TASK_PP(16'hFC28,4);
TASK_PP(16'hFC29,4);
TASK_PP(16'hFC2A,4);
TASK_PP(16'hFC2B,4);
TASK_PP(16'hFC2C,4);
TASK_PP(16'hFC2D,4);
TASK_PP(16'hFC2E,4);
TASK_PP(16'hFC2F,4);
TASK_PP(16'hFC30,4);
TASK_PP(16'hFC31,4);
TASK_PP(16'hFC32,4);
TASK_PP(16'hFC33,4);
TASK_PP(16'hFC34,4);
TASK_PP(16'hFC35,4);
TASK_PP(16'hFC36,4);
TASK_PP(16'hFC37,4);
TASK_PP(16'hFC38,4);
TASK_PP(16'hFC39,4);
TASK_PP(16'hFC3A,4);
TASK_PP(16'hFC3B,4);
TASK_PP(16'hFC3C,4);
TASK_PP(16'hFC3D,4);
TASK_PP(16'hFC3E,4);
TASK_PP(16'hFC3F,4);
TASK_PP(16'hFC40,4);
TASK_PP(16'hFC41,4);
TASK_PP(16'hFC42,4);
TASK_PP(16'hFC43,4);
TASK_PP(16'hFC44,4);
TASK_PP(16'hFC45,4);
TASK_PP(16'hFC46,4);
TASK_PP(16'hFC47,4);
TASK_PP(16'hFC48,4);
TASK_PP(16'hFC49,4);
TASK_PP(16'hFC4A,4);
TASK_PP(16'hFC4B,4);
TASK_PP(16'hFC4C,4);
TASK_PP(16'hFC4D,4);
TASK_PP(16'hFC4E,4);
TASK_PP(16'hFC4F,4);
TASK_PP(16'hFC50,4);
TASK_PP(16'hFC51,4);
TASK_PP(16'hFC52,4);
TASK_PP(16'hFC53,4);
TASK_PP(16'hFC54,4);
TASK_PP(16'hFC55,4);
TASK_PP(16'hFC56,4);
TASK_PP(16'hFC57,4);
TASK_PP(16'hFC58,4);
TASK_PP(16'hFC59,4);
TASK_PP(16'hFC5A,4);
TASK_PP(16'hFC5B,4);
TASK_PP(16'hFC5C,4);
TASK_PP(16'hFC5D,4);
TASK_PP(16'hFC5E,4);
TASK_PP(16'hFC5F,4);
TASK_PP(16'hFC60,4);
TASK_PP(16'hFC61,4);
TASK_PP(16'hFC62,4);
TASK_PP(16'hFC63,4);
TASK_PP(16'hFC64,4);
TASK_PP(16'hFC65,4);
TASK_PP(16'hFC66,4);
TASK_PP(16'hFC67,4);
TASK_PP(16'hFC68,4);
TASK_PP(16'hFC69,4);
TASK_PP(16'hFC6A,4);
TASK_PP(16'hFC6B,4);
TASK_PP(16'hFC6C,4);
TASK_PP(16'hFC6D,4);
TASK_PP(16'hFC6E,4);
TASK_PP(16'hFC6F,4);
TASK_PP(16'hFC70,4);
TASK_PP(16'hFC71,4);
TASK_PP(16'hFC72,4);
TASK_PP(16'hFC73,4);
TASK_PP(16'hFC74,4);
TASK_PP(16'hFC75,4);
TASK_PP(16'hFC76,4);
TASK_PP(16'hFC77,4);
TASK_PP(16'hFC78,4);
TASK_PP(16'hFC79,4);
TASK_PP(16'hFC7A,4);
TASK_PP(16'hFC7B,4);
TASK_PP(16'hFC7C,4);
TASK_PP(16'hFC7D,4);
TASK_PP(16'hFC7E,4);
TASK_PP(16'hFC7F,4);
TASK_PP(16'hFC80,4);
TASK_PP(16'hFC81,4);
TASK_PP(16'hFC82,4);
TASK_PP(16'hFC83,4);
TASK_PP(16'hFC84,4);
TASK_PP(16'hFC85,4);
TASK_PP(16'hFC86,4);
TASK_PP(16'hFC87,4);
TASK_PP(16'hFC88,4);
TASK_PP(16'hFC89,4);
TASK_PP(16'hFC8A,4);
TASK_PP(16'hFC8B,4);
TASK_PP(16'hFC8C,4);
TASK_PP(16'hFC8D,4);
TASK_PP(16'hFC8E,4);
TASK_PP(16'hFC8F,4);
TASK_PP(16'hFC90,4);
TASK_PP(16'hFC91,4);
TASK_PP(16'hFC92,4);
TASK_PP(16'hFC93,4);
TASK_PP(16'hFC94,4);
TASK_PP(16'hFC95,4);
TASK_PP(16'hFC96,4);
TASK_PP(16'hFC97,4);
TASK_PP(16'hFC98,4);
TASK_PP(16'hFC99,4);
TASK_PP(16'hFC9A,4);
TASK_PP(16'hFC9B,4);
TASK_PP(16'hFC9C,4);
TASK_PP(16'hFC9D,4);
TASK_PP(16'hFC9E,4);
TASK_PP(16'hFC9F,4);
TASK_PP(16'hFCA0,4);
TASK_PP(16'hFCA1,4);
TASK_PP(16'hFCA2,4);
TASK_PP(16'hFCA3,4);
TASK_PP(16'hFCA4,4);
TASK_PP(16'hFCA5,4);
TASK_PP(16'hFCA6,4);
TASK_PP(16'hFCA7,4);
TASK_PP(16'hFCA8,4);
TASK_PP(16'hFCA9,4);
TASK_PP(16'hFCAA,4);
TASK_PP(16'hFCAB,4);
TASK_PP(16'hFCAC,4);
TASK_PP(16'hFCAD,4);
TASK_PP(16'hFCAE,4);
TASK_PP(16'hFCAF,4);
TASK_PP(16'hFCB0,4);
TASK_PP(16'hFCB1,4);
TASK_PP(16'hFCB2,4);
TASK_PP(16'hFCB3,4);
TASK_PP(16'hFCB4,4);
TASK_PP(16'hFCB5,4);
TASK_PP(16'hFCB6,4);
TASK_PP(16'hFCB7,4);
TASK_PP(16'hFCB8,4);
TASK_PP(16'hFCB9,4);
TASK_PP(16'hFCBA,4);
TASK_PP(16'hFCBB,4);
TASK_PP(16'hFCBC,4);
TASK_PP(16'hFCBD,4);
TASK_PP(16'hFCBE,4);
TASK_PP(16'hFCBF,4);
TASK_PP(16'hFCC0,4);
TASK_PP(16'hFCC1,4);
TASK_PP(16'hFCC2,4);
TASK_PP(16'hFCC3,4);
TASK_PP(16'hFCC4,4);
TASK_PP(16'hFCC5,4);
TASK_PP(16'hFCC6,4);
TASK_PP(16'hFCC7,4);
TASK_PP(16'hFCC8,4);
TASK_PP(16'hFCC9,4);
TASK_PP(16'hFCCA,4);
TASK_PP(16'hFCCB,4);
TASK_PP(16'hFCCC,4);
TASK_PP(16'hFCCD,4);
TASK_PP(16'hFCCE,4);
TASK_PP(16'hFCCF,4);
TASK_PP(16'hFCD0,4);
TASK_PP(16'hFCD1,4);
TASK_PP(16'hFCD2,4);
TASK_PP(16'hFCD3,4);
TASK_PP(16'hFCD4,4);
TASK_PP(16'hFCD5,4);
TASK_PP(16'hFCD6,4);
TASK_PP(16'hFCD7,4);
TASK_PP(16'hFCD8,4);
TASK_PP(16'hFCD9,4);
TASK_PP(16'hFCDA,4);
TASK_PP(16'hFCDB,4);
TASK_PP(16'hFCDC,4);
TASK_PP(16'hFCDD,4);
TASK_PP(16'hFCDE,4);
TASK_PP(16'hFCDF,4);
TASK_PP(16'hFCE0,4);
TASK_PP(16'hFCE1,4);
TASK_PP(16'hFCE2,4);
TASK_PP(16'hFCE3,4);
TASK_PP(16'hFCE4,4);
TASK_PP(16'hFCE5,4);
TASK_PP(16'hFCE6,4);
TASK_PP(16'hFCE7,4);
TASK_PP(16'hFCE8,4);
TASK_PP(16'hFCE9,4);
TASK_PP(16'hFCEA,4);
TASK_PP(16'hFCEB,4);
TASK_PP(16'hFCEC,4);
TASK_PP(16'hFCED,4);
TASK_PP(16'hFCEE,4);
TASK_PP(16'hFCEF,4);
TASK_PP(16'hFCF0,4);
TASK_PP(16'hFCF1,4);
TASK_PP(16'hFCF2,4);
TASK_PP(16'hFCF3,4);
TASK_PP(16'hFCF4,4);
TASK_PP(16'hFCF5,4);
TASK_PP(16'hFCF6,4);
TASK_PP(16'hFCF7,4);
TASK_PP(16'hFCF8,4);
TASK_PP(16'hFCF9,4);
TASK_PP(16'hFCFA,4);
TASK_PP(16'hFCFB,4);
TASK_PP(16'hFCFC,4);
TASK_PP(16'hFCFD,4);
TASK_PP(16'hFCFE,4);
TASK_PP(16'hFCFF,4);
TASK_PP(16'hFD00,4);
TASK_PP(16'hFD01,4);
TASK_PP(16'hFD02,4);
TASK_PP(16'hFD03,4);
TASK_PP(16'hFD04,4);
TASK_PP(16'hFD05,4);
TASK_PP(16'hFD06,4);
TASK_PP(16'hFD07,4);
TASK_PP(16'hFD08,4);
TASK_PP(16'hFD09,4);
TASK_PP(16'hFD0A,4);
TASK_PP(16'hFD0B,4);
TASK_PP(16'hFD0C,4);
TASK_PP(16'hFD0D,4);
TASK_PP(16'hFD0E,4);
TASK_PP(16'hFD0F,4);
TASK_PP(16'hFD10,4);
TASK_PP(16'hFD11,4);
TASK_PP(16'hFD12,4);
TASK_PP(16'hFD13,4);
TASK_PP(16'hFD14,4);
TASK_PP(16'hFD15,4);
TASK_PP(16'hFD16,4);
TASK_PP(16'hFD17,4);
TASK_PP(16'hFD18,4);
TASK_PP(16'hFD19,4);
TASK_PP(16'hFD1A,4);
TASK_PP(16'hFD1B,4);
TASK_PP(16'hFD1C,4);
TASK_PP(16'hFD1D,4);
TASK_PP(16'hFD1E,4);
TASK_PP(16'hFD1F,4);
TASK_PP(16'hFD20,4);
TASK_PP(16'hFD21,4);
TASK_PP(16'hFD22,4);
TASK_PP(16'hFD23,4);
TASK_PP(16'hFD24,4);
TASK_PP(16'hFD25,4);
TASK_PP(16'hFD26,4);
TASK_PP(16'hFD27,4);
TASK_PP(16'hFD28,4);
TASK_PP(16'hFD29,4);
TASK_PP(16'hFD2A,4);
TASK_PP(16'hFD2B,4);
TASK_PP(16'hFD2C,4);
TASK_PP(16'hFD2D,4);
TASK_PP(16'hFD2E,4);
TASK_PP(16'hFD2F,4);
TASK_PP(16'hFD30,4);
TASK_PP(16'hFD31,4);
TASK_PP(16'hFD32,4);
TASK_PP(16'hFD33,4);
TASK_PP(16'hFD34,4);
TASK_PP(16'hFD35,4);
TASK_PP(16'hFD36,4);
TASK_PP(16'hFD37,4);
TASK_PP(16'hFD38,4);
TASK_PP(16'hFD39,4);
TASK_PP(16'hFD3A,4);
TASK_PP(16'hFD3B,4);
TASK_PP(16'hFD3C,4);
TASK_PP(16'hFD3D,4);
TASK_PP(16'hFD3E,4);
TASK_PP(16'hFD3F,4);
TASK_PP(16'hFD40,4);
TASK_PP(16'hFD41,4);
TASK_PP(16'hFD42,4);
TASK_PP(16'hFD43,4);
TASK_PP(16'hFD44,4);
TASK_PP(16'hFD45,4);
TASK_PP(16'hFD46,4);
TASK_PP(16'hFD47,4);
TASK_PP(16'hFD48,4);
TASK_PP(16'hFD49,4);
TASK_PP(16'hFD4A,4);
TASK_PP(16'hFD4B,4);
TASK_PP(16'hFD4C,4);
TASK_PP(16'hFD4D,4);
TASK_PP(16'hFD4E,4);
TASK_PP(16'hFD4F,4);
TASK_PP(16'hFD50,4);
TASK_PP(16'hFD51,4);
TASK_PP(16'hFD52,4);
TASK_PP(16'hFD53,4);
TASK_PP(16'hFD54,4);
TASK_PP(16'hFD55,4);
TASK_PP(16'hFD56,4);
TASK_PP(16'hFD57,4);
TASK_PP(16'hFD58,4);
TASK_PP(16'hFD59,4);
TASK_PP(16'hFD5A,4);
TASK_PP(16'hFD5B,4);
TASK_PP(16'hFD5C,4);
TASK_PP(16'hFD5D,4);
TASK_PP(16'hFD5E,4);
TASK_PP(16'hFD5F,4);
TASK_PP(16'hFD60,4);
TASK_PP(16'hFD61,4);
TASK_PP(16'hFD62,4);
TASK_PP(16'hFD63,4);
TASK_PP(16'hFD64,4);
TASK_PP(16'hFD65,4);
TASK_PP(16'hFD66,4);
TASK_PP(16'hFD67,4);
TASK_PP(16'hFD68,4);
TASK_PP(16'hFD69,4);
TASK_PP(16'hFD6A,4);
TASK_PP(16'hFD6B,4);
TASK_PP(16'hFD6C,4);
TASK_PP(16'hFD6D,4);
TASK_PP(16'hFD6E,4);
TASK_PP(16'hFD6F,4);
TASK_PP(16'hFD70,4);
TASK_PP(16'hFD71,4);
TASK_PP(16'hFD72,4);
TASK_PP(16'hFD73,4);
TASK_PP(16'hFD74,4);
TASK_PP(16'hFD75,4);
TASK_PP(16'hFD76,4);
TASK_PP(16'hFD77,4);
TASK_PP(16'hFD78,4);
TASK_PP(16'hFD79,4);
TASK_PP(16'hFD7A,4);
TASK_PP(16'hFD7B,4);
TASK_PP(16'hFD7C,4);
TASK_PP(16'hFD7D,4);
TASK_PP(16'hFD7E,4);
TASK_PP(16'hFD7F,4);
TASK_PP(16'hFD80,4);
TASK_PP(16'hFD81,4);
TASK_PP(16'hFD82,4);
TASK_PP(16'hFD83,4);
TASK_PP(16'hFD84,4);
TASK_PP(16'hFD85,4);
TASK_PP(16'hFD86,4);
TASK_PP(16'hFD87,4);
TASK_PP(16'hFD88,4);
TASK_PP(16'hFD89,4);
TASK_PP(16'hFD8A,4);
TASK_PP(16'hFD8B,4);
TASK_PP(16'hFD8C,4);
TASK_PP(16'hFD8D,4);
TASK_PP(16'hFD8E,4);
TASK_PP(16'hFD8F,4);
TASK_PP(16'hFD90,4);
TASK_PP(16'hFD91,4);
TASK_PP(16'hFD92,4);
TASK_PP(16'hFD93,4);
TASK_PP(16'hFD94,4);
TASK_PP(16'hFD95,4);
TASK_PP(16'hFD96,4);
TASK_PP(16'hFD97,4);
TASK_PP(16'hFD98,4);
TASK_PP(16'hFD99,4);
TASK_PP(16'hFD9A,4);
TASK_PP(16'hFD9B,4);
TASK_PP(16'hFD9C,4);
TASK_PP(16'hFD9D,4);
TASK_PP(16'hFD9E,4);
TASK_PP(16'hFD9F,4);
TASK_PP(16'hFDA0,4);
TASK_PP(16'hFDA1,4);
TASK_PP(16'hFDA2,4);
TASK_PP(16'hFDA3,4);
TASK_PP(16'hFDA4,4);
TASK_PP(16'hFDA5,4);
TASK_PP(16'hFDA6,4);
TASK_PP(16'hFDA7,4);
TASK_PP(16'hFDA8,4);
TASK_PP(16'hFDA9,4);
TASK_PP(16'hFDAA,4);
TASK_PP(16'hFDAB,4);
TASK_PP(16'hFDAC,4);
TASK_PP(16'hFDAD,4);
TASK_PP(16'hFDAE,4);
TASK_PP(16'hFDAF,4);
TASK_PP(16'hFDB0,4);
TASK_PP(16'hFDB1,4);
TASK_PP(16'hFDB2,4);
TASK_PP(16'hFDB3,4);
TASK_PP(16'hFDB4,4);
TASK_PP(16'hFDB5,4);
TASK_PP(16'hFDB6,4);
TASK_PP(16'hFDB7,4);
TASK_PP(16'hFDB8,4);
TASK_PP(16'hFDB9,4);
TASK_PP(16'hFDBA,4);
TASK_PP(16'hFDBB,4);
TASK_PP(16'hFDBC,4);
TASK_PP(16'hFDBD,4);
TASK_PP(16'hFDBE,4);
TASK_PP(16'hFDBF,4);
TASK_PP(16'hFDC0,4);
TASK_PP(16'hFDC1,4);
TASK_PP(16'hFDC2,4);
TASK_PP(16'hFDC3,4);
TASK_PP(16'hFDC4,4);
TASK_PP(16'hFDC5,4);
TASK_PP(16'hFDC6,4);
TASK_PP(16'hFDC7,4);
TASK_PP(16'hFDC8,4);
TASK_PP(16'hFDC9,4);
TASK_PP(16'hFDCA,4);
TASK_PP(16'hFDCB,4);
TASK_PP(16'hFDCC,4);
TASK_PP(16'hFDCD,4);
TASK_PP(16'hFDCE,4);
TASK_PP(16'hFDCF,4);
TASK_PP(16'hFDD0,4);
TASK_PP(16'hFDD1,4);
TASK_PP(16'hFDD2,4);
TASK_PP(16'hFDD3,4);
TASK_PP(16'hFDD4,4);
TASK_PP(16'hFDD5,4);
TASK_PP(16'hFDD6,4);
TASK_PP(16'hFDD7,4);
TASK_PP(16'hFDD8,4);
TASK_PP(16'hFDD9,4);
TASK_PP(16'hFDDA,4);
TASK_PP(16'hFDDB,4);
TASK_PP(16'hFDDC,4);
TASK_PP(16'hFDDD,4);
TASK_PP(16'hFDDE,4);
TASK_PP(16'hFDDF,4);
TASK_PP(16'hFDE0,4);
TASK_PP(16'hFDE1,4);
TASK_PP(16'hFDE2,4);
TASK_PP(16'hFDE3,4);
TASK_PP(16'hFDE4,4);
TASK_PP(16'hFDE5,4);
TASK_PP(16'hFDE6,4);
TASK_PP(16'hFDE7,4);
TASK_PP(16'hFDE8,4);
TASK_PP(16'hFDE9,4);
TASK_PP(16'hFDEA,4);
TASK_PP(16'hFDEB,4);
TASK_PP(16'hFDEC,4);
TASK_PP(16'hFDED,4);
TASK_PP(16'hFDEE,4);
TASK_PP(16'hFDEF,4);
TASK_PP(16'hFDF0,4);
TASK_PP(16'hFDF1,4);
TASK_PP(16'hFDF2,4);
TASK_PP(16'hFDF3,4);
TASK_PP(16'hFDF4,4);
TASK_PP(16'hFDF5,4);
TASK_PP(16'hFDF6,4);
TASK_PP(16'hFDF7,4);
TASK_PP(16'hFDF8,4);
TASK_PP(16'hFDF9,4);
TASK_PP(16'hFDFA,4);
TASK_PP(16'hFDFB,4);
TASK_PP(16'hFDFC,4);
TASK_PP(16'hFDFD,4);
TASK_PP(16'hFDFE,4);
TASK_PP(16'hFDFF,4);
TASK_PP(16'hFE00,4);
TASK_PP(16'hFE01,4);
TASK_PP(16'hFE02,4);
TASK_PP(16'hFE03,4);
TASK_PP(16'hFE04,4);
TASK_PP(16'hFE05,4);
TASK_PP(16'hFE06,4);
TASK_PP(16'hFE07,4);
TASK_PP(16'hFE08,4);
TASK_PP(16'hFE09,4);
TASK_PP(16'hFE0A,4);
TASK_PP(16'hFE0B,4);
TASK_PP(16'hFE0C,4);
TASK_PP(16'hFE0D,4);
TASK_PP(16'hFE0E,4);
TASK_PP(16'hFE0F,4);
TASK_PP(16'hFE10,4);
TASK_PP(16'hFE11,4);
TASK_PP(16'hFE12,4);
TASK_PP(16'hFE13,4);
TASK_PP(16'hFE14,4);
TASK_PP(16'hFE15,4);
TASK_PP(16'hFE16,4);
TASK_PP(16'hFE17,4);
TASK_PP(16'hFE18,4);
TASK_PP(16'hFE19,4);
TASK_PP(16'hFE1A,4);
TASK_PP(16'hFE1B,4);
TASK_PP(16'hFE1C,4);
TASK_PP(16'hFE1D,4);
TASK_PP(16'hFE1E,4);
TASK_PP(16'hFE1F,4);
TASK_PP(16'hFE20,4);
TASK_PP(16'hFE21,4);
TASK_PP(16'hFE22,4);
TASK_PP(16'hFE23,4);
TASK_PP(16'hFE24,4);
TASK_PP(16'hFE25,4);
TASK_PP(16'hFE26,4);
TASK_PP(16'hFE27,4);
TASK_PP(16'hFE28,4);
TASK_PP(16'hFE29,4);
TASK_PP(16'hFE2A,4);
TASK_PP(16'hFE2B,4);
TASK_PP(16'hFE2C,4);
TASK_PP(16'hFE2D,4);
TASK_PP(16'hFE2E,4);
TASK_PP(16'hFE2F,4);
TASK_PP(16'hFE30,4);
TASK_PP(16'hFE31,4);
TASK_PP(16'hFE32,4);
TASK_PP(16'hFE33,4);
TASK_PP(16'hFE34,4);
TASK_PP(16'hFE35,4);
TASK_PP(16'hFE36,4);
TASK_PP(16'hFE37,4);
TASK_PP(16'hFE38,4);
TASK_PP(16'hFE39,4);
TASK_PP(16'hFE3A,4);
TASK_PP(16'hFE3B,4);
TASK_PP(16'hFE3C,4);
TASK_PP(16'hFE3D,4);
TASK_PP(16'hFE3E,4);
TASK_PP(16'hFE3F,4);
TASK_PP(16'hFE40,4);
TASK_PP(16'hFE41,4);
TASK_PP(16'hFE42,4);
TASK_PP(16'hFE43,4);
TASK_PP(16'hFE44,4);
TASK_PP(16'hFE45,4);
TASK_PP(16'hFE46,4);
TASK_PP(16'hFE47,4);
TASK_PP(16'hFE48,4);
TASK_PP(16'hFE49,4);
TASK_PP(16'hFE4A,4);
TASK_PP(16'hFE4B,4);
TASK_PP(16'hFE4C,4);
TASK_PP(16'hFE4D,4);
TASK_PP(16'hFE4E,4);
TASK_PP(16'hFE4F,4);
TASK_PP(16'hFE50,4);
TASK_PP(16'hFE51,4);
TASK_PP(16'hFE52,4);
TASK_PP(16'hFE53,4);
TASK_PP(16'hFE54,4);
TASK_PP(16'hFE55,4);
TASK_PP(16'hFE56,4);
TASK_PP(16'hFE57,4);
TASK_PP(16'hFE58,4);
TASK_PP(16'hFE59,4);
TASK_PP(16'hFE5A,4);
TASK_PP(16'hFE5B,4);
TASK_PP(16'hFE5C,4);
TASK_PP(16'hFE5D,4);
TASK_PP(16'hFE5E,4);
TASK_PP(16'hFE5F,4);
TASK_PP(16'hFE60,4);
TASK_PP(16'hFE61,4);
TASK_PP(16'hFE62,4);
TASK_PP(16'hFE63,4);
TASK_PP(16'hFE64,4);
TASK_PP(16'hFE65,4);
TASK_PP(16'hFE66,4);
TASK_PP(16'hFE67,4);
TASK_PP(16'hFE68,4);
TASK_PP(16'hFE69,4);
TASK_PP(16'hFE6A,4);
TASK_PP(16'hFE6B,4);
TASK_PP(16'hFE6C,4);
TASK_PP(16'hFE6D,4);
TASK_PP(16'hFE6E,4);
TASK_PP(16'hFE6F,4);
TASK_PP(16'hFE70,4);
TASK_PP(16'hFE71,4);
TASK_PP(16'hFE72,4);
TASK_PP(16'hFE73,4);
TASK_PP(16'hFE74,4);
TASK_PP(16'hFE75,4);
TASK_PP(16'hFE76,4);
TASK_PP(16'hFE77,4);
TASK_PP(16'hFE78,4);
TASK_PP(16'hFE79,4);
TASK_PP(16'hFE7A,4);
TASK_PP(16'hFE7B,4);
TASK_PP(16'hFE7C,4);
TASK_PP(16'hFE7D,4);
TASK_PP(16'hFE7E,4);
TASK_PP(16'hFE7F,4);
TASK_PP(16'hFE80,4);
TASK_PP(16'hFE81,4);
TASK_PP(16'hFE82,4);
TASK_PP(16'hFE83,4);
TASK_PP(16'hFE84,4);
TASK_PP(16'hFE85,4);
TASK_PP(16'hFE86,4);
TASK_PP(16'hFE87,4);
TASK_PP(16'hFE88,4);
TASK_PP(16'hFE89,4);
TASK_PP(16'hFE8A,4);
TASK_PP(16'hFE8B,4);
TASK_PP(16'hFE8C,4);
TASK_PP(16'hFE8D,4);
TASK_PP(16'hFE8E,4);
TASK_PP(16'hFE8F,4);
TASK_PP(16'hFE90,4);
TASK_PP(16'hFE91,4);
TASK_PP(16'hFE92,4);
TASK_PP(16'hFE93,4);
TASK_PP(16'hFE94,4);
TASK_PP(16'hFE95,4);
TASK_PP(16'hFE96,4);
TASK_PP(16'hFE97,4);
TASK_PP(16'hFE98,4);
TASK_PP(16'hFE99,4);
TASK_PP(16'hFE9A,4);
TASK_PP(16'hFE9B,4);
TASK_PP(16'hFE9C,4);
TASK_PP(16'hFE9D,4);
TASK_PP(16'hFE9E,4);
TASK_PP(16'hFE9F,4);
TASK_PP(16'hFEA0,4);
TASK_PP(16'hFEA1,4);
TASK_PP(16'hFEA2,4);
TASK_PP(16'hFEA3,4);
TASK_PP(16'hFEA4,4);
TASK_PP(16'hFEA5,4);
TASK_PP(16'hFEA6,4);
TASK_PP(16'hFEA7,4);
TASK_PP(16'hFEA8,4);
TASK_PP(16'hFEA9,4);
TASK_PP(16'hFEAA,4);
TASK_PP(16'hFEAB,4);
TASK_PP(16'hFEAC,4);
TASK_PP(16'hFEAD,4);
TASK_PP(16'hFEAE,4);
TASK_PP(16'hFEAF,4);
TASK_PP(16'hFEB0,4);
TASK_PP(16'hFEB1,4);
TASK_PP(16'hFEB2,4);
TASK_PP(16'hFEB3,4);
TASK_PP(16'hFEB4,4);
TASK_PP(16'hFEB5,4);
TASK_PP(16'hFEB6,4);
TASK_PP(16'hFEB7,4);
TASK_PP(16'hFEB8,4);
TASK_PP(16'hFEB9,4);
TASK_PP(16'hFEBA,4);
TASK_PP(16'hFEBB,4);
TASK_PP(16'hFEBC,4);
TASK_PP(16'hFEBD,4);
TASK_PP(16'hFEBE,4);
TASK_PP(16'hFEBF,4);
TASK_PP(16'hFEC0,4);
TASK_PP(16'hFEC1,4);
TASK_PP(16'hFEC2,4);
TASK_PP(16'hFEC3,4);
TASK_PP(16'hFEC4,4);
TASK_PP(16'hFEC5,4);
TASK_PP(16'hFEC6,4);
TASK_PP(16'hFEC7,4);
TASK_PP(16'hFEC8,4);
TASK_PP(16'hFEC9,4);
TASK_PP(16'hFECA,4);
TASK_PP(16'hFECB,4);
TASK_PP(16'hFECC,4);
TASK_PP(16'hFECD,4);
TASK_PP(16'hFECE,4);
TASK_PP(16'hFECF,4);
TASK_PP(16'hFED0,4);
TASK_PP(16'hFED1,4);
TASK_PP(16'hFED2,4);
TASK_PP(16'hFED3,4);
TASK_PP(16'hFED4,4);
TASK_PP(16'hFED5,4);
TASK_PP(16'hFED6,4);
TASK_PP(16'hFED7,4);
TASK_PP(16'hFED8,4);
TASK_PP(16'hFED9,4);
TASK_PP(16'hFEDA,4);
TASK_PP(16'hFEDB,4);
TASK_PP(16'hFEDC,4);
TASK_PP(16'hFEDD,4);
TASK_PP(16'hFEDE,4);
TASK_PP(16'hFEDF,4);
TASK_PP(16'hFEE0,4);
TASK_PP(16'hFEE1,4);
TASK_PP(16'hFEE2,4);
TASK_PP(16'hFEE3,4);
TASK_PP(16'hFEE4,4);
TASK_PP(16'hFEE5,4);
TASK_PP(16'hFEE6,4);
TASK_PP(16'hFEE7,4);
TASK_PP(16'hFEE8,4);
TASK_PP(16'hFEE9,4);
TASK_PP(16'hFEEA,4);
TASK_PP(16'hFEEB,4);
TASK_PP(16'hFEEC,4);
TASK_PP(16'hFEED,4);
TASK_PP(16'hFEEE,4);
TASK_PP(16'hFEEF,4);
TASK_PP(16'hFEF0,4);
TASK_PP(16'hFEF1,4);
TASK_PP(16'hFEF2,4);
TASK_PP(16'hFEF3,4);
TASK_PP(16'hFEF4,4);
TASK_PP(16'hFEF5,4);
TASK_PP(16'hFEF6,4);
TASK_PP(16'hFEF7,4);
TASK_PP(16'hFEF8,4);
TASK_PP(16'hFEF9,4);
TASK_PP(16'hFEFA,4);
TASK_PP(16'hFEFB,4);
TASK_PP(16'hFEFC,4);
TASK_PP(16'hFEFD,4);
TASK_PP(16'hFEFE,4);
TASK_PP(16'hFEFF,4);
TASK_PP(16'hFF00,4);
TASK_PP(16'hFF01,4);
TASK_PP(16'hFF02,4);
TASK_PP(16'hFF03,4);
TASK_PP(16'hFF04,4);
TASK_PP(16'hFF05,4);
TASK_PP(16'hFF06,4);
TASK_PP(16'hFF07,4);
TASK_PP(16'hFF08,4);
TASK_PP(16'hFF09,4);
TASK_PP(16'hFF0A,4);
TASK_PP(16'hFF0B,4);
TASK_PP(16'hFF0C,4);
TASK_PP(16'hFF0D,4);
TASK_PP(16'hFF0E,4);
TASK_PP(16'hFF0F,4);
TASK_PP(16'hFF10,4);
TASK_PP(16'hFF11,4);
TASK_PP(16'hFF12,4);
TASK_PP(16'hFF13,4);
TASK_PP(16'hFF14,4);
TASK_PP(16'hFF15,4);
TASK_PP(16'hFF16,4);
TASK_PP(16'hFF17,4);
TASK_PP(16'hFF18,4);
TASK_PP(16'hFF19,4);
TASK_PP(16'hFF1A,4);
TASK_PP(16'hFF1B,4);
TASK_PP(16'hFF1C,4);
TASK_PP(16'hFF1D,4);
TASK_PP(16'hFF1E,4);
TASK_PP(16'hFF1F,4);
TASK_PP(16'hFF20,4);
TASK_PP(16'hFF21,4);
TASK_PP(16'hFF22,4);
TASK_PP(16'hFF23,4);
TASK_PP(16'hFF24,4);
TASK_PP(16'hFF25,4);
TASK_PP(16'hFF26,4);
TASK_PP(16'hFF27,4);
TASK_PP(16'hFF28,4);
TASK_PP(16'hFF29,4);
TASK_PP(16'hFF2A,4);
TASK_PP(16'hFF2B,4);
TASK_PP(16'hFF2C,4);
TASK_PP(16'hFF2D,4);
TASK_PP(16'hFF2E,4);
TASK_PP(16'hFF2F,4);
TASK_PP(16'hFF30,4);
TASK_PP(16'hFF31,4);
TASK_PP(16'hFF32,4);
TASK_PP(16'hFF33,4);
TASK_PP(16'hFF34,4);
TASK_PP(16'hFF35,4);
TASK_PP(16'hFF36,4);
TASK_PP(16'hFF37,4);
TASK_PP(16'hFF38,4);
TASK_PP(16'hFF39,4);
TASK_PP(16'hFF3A,4);
TASK_PP(16'hFF3B,4);
TASK_PP(16'hFF3C,4);
TASK_PP(16'hFF3D,4);
TASK_PP(16'hFF3E,4);
TASK_PP(16'hFF3F,4);
TASK_PP(16'hFF40,4);
TASK_PP(16'hFF41,4);
TASK_PP(16'hFF42,4);
TASK_PP(16'hFF43,4);
TASK_PP(16'hFF44,4);
TASK_PP(16'hFF45,4);
TASK_PP(16'hFF46,4);
TASK_PP(16'hFF47,4);
TASK_PP(16'hFF48,4);
TASK_PP(16'hFF49,4);
TASK_PP(16'hFF4A,4);
TASK_PP(16'hFF4B,4);
TASK_PP(16'hFF4C,4);
TASK_PP(16'hFF4D,4);
TASK_PP(16'hFF4E,4);
TASK_PP(16'hFF4F,4);
TASK_PP(16'hFF50,4);
TASK_PP(16'hFF51,4);
TASK_PP(16'hFF52,4);
TASK_PP(16'hFF53,4);
TASK_PP(16'hFF54,4);
TASK_PP(16'hFF55,4);
TASK_PP(16'hFF56,4);
TASK_PP(16'hFF57,4);
TASK_PP(16'hFF58,4);
TASK_PP(16'hFF59,4);
TASK_PP(16'hFF5A,4);
TASK_PP(16'hFF5B,4);
TASK_PP(16'hFF5C,4);
TASK_PP(16'hFF5D,4);
TASK_PP(16'hFF5E,4);
TASK_PP(16'hFF5F,4);
TASK_PP(16'hFF60,4);
TASK_PP(16'hFF61,4);
TASK_PP(16'hFF62,4);
TASK_PP(16'hFF63,4);
TASK_PP(16'hFF64,4);
TASK_PP(16'hFF65,4);
TASK_PP(16'hFF66,4);
TASK_PP(16'hFF67,4);
TASK_PP(16'hFF68,4);
TASK_PP(16'hFF69,4);
TASK_PP(16'hFF6A,4);
TASK_PP(16'hFF6B,4);
TASK_PP(16'hFF6C,4);
TASK_PP(16'hFF6D,4);
TASK_PP(16'hFF6E,4);
TASK_PP(16'hFF6F,4);
TASK_PP(16'hFF70,4);
TASK_PP(16'hFF71,4);
TASK_PP(16'hFF72,4);
TASK_PP(16'hFF73,4);
TASK_PP(16'hFF74,4);
TASK_PP(16'hFF75,4);
TASK_PP(16'hFF76,4);
TASK_PP(16'hFF77,4);
TASK_PP(16'hFF78,4);
TASK_PP(16'hFF79,4);
TASK_PP(16'hFF7A,4);
TASK_PP(16'hFF7B,4);
TASK_PP(16'hFF7C,4);
TASK_PP(16'hFF7D,4);
TASK_PP(16'hFF7E,4);
TASK_PP(16'hFF7F,4);
TASK_PP(16'hFF80,4);
TASK_PP(16'hFF81,4);
TASK_PP(16'hFF82,4);
TASK_PP(16'hFF83,4);
TASK_PP(16'hFF84,4);
TASK_PP(16'hFF85,4);
TASK_PP(16'hFF86,4);
TASK_PP(16'hFF87,4);
TASK_PP(16'hFF88,4);
TASK_PP(16'hFF89,4);
TASK_PP(16'hFF8A,4);
TASK_PP(16'hFF8B,4);
TASK_PP(16'hFF8C,4);
TASK_PP(16'hFF8D,4);
TASK_PP(16'hFF8E,4);
TASK_PP(16'hFF8F,4);
TASK_PP(16'hFF90,4);
TASK_PP(16'hFF91,4);
TASK_PP(16'hFF92,4);
TASK_PP(16'hFF93,4);
TASK_PP(16'hFF94,4);
TASK_PP(16'hFF95,4);
TASK_PP(16'hFF96,4);
TASK_PP(16'hFF97,4);
TASK_PP(16'hFF98,4);
TASK_PP(16'hFF99,4);
TASK_PP(16'hFF9A,4);
TASK_PP(16'hFF9B,4);
TASK_PP(16'hFF9C,4);
TASK_PP(16'hFF9D,4);
TASK_PP(16'hFF9E,4);
TASK_PP(16'hFF9F,4);
TASK_PP(16'hFFA0,4);
TASK_PP(16'hFFA1,4);
TASK_PP(16'hFFA2,4);
TASK_PP(16'hFFA3,4);
TASK_PP(16'hFFA4,4);
TASK_PP(16'hFFA5,4);
TASK_PP(16'hFFA6,4);
TASK_PP(16'hFFA7,4);
TASK_PP(16'hFFA8,4);
TASK_PP(16'hFFA9,4);
TASK_PP(16'hFFAA,4);
TASK_PP(16'hFFAB,4);
TASK_PP(16'hFFAC,4);
TASK_PP(16'hFFAD,4);
TASK_PP(16'hFFAE,4);
TASK_PP(16'hFFAF,4);
TASK_PP(16'hFFB0,4);
TASK_PP(16'hFFB1,4);
TASK_PP(16'hFFB2,4);
TASK_PP(16'hFFB3,4);
TASK_PP(16'hFFB4,4);
TASK_PP(16'hFFB5,4);
TASK_PP(16'hFFB6,4);
TASK_PP(16'hFFB7,4);
TASK_PP(16'hFFB8,4);
TASK_PP(16'hFFB9,4);
TASK_PP(16'hFFBA,4);
TASK_PP(16'hFFBB,4);
TASK_PP(16'hFFBC,4);
TASK_PP(16'hFFBD,4);
TASK_PP(16'hFFBE,4);
TASK_PP(16'hFFBF,4);
TASK_PP(16'hFFC0,4);
TASK_PP(16'hFFC1,4);
TASK_PP(16'hFFC2,4);
TASK_PP(16'hFFC3,4);
TASK_PP(16'hFFC4,4);
TASK_PP(16'hFFC5,4);
TASK_PP(16'hFFC6,4);
TASK_PP(16'hFFC7,4);
TASK_PP(16'hFFC8,4);
TASK_PP(16'hFFC9,4);
TASK_PP(16'hFFCA,4);
TASK_PP(16'hFFCB,4);
TASK_PP(16'hFFCC,4);
TASK_PP(16'hFFCD,4);
TASK_PP(16'hFFCE,4);
TASK_PP(16'hFFCF,4);
TASK_PP(16'hFFD0,4);
TASK_PP(16'hFFD1,4);
TASK_PP(16'hFFD2,4);
TASK_PP(16'hFFD3,4);
TASK_PP(16'hFFD4,4);
TASK_PP(16'hFFD5,4);
TASK_PP(16'hFFD6,4);
TASK_PP(16'hFFD7,4);
TASK_PP(16'hFFD8,4);
TASK_PP(16'hFFD9,4);
TASK_PP(16'hFFDA,4);
TASK_PP(16'hFFDB,4);
TASK_PP(16'hFFDC,4);
TASK_PP(16'hFFDD,4);
TASK_PP(16'hFFDE,4);
TASK_PP(16'hFFDF,4);
TASK_PP(16'hFFE0,4);
TASK_PP(16'hFFE1,4);
TASK_PP(16'hFFE2,4);
TASK_PP(16'hFFE3,4);
TASK_PP(16'hFFE4,4);
TASK_PP(16'hFFE5,4);
TASK_PP(16'hFFE6,4);
TASK_PP(16'hFFE7,4);
TASK_PP(16'hFFE8,4);
TASK_PP(16'hFFE9,4);
TASK_PP(16'hFFEA,4);
TASK_PP(16'hFFEB,4);
TASK_PP(16'hFFEC,4);
TASK_PP(16'hFFED,4);
TASK_PP(16'hFFEE,4);
TASK_PP(16'hFFEF,4);
TASK_PP(16'hFFF0,4);
TASK_PP(16'hFFF1,4);
TASK_PP(16'hFFF2,4);
TASK_PP(16'hFFF3,4);
TASK_PP(16'hFFF4,4);
TASK_PP(16'hFFF5,4);
TASK_PP(16'hFFF6,4);
TASK_PP(16'hFFF7,4);
TASK_PP(16'hFFF8,4);
TASK_PP(16'hFFF9,4);
TASK_PP(16'hFFFA,4);
TASK_PP(16'hFFFB,4);
TASK_PP(16'hFFFC,4);
TASK_PP(16'hFFFD,4);
TASK_PP(16'hFFFE,4);
TASK_PP(16'hFFFF,4);
TASK_PP(16'h10000,4);
TASK_PP(16'h10001,4);
TASK_PP(16'h10002,4);
TASK_PP(16'h10003,4);
TASK_PP(16'h10004,4);
TASK_PP(16'h10005,4);
TASK_PP(16'h10006,4);
TASK_PP(16'h10007,4);
TASK_PP(16'h10008,4);
TASK_PP(16'h10009,4);
TASK_PP(16'h1000A,4);
TASK_PP(16'h1000B,4);
TASK_PP(16'h1000C,4);
TASK_PP(16'h1000D,4);
TASK_PP(16'h1000E,4);
TASK_PP(16'h1000F,4);
TASK_PP(16'h10010,4);
TASK_PP(16'h10011,4);
TASK_PP(16'h10012,4);
TASK_PP(16'h10013,4);
TASK_PP(16'h10014,4);
TASK_PP(16'h10015,4);
TASK_PP(16'h10016,4);
TASK_PP(16'h10017,4);
TASK_PP(16'h10018,4);
TASK_PP(16'h10019,4);
TASK_PP(16'h1001A,4);
TASK_PP(16'h1001B,4);
TASK_PP(16'h1001C,4);
TASK_PP(16'h1001D,4);
TASK_PP(16'h1001E,4);
TASK_PP(16'h1001F,4);
TASK_PP(16'h10020,4);
TASK_PP(16'h10021,4);
TASK_PP(16'h10022,4);
TASK_PP(16'h10023,4);
TASK_PP(16'h10024,4);
TASK_PP(16'h10025,4);
TASK_PP(16'h10026,4);
TASK_PP(16'h10027,4);
TASK_PP(16'h10028,4);
TASK_PP(16'h10029,4);
TASK_PP(16'h1002A,4);
TASK_PP(16'h1002B,4);
TASK_PP(16'h1002C,4);
TASK_PP(16'h1002D,4);
TASK_PP(16'h1002E,4);
TASK_PP(16'h1002F,4);
TASK_PP(16'h10030,4);
TASK_PP(16'h10031,4);
TASK_PP(16'h10032,4);
TASK_PP(16'h10033,4);
TASK_PP(16'h10034,4);
TASK_PP(16'h10035,4);
TASK_PP(16'h10036,4);
TASK_PP(16'h10037,4);
TASK_PP(16'h10038,4);
TASK_PP(16'h10039,4);
TASK_PP(16'h1003A,4);
TASK_PP(16'h1003B,4);
TASK_PP(16'h1003C,4);
TASK_PP(16'h1003D,4);
TASK_PP(16'h1003E,4);
TASK_PP(16'h1003F,4);
TASK_PP(16'h10040,4);
TASK_PP(16'h10041,4);
TASK_PP(16'h10042,4);
TASK_PP(16'h10043,4);
TASK_PP(16'h10044,4);
TASK_PP(16'h10045,4);
TASK_PP(16'h10046,4);
TASK_PP(16'h10047,4);
TASK_PP(16'h10048,4);
TASK_PP(16'h10049,4);
TASK_PP(16'h1004A,4);
TASK_PP(16'h1004B,4);
TASK_PP(16'h1004C,4);
TASK_PP(16'h1004D,4);
TASK_PP(16'h1004E,4);
TASK_PP(16'h1004F,4);
TASK_PP(16'h10050,4);
TASK_PP(16'h10051,4);
TASK_PP(16'h10052,4);
TASK_PP(16'h10053,4);
TASK_PP(16'h10054,4);
TASK_PP(16'h10055,4);
TASK_PP(16'h10056,4);
TASK_PP(16'h10057,4);
TASK_PP(16'h10058,4);
TASK_PP(16'h10059,4);
TASK_PP(16'h1005A,4);
TASK_PP(16'h1005B,4);
TASK_PP(16'h1005C,4);
TASK_PP(16'h1005D,4);
TASK_PP(16'h1005E,4);
TASK_PP(16'h1005F,4);
TASK_PP(16'h10060,4);
TASK_PP(16'h10061,4);
TASK_PP(16'h10062,4);
TASK_PP(16'h10063,4);
TASK_PP(16'h10064,4);
TASK_PP(16'h10065,4);
TASK_PP(16'h10066,4);
TASK_PP(16'h10067,4);
TASK_PP(16'h10068,4);
TASK_PP(16'h10069,4);
TASK_PP(16'h1006A,4);
TASK_PP(16'h1006B,4);
TASK_PP(16'h1006C,4);
TASK_PP(16'h1006D,4);
TASK_PP(16'h1006E,4);
TASK_PP(16'h1006F,4);
TASK_PP(16'h10070,4);
TASK_PP(16'h10071,4);
TASK_PP(16'h10072,4);
TASK_PP(16'h10073,4);
TASK_PP(16'h10074,4);
TASK_PP(16'h10075,4);
TASK_PP(16'h10076,4);
TASK_PP(16'h10077,4);
TASK_PP(16'h10078,4);
TASK_PP(16'h10079,4);
TASK_PP(16'h1007A,4);
TASK_PP(16'h1007B,4);
TASK_PP(16'h1007C,4);
TASK_PP(16'h1007D,4);
TASK_PP(16'h1007E,4);
TASK_PP(16'h1007F,4);
TASK_PP(16'h10080,4);
TASK_PP(16'h10081,4);
TASK_PP(16'h10082,4);
TASK_PP(16'h10083,4);
TASK_PP(16'h10084,4);
TASK_PP(16'h10085,4);
TASK_PP(16'h10086,4);
TASK_PP(16'h10087,4);
TASK_PP(16'h10088,4);
TASK_PP(16'h10089,4);
TASK_PP(16'h1008A,4);
TASK_PP(16'h1008B,4);
TASK_PP(16'h1008C,4);
TASK_PP(16'h1008D,4);
TASK_PP(16'h1008E,4);
TASK_PP(16'h1008F,4);
TASK_PP(16'h10090,4);
TASK_PP(16'h10091,4);
TASK_PP(16'h10092,4);
TASK_PP(16'h10093,4);
TASK_PP(16'h10094,4);
TASK_PP(16'h10095,4);
TASK_PP(16'h10096,4);
TASK_PP(16'h10097,4);
TASK_PP(16'h10098,4);
TASK_PP(16'h10099,4);
TASK_PP(16'h1009A,4);
TASK_PP(16'h1009B,4);
TASK_PP(16'h1009C,4);
TASK_PP(16'h1009D,4);
TASK_PP(16'h1009E,4);
TASK_PP(16'h1009F,4);
TASK_PP(16'h100A0,4);
TASK_PP(16'h100A1,4);
TASK_PP(16'h100A2,4);
TASK_PP(16'h100A3,4);
TASK_PP(16'h100A4,4);
TASK_PP(16'h100A5,4);
TASK_PP(16'h100A6,4);
TASK_PP(16'h100A7,4);
TASK_PP(16'h100A8,4);
TASK_PP(16'h100A9,4);
TASK_PP(16'h100AA,4);
TASK_PP(16'h100AB,4);
TASK_PP(16'h100AC,4);
TASK_PP(16'h100AD,4);
TASK_PP(16'h100AE,4);
TASK_PP(16'h100AF,4);
TASK_PP(16'h100B0,4);
TASK_PP(16'h100B1,4);
TASK_PP(16'h100B2,4);
TASK_PP(16'h100B3,4);
TASK_PP(16'h100B4,4);
TASK_PP(16'h100B5,4);
TASK_PP(16'h100B6,4);
TASK_PP(16'h100B7,4);
TASK_PP(16'h100B8,4);
TASK_PP(16'h100B9,4);
TASK_PP(16'h100BA,4);
TASK_PP(16'h100BB,4);
TASK_PP(16'h100BC,4);
TASK_PP(16'h100BD,4);
TASK_PP(16'h100BE,4);
TASK_PP(16'h100BF,4);
TASK_PP(16'h100C0,4);
TASK_PP(16'h100C1,4);
TASK_PP(16'h100C2,4);
TASK_PP(16'h100C3,4);
TASK_PP(16'h100C4,4);
TASK_PP(16'h100C5,4);
TASK_PP(16'h100C6,4);
TASK_PP(16'h100C7,4);
TASK_PP(16'h100C8,4);
TASK_PP(16'h100C9,4);
TASK_PP(16'h100CA,4);
TASK_PP(16'h100CB,4);
TASK_PP(16'h100CC,4);
TASK_PP(16'h100CD,4);
TASK_PP(16'h100CE,4);
TASK_PP(16'h100CF,4);
TASK_PP(16'h100D0,4);
TASK_PP(16'h100D1,4);
TASK_PP(16'h100D2,4);
TASK_PP(16'h100D3,4);
TASK_PP(16'h100D4,4);
TASK_PP(16'h100D5,4);
TASK_PP(16'h100D6,4);
TASK_PP(16'h100D7,4);
TASK_PP(16'h100D8,4);
TASK_PP(16'h100D9,4);
TASK_PP(16'h100DA,4);
TASK_PP(16'h100DB,4);
TASK_PP(16'h100DC,4);
TASK_PP(16'h100DD,4);
TASK_PP(16'h100DE,4);
TASK_PP(16'h100DF,4);
TASK_PP(16'h100E0,4);
TASK_PP(16'h100E1,4);
TASK_PP(16'h100E2,4);
TASK_PP(16'h100E3,4);
TASK_PP(16'h100E4,4);
TASK_PP(16'h100E5,4);
TASK_PP(16'h100E6,4);
TASK_PP(16'h100E7,4);
TASK_PP(16'h100E8,4);
TASK_PP(16'h100E9,4);
TASK_PP(16'h100EA,4);
TASK_PP(16'h100EB,4);
TASK_PP(16'h100EC,4);
TASK_PP(16'h100ED,4);
TASK_PP(16'h100EE,4);
TASK_PP(16'h100EF,4);
TASK_PP(16'h100F0,4);
TASK_PP(16'h100F1,4);
TASK_PP(16'h100F2,4);
TASK_PP(16'h100F3,4);
TASK_PP(16'h100F4,4);
TASK_PP(16'h100F5,4);
TASK_PP(16'h100F6,4);
TASK_PP(16'h100F7,4);
TASK_PP(16'h100F8,4);
TASK_PP(16'h100F9,4);
TASK_PP(16'h100FA,4);
TASK_PP(16'h100FB,4);
TASK_PP(16'h100FC,4);
TASK_PP(16'h100FD,4);
TASK_PP(16'h100FE,4);
TASK_PP(16'h100FF,4);
TASK_PP(16'h10100,4);
TASK_PP(16'h10101,4);
TASK_PP(16'h10102,4);
TASK_PP(16'h10103,4);
TASK_PP(16'h10104,4);
TASK_PP(16'h10105,4);
TASK_PP(16'h10106,4);
TASK_PP(16'h10107,4);
TASK_PP(16'h10108,4);
TASK_PP(16'h10109,4);
TASK_PP(16'h1010A,4);
TASK_PP(16'h1010B,4);
TASK_PP(16'h1010C,4);
TASK_PP(16'h1010D,4);
TASK_PP(16'h1010E,4);
TASK_PP(16'h1010F,4);
TASK_PP(16'h10110,4);
TASK_PP(16'h10111,4);
TASK_PP(16'h10112,4);
TASK_PP(16'h10113,4);
TASK_PP(16'h10114,4);
TASK_PP(16'h10115,4);
TASK_PP(16'h10116,4);
TASK_PP(16'h10117,4);
TASK_PP(16'h10118,4);
TASK_PP(16'h10119,4);
TASK_PP(16'h1011A,4);
TASK_PP(16'h1011B,4);
TASK_PP(16'h1011C,4);
TASK_PP(16'h1011D,4);
TASK_PP(16'h1011E,4);
TASK_PP(16'h1011F,4);
TASK_PP(16'h10120,4);
TASK_PP(16'h10121,4);
TASK_PP(16'h10122,4);
TASK_PP(16'h10123,4);
TASK_PP(16'h10124,4);
TASK_PP(16'h10125,4);
TASK_PP(16'h10126,4);
TASK_PP(16'h10127,4);
TASK_PP(16'h10128,4);
TASK_PP(16'h10129,4);
TASK_PP(16'h1012A,4);
TASK_PP(16'h1012B,4);
TASK_PP(16'h1012C,4);
TASK_PP(16'h1012D,4);
TASK_PP(16'h1012E,4);
TASK_PP(16'h1012F,4);
TASK_PP(16'h10130,4);
TASK_PP(16'h10131,4);
TASK_PP(16'h10132,4);
TASK_PP(16'h10133,4);
TASK_PP(16'h10134,4);
TASK_PP(16'h10135,4);
TASK_PP(16'h10136,4);
TASK_PP(16'h10137,4);
TASK_PP(16'h10138,4);
TASK_PP(16'h10139,4);
TASK_PP(16'h1013A,4);
TASK_PP(16'h1013B,4);
TASK_PP(16'h1013C,4);
TASK_PP(16'h1013D,4);
TASK_PP(16'h1013E,4);
TASK_PP(16'h1013F,4);
TASK_PP(16'h10140,4);
TASK_PP(16'h10141,4);
TASK_PP(16'h10142,4);
TASK_PP(16'h10143,4);
TASK_PP(16'h10144,4);
TASK_PP(16'h10145,4);
TASK_PP(16'h10146,4);
TASK_PP(16'h10147,4);
TASK_PP(16'h10148,4);
TASK_PP(16'h10149,4);
TASK_PP(16'h1014A,4);
TASK_PP(16'h1014B,4);
TASK_PP(16'h1014C,4);
TASK_PP(16'h1014D,4);
TASK_PP(16'h1014E,4);
TASK_PP(16'h1014F,4);
TASK_PP(16'h10150,4);
TASK_PP(16'h10151,4);
TASK_PP(16'h10152,4);
TASK_PP(16'h10153,4);
TASK_PP(16'h10154,4);
TASK_PP(16'h10155,4);
TASK_PP(16'h10156,4);
TASK_PP(16'h10157,4);
TASK_PP(16'h10158,4);
TASK_PP(16'h10159,4);
TASK_PP(16'h1015A,4);
TASK_PP(16'h1015B,4);
TASK_PP(16'h1015C,4);
TASK_PP(16'h1015D,4);
TASK_PP(16'h1015E,4);
TASK_PP(16'h1015F,4);
TASK_PP(16'h10160,4);
TASK_PP(16'h10161,4);
TASK_PP(16'h10162,4);
TASK_PP(16'h10163,4);
TASK_PP(16'h10164,4);
TASK_PP(16'h10165,4);
TASK_PP(16'h10166,4);
TASK_PP(16'h10167,4);
TASK_PP(16'h10168,4);
TASK_PP(16'h10169,4);
TASK_PP(16'h1016A,4);
TASK_PP(16'h1016B,4);
TASK_PP(16'h1016C,4);
TASK_PP(16'h1016D,4);
TASK_PP(16'h1016E,4);
TASK_PP(16'h1016F,4);
TASK_PP(16'h10170,4);
TASK_PP(16'h10171,4);
TASK_PP(16'h10172,4);
TASK_PP(16'h10173,4);
TASK_PP(16'h10174,4);
TASK_PP(16'h10175,4);
TASK_PP(16'h10176,4);
TASK_PP(16'h10177,4);
TASK_PP(16'h10178,4);
TASK_PP(16'h10179,4);
TASK_PP(16'h1017A,4);
TASK_PP(16'h1017B,4);
TASK_PP(16'h1017C,4);
TASK_PP(16'h1017D,4);
TASK_PP(16'h1017E,4);
TASK_PP(16'h1017F,4);
TASK_PP(16'h10180,4);
TASK_PP(16'h10181,4);
TASK_PP(16'h10182,4);
TASK_PP(16'h10183,4);
TASK_PP(16'h10184,4);
TASK_PP(16'h10185,4);
TASK_PP(16'h10186,4);
TASK_PP(16'h10187,4);
TASK_PP(16'h10188,4);
TASK_PP(16'h10189,4);
TASK_PP(16'h1018A,4);
TASK_PP(16'h1018B,4);
TASK_PP(16'h1018C,4);
TASK_PP(16'h1018D,4);
TASK_PP(16'h1018E,4);
TASK_PP(16'h1018F,4);
TASK_PP(16'h10190,4);
TASK_PP(16'h10191,4);
TASK_PP(16'h10192,4);
TASK_PP(16'h10193,4);
TASK_PP(16'h10194,4);
TASK_PP(16'h10195,4);
TASK_PP(16'h10196,4);
TASK_PP(16'h10197,4);
TASK_PP(16'h10198,4);
TASK_PP(16'h10199,4);
TASK_PP(16'h1019A,4);
TASK_PP(16'h1019B,4);
TASK_PP(16'h1019C,4);
TASK_PP(16'h1019D,4);
TASK_PP(16'h1019E,4);
TASK_PP(16'h1019F,4);
TASK_PP(16'h101A0,4);
TASK_PP(16'h101A1,4);
TASK_PP(16'h101A2,4);
TASK_PP(16'h101A3,4);
TASK_PP(16'h101A4,4);
TASK_PP(16'h101A5,4);
TASK_PP(16'h101A6,4);
TASK_PP(16'h101A7,4);
TASK_PP(16'h101A8,4);
TASK_PP(16'h101A9,4);
TASK_PP(16'h101AA,4);
TASK_PP(16'h101AB,4);
TASK_PP(16'h101AC,4);
TASK_PP(16'h101AD,4);
TASK_PP(16'h101AE,4);
TASK_PP(16'h101AF,4);
TASK_PP(16'h101B0,4);
TASK_PP(16'h101B1,4);
TASK_PP(16'h101B2,4);
TASK_PP(16'h101B3,4);
TASK_PP(16'h101B4,4);
TASK_PP(16'h101B5,4);
TASK_PP(16'h101B6,4);
TASK_PP(16'h101B7,4);
TASK_PP(16'h101B8,4);
TASK_PP(16'h101B9,4);
TASK_PP(16'h101BA,4);
TASK_PP(16'h101BB,4);
TASK_PP(16'h101BC,4);
TASK_PP(16'h101BD,4);
TASK_PP(16'h101BE,4);
TASK_PP(16'h101BF,4);
TASK_PP(16'h101C0,4);
TASK_PP(16'h101C1,4);
TASK_PP(16'h101C2,4);
TASK_PP(16'h101C3,4);
TASK_PP(16'h101C4,4);
TASK_PP(16'h101C5,4);
TASK_PP(16'h101C6,4);
TASK_PP(16'h101C7,4);
TASK_PP(16'h101C8,4);
TASK_PP(16'h101C9,4);
TASK_PP(16'h101CA,4);
TASK_PP(16'h101CB,4);
TASK_PP(16'h101CC,4);
TASK_PP(16'h101CD,4);
TASK_PP(16'h101CE,4);
TASK_PP(16'h101CF,4);
TASK_PP(16'h101D0,4);
TASK_PP(16'h101D1,4);
TASK_PP(16'h101D2,4);
TASK_PP(16'h101D3,4);
TASK_PP(16'h101D4,4);
TASK_PP(16'h101D5,4);
TASK_PP(16'h101D6,4);
TASK_PP(16'h101D7,4);
TASK_PP(16'h101D8,4);
TASK_PP(16'h101D9,4);
TASK_PP(16'h101DA,4);
TASK_PP(16'h101DB,4);
TASK_PP(16'h101DC,4);
TASK_PP(16'h101DD,4);
TASK_PP(16'h101DE,4);
TASK_PP(16'h101DF,4);
TASK_PP(16'h101E0,4);
TASK_PP(16'h101E1,4);
TASK_PP(16'h101E2,4);
TASK_PP(16'h101E3,4);
TASK_PP(16'h101E4,4);
TASK_PP(16'h101E5,4);
TASK_PP(16'h101E6,4);
TASK_PP(16'h101E7,4);
TASK_PP(16'h101E8,4);
TASK_PP(16'h101E9,4);
TASK_PP(16'h101EA,4);
TASK_PP(16'h101EB,4);
TASK_PP(16'h101EC,4);
TASK_PP(16'h101ED,4);
TASK_PP(16'h101EE,4);
TASK_PP(16'h101EF,4);
TASK_PP(16'h101F0,4);
TASK_PP(16'h101F1,4);
TASK_PP(16'h101F2,4);
TASK_PP(16'h101F3,4);
TASK_PP(16'h101F4,4);
TASK_PP(16'h101F5,4);
TASK_PP(16'h101F6,4);
TASK_PP(16'h101F7,4);
TASK_PP(16'h101F8,4);
TASK_PP(16'h101F9,4);
TASK_PP(16'h101FA,4);
TASK_PP(16'h101FB,4);
TASK_PP(16'h101FC,4);
TASK_PP(16'h101FD,4);
TASK_PP(16'h101FE,4);
TASK_PP(16'h101FF,4);
TASK_PP(16'h10200,4);
TASK_PP(16'h10201,4);
TASK_PP(16'h10202,4);
TASK_PP(16'h10203,4);
TASK_PP(16'h10204,4);
TASK_PP(16'h10205,4);
TASK_PP(16'h10206,4);
TASK_PP(16'h10207,4);
TASK_PP(16'h10208,4);
TASK_PP(16'h10209,4);
TASK_PP(16'h1020A,4);
TASK_PP(16'h1020B,4);
TASK_PP(16'h1020C,4);
TASK_PP(16'h1020D,4);
TASK_PP(16'h1020E,4);
TASK_PP(16'h1020F,4);
TASK_PP(16'h10210,4);
TASK_PP(16'h10211,4);
TASK_PP(16'h10212,4);
TASK_PP(16'h10213,4);
TASK_PP(16'h10214,4);
TASK_PP(16'h10215,4);
TASK_PP(16'h10216,4);
TASK_PP(16'h10217,4);
TASK_PP(16'h10218,4);
TASK_PP(16'h10219,4);
TASK_PP(16'h1021A,4);
TASK_PP(16'h1021B,4);
TASK_PP(16'h1021C,4);
TASK_PP(16'h1021D,4);
TASK_PP(16'h1021E,4);
TASK_PP(16'h1021F,4);
TASK_PP(16'h10220,4);
TASK_PP(16'h10221,4);
TASK_PP(16'h10222,4);
TASK_PP(16'h10223,4);
TASK_PP(16'h10224,4);
TASK_PP(16'h10225,4);
TASK_PP(16'h10226,4);
TASK_PP(16'h10227,4);
TASK_PP(16'h10228,4);
TASK_PP(16'h10229,4);
TASK_PP(16'h1022A,4);
TASK_PP(16'h1022B,4);
TASK_PP(16'h1022C,4);
TASK_PP(16'h1022D,4);
TASK_PP(16'h1022E,4);
TASK_PP(16'h1022F,4);
TASK_PP(16'h10230,4);
TASK_PP(16'h10231,4);
TASK_PP(16'h10232,4);
TASK_PP(16'h10233,4);
TASK_PP(16'h10234,4);
TASK_PP(16'h10235,4);
TASK_PP(16'h10236,4);
TASK_PP(16'h10237,4);
TASK_PP(16'h10238,4);
TASK_PP(16'h10239,4);
TASK_PP(16'h1023A,4);
TASK_PP(16'h1023B,4);
TASK_PP(16'h1023C,4);
TASK_PP(16'h1023D,4);
TASK_PP(16'h1023E,4);
TASK_PP(16'h1023F,4);
TASK_PP(16'h10240,4);
TASK_PP(16'h10241,4);
TASK_PP(16'h10242,4);
TASK_PP(16'h10243,4);
TASK_PP(16'h10244,4);
TASK_PP(16'h10245,4);
TASK_PP(16'h10246,4);
TASK_PP(16'h10247,4);
TASK_PP(16'h10248,4);
TASK_PP(16'h10249,4);
TASK_PP(16'h1024A,4);
TASK_PP(16'h1024B,4);
TASK_PP(16'h1024C,4);
TASK_PP(16'h1024D,4);
TASK_PP(16'h1024E,4);
TASK_PP(16'h1024F,4);
TASK_PP(16'h10250,4);
TASK_PP(16'h10251,4);
TASK_PP(16'h10252,4);
TASK_PP(16'h10253,4);
TASK_PP(16'h10254,4);
TASK_PP(16'h10255,4);
TASK_PP(16'h10256,4);
TASK_PP(16'h10257,4);
TASK_PP(16'h10258,4);
TASK_PP(16'h10259,4);
TASK_PP(16'h1025A,4);
TASK_PP(16'h1025B,4);
TASK_PP(16'h1025C,4);
TASK_PP(16'h1025D,4);
TASK_PP(16'h1025E,4);
TASK_PP(16'h1025F,4);
TASK_PP(16'h10260,4);
TASK_PP(16'h10261,4);
TASK_PP(16'h10262,4);
TASK_PP(16'h10263,4);
TASK_PP(16'h10264,4);
TASK_PP(16'h10265,4);
TASK_PP(16'h10266,4);
TASK_PP(16'h10267,4);
TASK_PP(16'h10268,4);
TASK_PP(16'h10269,4);
TASK_PP(16'h1026A,4);
TASK_PP(16'h1026B,4);
TASK_PP(16'h1026C,4);
TASK_PP(16'h1026D,4);
TASK_PP(16'h1026E,4);
TASK_PP(16'h1026F,4);
TASK_PP(16'h10270,4);
TASK_PP(16'h10271,4);
TASK_PP(16'h10272,4);
TASK_PP(16'h10273,4);
TASK_PP(16'h10274,4);
TASK_PP(16'h10275,4);
TASK_PP(16'h10276,4);
TASK_PP(16'h10277,4);
TASK_PP(16'h10278,4);
TASK_PP(16'h10279,4);
TASK_PP(16'h1027A,4);
TASK_PP(16'h1027B,4);
TASK_PP(16'h1027C,4);
TASK_PP(16'h1027D,4);
TASK_PP(16'h1027E,4);
TASK_PP(16'h1027F,4);
TASK_PP(16'h10280,4);
TASK_PP(16'h10281,4);
TASK_PP(16'h10282,4);
TASK_PP(16'h10283,4);
TASK_PP(16'h10284,4);
TASK_PP(16'h10285,4);
TASK_PP(16'h10286,4);
TASK_PP(16'h10287,4);
TASK_PP(16'h10288,4);
TASK_PP(16'h10289,4);
TASK_PP(16'h1028A,4);
TASK_PP(16'h1028B,4);
TASK_PP(16'h1028C,4);
TASK_PP(16'h1028D,4);
TASK_PP(16'h1028E,4);
TASK_PP(16'h1028F,4);
TASK_PP(16'h10290,4);
TASK_PP(16'h10291,4);
TASK_PP(16'h10292,4);
TASK_PP(16'h10293,4);
TASK_PP(16'h10294,4);
TASK_PP(16'h10295,4);
TASK_PP(16'h10296,4);
TASK_PP(16'h10297,4);
TASK_PP(16'h10298,4);
TASK_PP(16'h10299,4);
TASK_PP(16'h1029A,4);
TASK_PP(16'h1029B,4);
TASK_PP(16'h1029C,4);
TASK_PP(16'h1029D,4);
TASK_PP(16'h1029E,4);
TASK_PP(16'h1029F,4);
TASK_PP(16'h102A0,4);
TASK_PP(16'h102A1,4);
TASK_PP(16'h102A2,4);
TASK_PP(16'h102A3,4);
TASK_PP(16'h102A4,4);
TASK_PP(16'h102A5,4);
TASK_PP(16'h102A6,4);
TASK_PP(16'h102A7,4);
TASK_PP(16'h102A8,4);
TASK_PP(16'h102A9,4);
TASK_PP(16'h102AA,4);
TASK_PP(16'h102AB,4);
TASK_PP(16'h102AC,4);
TASK_PP(16'h102AD,4);
TASK_PP(16'h102AE,4);
TASK_PP(16'h102AF,4);
TASK_PP(16'h102B0,4);
TASK_PP(16'h102B1,4);
TASK_PP(16'h102B2,4);
TASK_PP(16'h102B3,4);
TASK_PP(16'h102B4,4);
TASK_PP(16'h102B5,4);
TASK_PP(16'h102B6,4);
TASK_PP(16'h102B7,4);
TASK_PP(16'h102B8,4);
TASK_PP(16'h102B9,4);
TASK_PP(16'h102BA,4);
TASK_PP(16'h102BB,4);
TASK_PP(16'h102BC,4);
TASK_PP(16'h102BD,4);
TASK_PP(16'h102BE,4);
TASK_PP(16'h102BF,4);
TASK_PP(16'h102C0,4);
TASK_PP(16'h102C1,4);
TASK_PP(16'h102C2,4);
TASK_PP(16'h102C3,4);
TASK_PP(16'h102C4,4);
TASK_PP(16'h102C5,4);
TASK_PP(16'h102C6,4);
TASK_PP(16'h102C7,4);
TASK_PP(16'h102C8,4);
TASK_PP(16'h102C9,4);
TASK_PP(16'h102CA,4);
TASK_PP(16'h102CB,4);
TASK_PP(16'h102CC,4);
TASK_PP(16'h102CD,4);
TASK_PP(16'h102CE,4);
TASK_PP(16'h102CF,4);
TASK_PP(16'h102D0,4);
TASK_PP(16'h102D1,4);
TASK_PP(16'h102D2,4);
TASK_PP(16'h102D3,4);
TASK_PP(16'h102D4,4);
TASK_PP(16'h102D5,4);
TASK_PP(16'h102D6,4);
TASK_PP(16'h102D7,4);
TASK_PP(16'h102D8,4);
TASK_PP(16'h102D9,4);
TASK_PP(16'h102DA,4);
TASK_PP(16'h102DB,4);
TASK_PP(16'h102DC,4);
TASK_PP(16'h102DD,4);
TASK_PP(16'h102DE,4);
TASK_PP(16'h102DF,4);
TASK_PP(16'h102E0,4);
TASK_PP(16'h102E1,4);
TASK_PP(16'h102E2,4);
TASK_PP(16'h102E3,4);
TASK_PP(16'h102E4,4);
TASK_PP(16'h102E5,4);
TASK_PP(16'h102E6,4);
TASK_PP(16'h102E7,4);
TASK_PP(16'h102E8,4);
TASK_PP(16'h102E9,4);
TASK_PP(16'h102EA,4);
TASK_PP(16'h102EB,4);
TASK_PP(16'h102EC,4);
TASK_PP(16'h102ED,4);
TASK_PP(16'h102EE,4);
TASK_PP(16'h102EF,4);
TASK_PP(16'h102F0,4);
TASK_PP(16'h102F1,4);
TASK_PP(16'h102F2,4);
TASK_PP(16'h102F3,4);
TASK_PP(16'h102F4,4);
TASK_PP(16'h102F5,4);
TASK_PP(16'h102F6,4);
TASK_PP(16'h102F7,4);
TASK_PP(16'h102F8,4);
TASK_PP(16'h102F9,4);
TASK_PP(16'h102FA,4);
TASK_PP(16'h102FB,4);
TASK_PP(16'h102FC,4);
TASK_PP(16'h102FD,4);
TASK_PP(16'h102FE,4);
TASK_PP(16'h102FF,4);
TASK_PP(16'h10300,4);
TASK_PP(16'h10301,4);
TASK_PP(16'h10302,4);
TASK_PP(16'h10303,4);
TASK_PP(16'h10304,4);
TASK_PP(16'h10305,4);
TASK_PP(16'h10306,4);
TASK_PP(16'h10307,4);
TASK_PP(16'h10308,4);
TASK_PP(16'h10309,4);
TASK_PP(16'h1030A,4);
TASK_PP(16'h1030B,4);
TASK_PP(16'h1030C,4);
TASK_PP(16'h1030D,4);
TASK_PP(16'h1030E,4);
TASK_PP(16'h1030F,4);
TASK_PP(16'h10310,4);
TASK_PP(16'h10311,4);
TASK_PP(16'h10312,4);
TASK_PP(16'h10313,4);
TASK_PP(16'h10314,4);
TASK_PP(16'h10315,4);
TASK_PP(16'h10316,4);
TASK_PP(16'h10317,4);
TASK_PP(16'h10318,4);
TASK_PP(16'h10319,4);
TASK_PP(16'h1031A,4);
TASK_PP(16'h1031B,4);
TASK_PP(16'h1031C,4);
TASK_PP(16'h1031D,4);
TASK_PP(16'h1031E,4);
TASK_PP(16'h1031F,4);
TASK_PP(16'h10320,4);
TASK_PP(16'h10321,4);
TASK_PP(16'h10322,4);
TASK_PP(16'h10323,4);
TASK_PP(16'h10324,4);
TASK_PP(16'h10325,4);
TASK_PP(16'h10326,4);
TASK_PP(16'h10327,4);
TASK_PP(16'h10328,4);
TASK_PP(16'h10329,4);
TASK_PP(16'h1032A,4);
TASK_PP(16'h1032B,4);
TASK_PP(16'h1032C,4);
TASK_PP(16'h1032D,4);
TASK_PP(16'h1032E,4);
TASK_PP(16'h1032F,4);
TASK_PP(16'h10330,4);
TASK_PP(16'h10331,4);
TASK_PP(16'h10332,4);
TASK_PP(16'h10333,4);
TASK_PP(16'h10334,4);
TASK_PP(16'h10335,4);
TASK_PP(16'h10336,4);
TASK_PP(16'h10337,4);
TASK_PP(16'h10338,4);
TASK_PP(16'h10339,4);
TASK_PP(16'h1033A,4);
TASK_PP(16'h1033B,4);
TASK_PP(16'h1033C,4);
TASK_PP(16'h1033D,4);
TASK_PP(16'h1033E,4);
TASK_PP(16'h1033F,4);
TASK_PP(16'h10340,4);
TASK_PP(16'h10341,4);
TASK_PP(16'h10342,4);
TASK_PP(16'h10343,4);
TASK_PP(16'h10344,4);
TASK_PP(16'h10345,4);
TASK_PP(16'h10346,4);
TASK_PP(16'h10347,4);
TASK_PP(16'h10348,4);
TASK_PP(16'h10349,4);
TASK_PP(16'h1034A,4);
TASK_PP(16'h1034B,4);
TASK_PP(16'h1034C,4);
TASK_PP(16'h1034D,4);
TASK_PP(16'h1034E,4);
TASK_PP(16'h1034F,4);
TASK_PP(16'h10350,4);
TASK_PP(16'h10351,4);
TASK_PP(16'h10352,4);
TASK_PP(16'h10353,4);
TASK_PP(16'h10354,4);
TASK_PP(16'h10355,4);
TASK_PP(16'h10356,4);
TASK_PP(16'h10357,4);
TASK_PP(16'h10358,4);
TASK_PP(16'h10359,4);
TASK_PP(16'h1035A,4);
TASK_PP(16'h1035B,4);
TASK_PP(16'h1035C,4);
TASK_PP(16'h1035D,4);
TASK_PP(16'h1035E,4);
TASK_PP(16'h1035F,4);
TASK_PP(16'h10360,4);
TASK_PP(16'h10361,4);
TASK_PP(16'h10362,4);
TASK_PP(16'h10363,4);
TASK_PP(16'h10364,4);
TASK_PP(16'h10365,4);
TASK_PP(16'h10366,4);
TASK_PP(16'h10367,4);
TASK_PP(16'h10368,4);
TASK_PP(16'h10369,4);
TASK_PP(16'h1036A,4);
TASK_PP(16'h1036B,4);
TASK_PP(16'h1036C,4);
TASK_PP(16'h1036D,4);
TASK_PP(16'h1036E,4);
TASK_PP(16'h1036F,4);
TASK_PP(16'h10370,4);
TASK_PP(16'h10371,4);
TASK_PP(16'h10372,4);
TASK_PP(16'h10373,4);
TASK_PP(16'h10374,4);
TASK_PP(16'h10375,4);
TASK_PP(16'h10376,4);
TASK_PP(16'h10377,4);
TASK_PP(16'h10378,4);
TASK_PP(16'h10379,4);
TASK_PP(16'h1037A,4);
TASK_PP(16'h1037B,4);
TASK_PP(16'h1037C,4);
TASK_PP(16'h1037D,4);
TASK_PP(16'h1037E,4);
TASK_PP(16'h1037F,4);
TASK_PP(16'h10380,4);
TASK_PP(16'h10381,4);
TASK_PP(16'h10382,4);
TASK_PP(16'h10383,4);
TASK_PP(16'h10384,4);
TASK_PP(16'h10385,4);
TASK_PP(16'h10386,4);
TASK_PP(16'h10387,4);
TASK_PP(16'h10388,4);
TASK_PP(16'h10389,4);
TASK_PP(16'h1038A,4);
TASK_PP(16'h1038B,4);
TASK_PP(16'h1038C,4);
TASK_PP(16'h1038D,4);
TASK_PP(16'h1038E,4);
TASK_PP(16'h1038F,4);
TASK_PP(16'h10390,4);
TASK_PP(16'h10391,4);
TASK_PP(16'h10392,4);
TASK_PP(16'h10393,4);
TASK_PP(16'h10394,4);
TASK_PP(16'h10395,4);
TASK_PP(16'h10396,4);
TASK_PP(16'h10397,4);
TASK_PP(16'h10398,4);
TASK_PP(16'h10399,4);
TASK_PP(16'h1039A,4);
TASK_PP(16'h1039B,4);
TASK_PP(16'h1039C,4);
TASK_PP(16'h1039D,4);
TASK_PP(16'h1039E,4);
TASK_PP(16'h1039F,4);
TASK_PP(16'h103A0,4);
TASK_PP(16'h103A1,4);
TASK_PP(16'h103A2,4);
TASK_PP(16'h103A3,4);
TASK_PP(16'h103A4,4);
TASK_PP(16'h103A5,4);
TASK_PP(16'h103A6,4);
TASK_PP(16'h103A7,4);
TASK_PP(16'h103A8,4);
TASK_PP(16'h103A9,4);
TASK_PP(16'h103AA,4);
TASK_PP(16'h103AB,4);
TASK_PP(16'h103AC,4);
TASK_PP(16'h103AD,4);
TASK_PP(16'h103AE,4);
TASK_PP(16'h103AF,4);
TASK_PP(16'h103B0,4);
TASK_PP(16'h103B1,4);
TASK_PP(16'h103B2,4);
TASK_PP(16'h103B3,4);
TASK_PP(16'h103B4,4);
TASK_PP(16'h103B5,4);
TASK_PP(16'h103B6,4);
TASK_PP(16'h103B7,4);
TASK_PP(16'h103B8,4);
TASK_PP(16'h103B9,4);
TASK_PP(16'h103BA,4);
TASK_PP(16'h103BB,4);
TASK_PP(16'h103BC,4);
TASK_PP(16'h103BD,4);
TASK_PP(16'h103BE,4);
TASK_PP(16'h103BF,4);
TASK_PP(16'h103C0,4);
TASK_PP(16'h103C1,4);
TASK_PP(16'h103C2,4);
TASK_PP(16'h103C3,4);
TASK_PP(16'h103C4,4);
TASK_PP(16'h103C5,4);
TASK_PP(16'h103C6,4);
TASK_PP(16'h103C7,4);
TASK_PP(16'h103C8,4);
TASK_PP(16'h103C9,4);
TASK_PP(16'h103CA,4);
TASK_PP(16'h103CB,4);
TASK_PP(16'h103CC,4);
TASK_PP(16'h103CD,4);
TASK_PP(16'h103CE,4);
TASK_PP(16'h103CF,4);
TASK_PP(16'h103D0,4);
TASK_PP(16'h103D1,4);
TASK_PP(16'h103D2,4);
TASK_PP(16'h103D3,4);
TASK_PP(16'h103D4,4);
TASK_PP(16'h103D5,4);
TASK_PP(16'h103D6,4);
TASK_PP(16'h103D7,4);
TASK_PP(16'h103D8,4);
TASK_PP(16'h103D9,4);
TASK_PP(16'h103DA,4);
TASK_PP(16'h103DB,4);
TASK_PP(16'h103DC,4);
TASK_PP(16'h103DD,4);
TASK_PP(16'h103DE,4);
TASK_PP(16'h103DF,4);
TASK_PP(16'h103E0,4);
TASK_PP(16'h103E1,4);
TASK_PP(16'h103E2,4);
TASK_PP(16'h103E3,4);
TASK_PP(16'h103E4,4);
TASK_PP(16'h103E5,4);
TASK_PP(16'h103E6,4);
TASK_PP(16'h103E7,4);
TASK_PP(16'h103E8,4);
TASK_PP(16'h103E9,4);
TASK_PP(16'h103EA,4);
TASK_PP(16'h103EB,4);
TASK_PP(16'h103EC,4);
TASK_PP(16'h103ED,4);
TASK_PP(16'h103EE,4);
TASK_PP(16'h103EF,4);
TASK_PP(16'h103F0,4);
TASK_PP(16'h103F1,4);
TASK_PP(16'h103F2,4);
TASK_PP(16'h103F3,4);
TASK_PP(16'h103F4,4);
TASK_PP(16'h103F5,4);
TASK_PP(16'h103F6,4);
TASK_PP(16'h103F7,4);
TASK_PP(16'h103F8,4);
TASK_PP(16'h103F9,4);
TASK_PP(16'h103FA,4);
TASK_PP(16'h103FB,4);
TASK_PP(16'h103FC,4);
TASK_PP(16'h103FD,4);
TASK_PP(16'h103FE,4);
TASK_PP(16'h103FF,4);
TASK_PP(16'h10400,4);
TASK_PP(16'h10401,4);
TASK_PP(16'h10402,4);
TASK_PP(16'h10403,4);
TASK_PP(16'h10404,4);
TASK_PP(16'h10405,4);
TASK_PP(16'h10406,4);
TASK_PP(16'h10407,4);
TASK_PP(16'h10408,4);
TASK_PP(16'h10409,4);
TASK_PP(16'h1040A,4);
TASK_PP(16'h1040B,4);
TASK_PP(16'h1040C,4);
TASK_PP(16'h1040D,4);
TASK_PP(16'h1040E,4);
TASK_PP(16'h1040F,4);
TASK_PP(16'h10410,4);
TASK_PP(16'h10411,4);
TASK_PP(16'h10412,4);
TASK_PP(16'h10413,4);
TASK_PP(16'h10414,4);
TASK_PP(16'h10415,4);
TASK_PP(16'h10416,4);
TASK_PP(16'h10417,4);
TASK_PP(16'h10418,4);
TASK_PP(16'h10419,4);
TASK_PP(16'h1041A,4);
TASK_PP(16'h1041B,4);
TASK_PP(16'h1041C,4);
TASK_PP(16'h1041D,4);
TASK_PP(16'h1041E,4);
TASK_PP(16'h1041F,4);
TASK_PP(16'h10420,4);
TASK_PP(16'h10421,4);
TASK_PP(16'h10422,4);
TASK_PP(16'h10423,4);
TASK_PP(16'h10424,4);
TASK_PP(16'h10425,4);
TASK_PP(16'h10426,4);
TASK_PP(16'h10427,4);
TASK_PP(16'h10428,4);
TASK_PP(16'h10429,4);
TASK_PP(16'h1042A,4);
TASK_PP(16'h1042B,4);
TASK_PP(16'h1042C,4);
TASK_PP(16'h1042D,4);
TASK_PP(16'h1042E,4);
TASK_PP(16'h1042F,4);
TASK_PP(16'h10430,4);
TASK_PP(16'h10431,4);
TASK_PP(16'h10432,4);
TASK_PP(16'h10433,4);
TASK_PP(16'h10434,4);
TASK_PP(16'h10435,4);
TASK_PP(16'h10436,4);
TASK_PP(16'h10437,4);
TASK_PP(16'h10438,4);
TASK_PP(16'h10439,4);
TASK_PP(16'h1043A,4);
TASK_PP(16'h1043B,4);
TASK_PP(16'h1043C,4);
TASK_PP(16'h1043D,4);
TASK_PP(16'h1043E,4);
TASK_PP(16'h1043F,4);
TASK_PP(16'h10440,4);
TASK_PP(16'h10441,4);
TASK_PP(16'h10442,4);
TASK_PP(16'h10443,4);
TASK_PP(16'h10444,4);
TASK_PP(16'h10445,4);
TASK_PP(16'h10446,4);
TASK_PP(16'h10447,4);
TASK_PP(16'h10448,4);
TASK_PP(16'h10449,4);
TASK_PP(16'h1044A,4);
TASK_PP(16'h1044B,4);
TASK_PP(16'h1044C,4);
TASK_PP(16'h1044D,4);
TASK_PP(16'h1044E,4);
TASK_PP(16'h1044F,4);
TASK_PP(16'h10450,4);
TASK_PP(16'h10451,4);
TASK_PP(16'h10452,4);
TASK_PP(16'h10453,4);
TASK_PP(16'h10454,4);
TASK_PP(16'h10455,4);
TASK_PP(16'h10456,4);
TASK_PP(16'h10457,4);
TASK_PP(16'h10458,4);
TASK_PP(16'h10459,4);
TASK_PP(16'h1045A,4);
TASK_PP(16'h1045B,4);
TASK_PP(16'h1045C,4);
TASK_PP(16'h1045D,4);
TASK_PP(16'h1045E,4);
TASK_PP(16'h1045F,4);
TASK_PP(16'h10460,4);
TASK_PP(16'h10461,4);
TASK_PP(16'h10462,4);
TASK_PP(16'h10463,4);
TASK_PP(16'h10464,4);
TASK_PP(16'h10465,4);
TASK_PP(16'h10466,4);
TASK_PP(16'h10467,4);
TASK_PP(16'h10468,4);
TASK_PP(16'h10469,4);
TASK_PP(16'h1046A,4);
TASK_PP(16'h1046B,4);
TASK_PP(16'h1046C,4);
TASK_PP(16'h1046D,4);
TASK_PP(16'h1046E,4);
TASK_PP(16'h1046F,4);
TASK_PP(16'h10470,4);
TASK_PP(16'h10471,4);
TASK_PP(16'h10472,4);
TASK_PP(16'h10473,4);
TASK_PP(16'h10474,4);
TASK_PP(16'h10475,4);
TASK_PP(16'h10476,4);
TASK_PP(16'h10477,4);
TASK_PP(16'h10478,4);
TASK_PP(16'h10479,4);
TASK_PP(16'h1047A,4);
TASK_PP(16'h1047B,4);
TASK_PP(16'h1047C,4);
TASK_PP(16'h1047D,4);
TASK_PP(16'h1047E,4);
TASK_PP(16'h1047F,4);
TASK_PP(16'h10480,4);
TASK_PP(16'h10481,4);
TASK_PP(16'h10482,4);
TASK_PP(16'h10483,4);
TASK_PP(16'h10484,4);
TASK_PP(16'h10485,4);
TASK_PP(16'h10486,4);
TASK_PP(16'h10487,4);
TASK_PP(16'h10488,4);
TASK_PP(16'h10489,4);
TASK_PP(16'h1048A,4);
TASK_PP(16'h1048B,4);
TASK_PP(16'h1048C,4);
TASK_PP(16'h1048D,4);
TASK_PP(16'h1048E,4);
TASK_PP(16'h1048F,4);
TASK_PP(16'h10490,4);
TASK_PP(16'h10491,4);
TASK_PP(16'h10492,4);
TASK_PP(16'h10493,4);
TASK_PP(16'h10494,4);
TASK_PP(16'h10495,4);
TASK_PP(16'h10496,4);
TASK_PP(16'h10497,4);
TASK_PP(16'h10498,4);
TASK_PP(16'h10499,4);
TASK_PP(16'h1049A,4);
TASK_PP(16'h1049B,4);
TASK_PP(16'h1049C,4);
TASK_PP(16'h1049D,4);
TASK_PP(16'h1049E,4);
TASK_PP(16'h1049F,4);
TASK_PP(16'h104A0,4);
TASK_PP(16'h104A1,4);
TASK_PP(16'h104A2,4);
TASK_PP(16'h104A3,4);
TASK_PP(16'h104A4,4);
TASK_PP(16'h104A5,4);
TASK_PP(16'h104A6,4);
TASK_PP(16'h104A7,4);
TASK_PP(16'h104A8,4);
TASK_PP(16'h104A9,4);
TASK_PP(16'h104AA,4);
TASK_PP(16'h104AB,4);
TASK_PP(16'h104AC,4);
TASK_PP(16'h104AD,4);
TASK_PP(16'h104AE,4);
TASK_PP(16'h104AF,4);
TASK_PP(16'h104B0,4);
TASK_PP(16'h104B1,4);
TASK_PP(16'h104B2,4);
TASK_PP(16'h104B3,4);
TASK_PP(16'h104B4,4);
TASK_PP(16'h104B5,4);
TASK_PP(16'h104B6,4);
TASK_PP(16'h104B7,4);
TASK_PP(16'h104B8,4);
TASK_PP(16'h104B9,4);
TASK_PP(16'h104BA,4);
TASK_PP(16'h104BB,4);
TASK_PP(16'h104BC,4);
TASK_PP(16'h104BD,4);
TASK_PP(16'h104BE,4);
TASK_PP(16'h104BF,4);
TASK_PP(16'h104C0,4);
TASK_PP(16'h104C1,4);
TASK_PP(16'h104C2,4);
TASK_PP(16'h104C3,4);
TASK_PP(16'h104C4,4);
TASK_PP(16'h104C5,4);
TASK_PP(16'h104C6,4);
TASK_PP(16'h104C7,4);
TASK_PP(16'h104C8,4);
TASK_PP(16'h104C9,4);
TASK_PP(16'h104CA,4);
TASK_PP(16'h104CB,4);
TASK_PP(16'h104CC,4);
TASK_PP(16'h104CD,4);
TASK_PP(16'h104CE,4);
TASK_PP(16'h104CF,4);
TASK_PP(16'h104D0,4);
TASK_PP(16'h104D1,4);
TASK_PP(16'h104D2,4);
TASK_PP(16'h104D3,4);
TASK_PP(16'h104D4,4);
TASK_PP(16'h104D5,4);
TASK_PP(16'h104D6,4);
TASK_PP(16'h104D7,4);
TASK_PP(16'h104D8,4);
TASK_PP(16'h104D9,4);
TASK_PP(16'h104DA,4);
TASK_PP(16'h104DB,4);
TASK_PP(16'h104DC,4);
TASK_PP(16'h104DD,4);
TASK_PP(16'h104DE,4);
TASK_PP(16'h104DF,4);
TASK_PP(16'h104E0,4);
TASK_PP(16'h104E1,4);
TASK_PP(16'h104E2,4);
TASK_PP(16'h104E3,4);
TASK_PP(16'h104E4,4);
TASK_PP(16'h104E5,4);
TASK_PP(16'h104E6,4);
TASK_PP(16'h104E7,4);
TASK_PP(16'h104E8,4);
TASK_PP(16'h104E9,4);
TASK_PP(16'h104EA,4);
TASK_PP(16'h104EB,4);
TASK_PP(16'h104EC,4);
TASK_PP(16'h104ED,4);
TASK_PP(16'h104EE,4);
TASK_PP(16'h104EF,4);
TASK_PP(16'h104F0,4);
TASK_PP(16'h104F1,4);
TASK_PP(16'h104F2,4);
TASK_PP(16'h104F3,4);
TASK_PP(16'h104F4,4);
TASK_PP(16'h104F5,4);
TASK_PP(16'h104F6,4);
TASK_PP(16'h104F7,4);
TASK_PP(16'h104F8,4);
TASK_PP(16'h104F9,4);
TASK_PP(16'h104FA,4);
TASK_PP(16'h104FB,4);
TASK_PP(16'h104FC,4);
TASK_PP(16'h104FD,4);
TASK_PP(16'h104FE,4);
TASK_PP(16'h104FF,4);
TASK_PP(16'h10500,4);
TASK_PP(16'h10501,4);
TASK_PP(16'h10502,4);
TASK_PP(16'h10503,4);
TASK_PP(16'h10504,4);
TASK_PP(16'h10505,4);
TASK_PP(16'h10506,4);
TASK_PP(16'h10507,4);
TASK_PP(16'h10508,4);
TASK_PP(16'h10509,4);
TASK_PP(16'h1050A,4);
TASK_PP(16'h1050B,4);
TASK_PP(16'h1050C,4);
TASK_PP(16'h1050D,4);
TASK_PP(16'h1050E,4);
TASK_PP(16'h1050F,4);
TASK_PP(16'h10510,4);
TASK_PP(16'h10511,4);
TASK_PP(16'h10512,4);
TASK_PP(16'h10513,4);
TASK_PP(16'h10514,4);
TASK_PP(16'h10515,4);
TASK_PP(16'h10516,4);
TASK_PP(16'h10517,4);
TASK_PP(16'h10518,4);
TASK_PP(16'h10519,4);
TASK_PP(16'h1051A,4);
TASK_PP(16'h1051B,4);
TASK_PP(16'h1051C,4);
TASK_PP(16'h1051D,4);
TASK_PP(16'h1051E,4);
TASK_PP(16'h1051F,4);
TASK_PP(16'h10520,4);
TASK_PP(16'h10521,4);
TASK_PP(16'h10522,4);
TASK_PP(16'h10523,4);
TASK_PP(16'h10524,4);
TASK_PP(16'h10525,4);
TASK_PP(16'h10526,4);
TASK_PP(16'h10527,4);
TASK_PP(16'h10528,4);
TASK_PP(16'h10529,4);
TASK_PP(16'h1052A,4);
TASK_PP(16'h1052B,4);
TASK_PP(16'h1052C,4);
TASK_PP(16'h1052D,4);
TASK_PP(16'h1052E,4);
TASK_PP(16'h1052F,4);
TASK_PP(16'h10530,4);
TASK_PP(16'h10531,4);
TASK_PP(16'h10532,4);
TASK_PP(16'h10533,4);
TASK_PP(16'h10534,4);
TASK_PP(16'h10535,4);
TASK_PP(16'h10536,4);
TASK_PP(16'h10537,4);
TASK_PP(16'h10538,4);
TASK_PP(16'h10539,4);
TASK_PP(16'h1053A,4);
TASK_PP(16'h1053B,4);
TASK_PP(16'h1053C,4);
TASK_PP(16'h1053D,4);
TASK_PP(16'h1053E,4);
TASK_PP(16'h1053F,4);
TASK_PP(16'h10540,4);
TASK_PP(16'h10541,4);
TASK_PP(16'h10542,4);
TASK_PP(16'h10543,4);
TASK_PP(16'h10544,4);
TASK_PP(16'h10545,4);
TASK_PP(16'h10546,4);
TASK_PP(16'h10547,4);
TASK_PP(16'h10548,4);
TASK_PP(16'h10549,4);
TASK_PP(16'h1054A,4);
TASK_PP(16'h1054B,4);
TASK_PP(16'h1054C,4);
TASK_PP(16'h1054D,4);
TASK_PP(16'h1054E,4);
TASK_PP(16'h1054F,4);
TASK_PP(16'h10550,4);
TASK_PP(16'h10551,4);
TASK_PP(16'h10552,4);
TASK_PP(16'h10553,4);
TASK_PP(16'h10554,4);
TASK_PP(16'h10555,4);
TASK_PP(16'h10556,4);
TASK_PP(16'h10557,4);
TASK_PP(16'h10558,4);
TASK_PP(16'h10559,4);
TASK_PP(16'h1055A,4);
TASK_PP(16'h1055B,4);
TASK_PP(16'h1055C,4);
TASK_PP(16'h1055D,4);
TASK_PP(16'h1055E,4);
TASK_PP(16'h1055F,4);
TASK_PP(16'h10560,4);
TASK_PP(16'h10561,4);
TASK_PP(16'h10562,4);
TASK_PP(16'h10563,4);
TASK_PP(16'h10564,4);
TASK_PP(16'h10565,4);
TASK_PP(16'h10566,4);
TASK_PP(16'h10567,4);
TASK_PP(16'h10568,4);
TASK_PP(16'h10569,4);
TASK_PP(16'h1056A,4);
TASK_PP(16'h1056B,4);
TASK_PP(16'h1056C,4);
TASK_PP(16'h1056D,4);
TASK_PP(16'h1056E,4);
TASK_PP(16'h1056F,4);
TASK_PP(16'h10570,4);
TASK_PP(16'h10571,4);
TASK_PP(16'h10572,4);
TASK_PP(16'h10573,4);
TASK_PP(16'h10574,4);
TASK_PP(16'h10575,4);
TASK_PP(16'h10576,4);
TASK_PP(16'h10577,4);
TASK_PP(16'h10578,4);
TASK_PP(16'h10579,4);
TASK_PP(16'h1057A,4);
TASK_PP(16'h1057B,4);
TASK_PP(16'h1057C,4);
TASK_PP(16'h1057D,4);
TASK_PP(16'h1057E,4);
TASK_PP(16'h1057F,4);
TASK_PP(16'h10580,4);
TASK_PP(16'h10581,4);
TASK_PP(16'h10582,4);
TASK_PP(16'h10583,4);
TASK_PP(16'h10584,4);
TASK_PP(16'h10585,4);
TASK_PP(16'h10586,4);
TASK_PP(16'h10587,4);
TASK_PP(16'h10588,4);
TASK_PP(16'h10589,4);
TASK_PP(16'h1058A,4);
TASK_PP(16'h1058B,4);
TASK_PP(16'h1058C,4);
TASK_PP(16'h1058D,4);
TASK_PP(16'h1058E,4);
TASK_PP(16'h1058F,4);
TASK_PP(16'h10590,4);
TASK_PP(16'h10591,4);
TASK_PP(16'h10592,4);
TASK_PP(16'h10593,4);
TASK_PP(16'h10594,4);
TASK_PP(16'h10595,4);
TASK_PP(16'h10596,4);
TASK_PP(16'h10597,4);
TASK_PP(16'h10598,4);
TASK_PP(16'h10599,4);
TASK_PP(16'h1059A,4);
TASK_PP(16'h1059B,4);
TASK_PP(16'h1059C,4);
TASK_PP(16'h1059D,4);
TASK_PP(16'h1059E,4);
TASK_PP(16'h1059F,4);
TASK_PP(16'h105A0,4);
TASK_PP(16'h105A1,4);
TASK_PP(16'h105A2,4);
TASK_PP(16'h105A3,4);
TASK_PP(16'h105A4,4);
TASK_PP(16'h105A5,4);
TASK_PP(16'h105A6,4);
TASK_PP(16'h105A7,4);
TASK_PP(16'h105A8,4);
TASK_PP(16'h105A9,4);
TASK_PP(16'h105AA,4);
TASK_PP(16'h105AB,4);
TASK_PP(16'h105AC,4);
TASK_PP(16'h105AD,4);
TASK_PP(16'h105AE,4);
TASK_PP(16'h105AF,4);
TASK_PP(16'h105B0,4);
TASK_PP(16'h105B1,4);
TASK_PP(16'h105B2,4);
TASK_PP(16'h105B3,4);
TASK_PP(16'h105B4,4);
TASK_PP(16'h105B5,4);
TASK_PP(16'h105B6,4);
TASK_PP(16'h105B7,4);
TASK_PP(16'h105B8,4);
TASK_PP(16'h105B9,4);
TASK_PP(16'h105BA,4);
TASK_PP(16'h105BB,4);
TASK_PP(16'h105BC,4);
TASK_PP(16'h105BD,4);
TASK_PP(16'h105BE,4);
TASK_PP(16'h105BF,4);
TASK_PP(16'h105C0,4);
TASK_PP(16'h105C1,4);
TASK_PP(16'h105C2,4);
TASK_PP(16'h105C3,4);
TASK_PP(16'h105C4,4);
TASK_PP(16'h105C5,4);
TASK_PP(16'h105C6,4);
TASK_PP(16'h105C7,4);
TASK_PP(16'h105C8,4);
TASK_PP(16'h105C9,4);
TASK_PP(16'h105CA,4);
TASK_PP(16'h105CB,4);
TASK_PP(16'h105CC,4);
TASK_PP(16'h105CD,4);
TASK_PP(16'h105CE,4);
TASK_PP(16'h105CF,4);
TASK_PP(16'h105D0,4);
TASK_PP(16'h105D1,4);
TASK_PP(16'h105D2,4);
TASK_PP(16'h105D3,4);
TASK_PP(16'h105D4,4);
TASK_PP(16'h105D5,4);
TASK_PP(16'h105D6,4);
TASK_PP(16'h105D7,4);
TASK_PP(16'h105D8,4);
TASK_PP(16'h105D9,4);
TASK_PP(16'h105DA,4);
TASK_PP(16'h105DB,4);
TASK_PP(16'h105DC,4);
TASK_PP(16'h105DD,4);
TASK_PP(16'h105DE,4);
TASK_PP(16'h105DF,4);
TASK_PP(16'h105E0,4);
TASK_PP(16'h105E1,4);
TASK_PP(16'h105E2,4);
TASK_PP(16'h105E3,4);
TASK_PP(16'h105E4,4);
TASK_PP(16'h105E5,4);
TASK_PP(16'h105E6,4);
TASK_PP(16'h105E7,4);
TASK_PP(16'h105E8,4);
TASK_PP(16'h105E9,4);
TASK_PP(16'h105EA,4);
TASK_PP(16'h105EB,4);
TASK_PP(16'h105EC,4);
TASK_PP(16'h105ED,4);
TASK_PP(16'h105EE,4);
TASK_PP(16'h105EF,4);
TASK_PP(16'h105F0,4);
TASK_PP(16'h105F1,4);
TASK_PP(16'h105F2,4);
TASK_PP(16'h105F3,4);
TASK_PP(16'h105F4,4);
TASK_PP(16'h105F5,4);
TASK_PP(16'h105F6,4);
TASK_PP(16'h105F7,4);
TASK_PP(16'h105F8,4);
TASK_PP(16'h105F9,4);
TASK_PP(16'h105FA,4);
TASK_PP(16'h105FB,4);
TASK_PP(16'h105FC,4);
TASK_PP(16'h105FD,4);
TASK_PP(16'h105FE,4);
TASK_PP(16'h105FF,4);
TASK_PP(16'h10600,4);
TASK_PP(16'h10601,4);
TASK_PP(16'h10602,4);
TASK_PP(16'h10603,4);
TASK_PP(16'h10604,4);
TASK_PP(16'h10605,4);
TASK_PP(16'h10606,4);
TASK_PP(16'h10607,4);
TASK_PP(16'h10608,4);
TASK_PP(16'h10609,4);
TASK_PP(16'h1060A,4);
TASK_PP(16'h1060B,4);
TASK_PP(16'h1060C,4);
TASK_PP(16'h1060D,4);
TASK_PP(16'h1060E,4);
TASK_PP(16'h1060F,4);
TASK_PP(16'h10610,4);
TASK_PP(16'h10611,4);
TASK_PP(16'h10612,4);
TASK_PP(16'h10613,4);
TASK_PP(16'h10614,4);
TASK_PP(16'h10615,4);
TASK_PP(16'h10616,4);
TASK_PP(16'h10617,4);
TASK_PP(16'h10618,4);
TASK_PP(16'h10619,4);
TASK_PP(16'h1061A,4);
TASK_PP(16'h1061B,4);
TASK_PP(16'h1061C,4);
TASK_PP(16'h1061D,4);
TASK_PP(16'h1061E,4);
TASK_PP(16'h1061F,4);
TASK_PP(16'h10620,4);
TASK_PP(16'h10621,4);
TASK_PP(16'h10622,4);
TASK_PP(16'h10623,4);
TASK_PP(16'h10624,4);
TASK_PP(16'h10625,4);
TASK_PP(16'h10626,4);
TASK_PP(16'h10627,4);
TASK_PP(16'h10628,4);
TASK_PP(16'h10629,4);
TASK_PP(16'h1062A,4);
TASK_PP(16'h1062B,4);
TASK_PP(16'h1062C,4);
TASK_PP(16'h1062D,4);
TASK_PP(16'h1062E,4);
TASK_PP(16'h1062F,4);
TASK_PP(16'h10630,4);
TASK_PP(16'h10631,4);
TASK_PP(16'h10632,4);
TASK_PP(16'h10633,4);
TASK_PP(16'h10634,4);
TASK_PP(16'h10635,4);
TASK_PP(16'h10636,4);
TASK_PP(16'h10637,4);
TASK_PP(16'h10638,4);
TASK_PP(16'h10639,4);
TASK_PP(16'h1063A,4);
TASK_PP(16'h1063B,4);
TASK_PP(16'h1063C,4);
TASK_PP(16'h1063D,4);
TASK_PP(16'h1063E,4);
TASK_PP(16'h1063F,4);
TASK_PP(16'h10640,4);
TASK_PP(16'h10641,4);
TASK_PP(16'h10642,4);
TASK_PP(16'h10643,4);
TASK_PP(16'h10644,4);
TASK_PP(16'h10645,4);
TASK_PP(16'h10646,4);
TASK_PP(16'h10647,4);
TASK_PP(16'h10648,4);
TASK_PP(16'h10649,4);
TASK_PP(16'h1064A,4);
TASK_PP(16'h1064B,4);
TASK_PP(16'h1064C,4);
TASK_PP(16'h1064D,4);
TASK_PP(16'h1064E,4);
TASK_PP(16'h1064F,4);
TASK_PP(16'h10650,4);
TASK_PP(16'h10651,4);
TASK_PP(16'h10652,4);
TASK_PP(16'h10653,4);
TASK_PP(16'h10654,4);
TASK_PP(16'h10655,4);
TASK_PP(16'h10656,4);
TASK_PP(16'h10657,4);
TASK_PP(16'h10658,4);
TASK_PP(16'h10659,4);
TASK_PP(16'h1065A,4);
TASK_PP(16'h1065B,4);
TASK_PP(16'h1065C,4);
TASK_PP(16'h1065D,4);
TASK_PP(16'h1065E,4);
TASK_PP(16'h1065F,4);
TASK_PP(16'h10660,4);
TASK_PP(16'h10661,4);
TASK_PP(16'h10662,4);
TASK_PP(16'h10663,4);
TASK_PP(16'h10664,4);
TASK_PP(16'h10665,4);
TASK_PP(16'h10666,4);
TASK_PP(16'h10667,4);
TASK_PP(16'h10668,4);
TASK_PP(16'h10669,4);
TASK_PP(16'h1066A,4);
TASK_PP(16'h1066B,4);
TASK_PP(16'h1066C,4);
TASK_PP(16'h1066D,4);
TASK_PP(16'h1066E,4);
TASK_PP(16'h1066F,4);
TASK_PP(16'h10670,4);
TASK_PP(16'h10671,4);
TASK_PP(16'h10672,4);
TASK_PP(16'h10673,4);
TASK_PP(16'h10674,4);
TASK_PP(16'h10675,4);
TASK_PP(16'h10676,4);
TASK_PP(16'h10677,4);
TASK_PP(16'h10678,4);
TASK_PP(16'h10679,4);
TASK_PP(16'h1067A,4);
TASK_PP(16'h1067B,4);
TASK_PP(16'h1067C,4);
TASK_PP(16'h1067D,4);
TASK_PP(16'h1067E,4);
TASK_PP(16'h1067F,4);
TASK_PP(16'h10680,4);
TASK_PP(16'h10681,4);
TASK_PP(16'h10682,4);
TASK_PP(16'h10683,4);
TASK_PP(16'h10684,4);
TASK_PP(16'h10685,4);
TASK_PP(16'h10686,4);
TASK_PP(16'h10687,4);
TASK_PP(16'h10688,4);
TASK_PP(16'h10689,4);
TASK_PP(16'h1068A,4);
TASK_PP(16'h1068B,4);
TASK_PP(16'h1068C,4);
TASK_PP(16'h1068D,4);
TASK_PP(16'h1068E,4);
TASK_PP(16'h1068F,4);
TASK_PP(16'h10690,4);
TASK_PP(16'h10691,4);
TASK_PP(16'h10692,4);
TASK_PP(16'h10693,4);
TASK_PP(16'h10694,4);
TASK_PP(16'h10695,4);
TASK_PP(16'h10696,4);
TASK_PP(16'h10697,4);
TASK_PP(16'h10698,4);
TASK_PP(16'h10699,4);
TASK_PP(16'h1069A,4);
TASK_PP(16'h1069B,4);
TASK_PP(16'h1069C,4);
TASK_PP(16'h1069D,4);
TASK_PP(16'h1069E,4);
TASK_PP(16'h1069F,4);
TASK_PP(16'h106A0,4);
TASK_PP(16'h106A1,4);
TASK_PP(16'h106A2,4);
TASK_PP(16'h106A3,4);
TASK_PP(16'h106A4,4);
TASK_PP(16'h106A5,4);
TASK_PP(16'h106A6,4);
TASK_PP(16'h106A7,4);
TASK_PP(16'h106A8,4);
TASK_PP(16'h106A9,4);
TASK_PP(16'h106AA,4);
TASK_PP(16'h106AB,4);
TASK_PP(16'h106AC,4);
TASK_PP(16'h106AD,4);
TASK_PP(16'h106AE,4);
TASK_PP(16'h106AF,4);
TASK_PP(16'h106B0,4);
TASK_PP(16'h106B1,4);
TASK_PP(16'h106B2,4);
TASK_PP(16'h106B3,4);
TASK_PP(16'h106B4,4);
TASK_PP(16'h106B5,4);
TASK_PP(16'h106B6,4);
TASK_PP(16'h106B7,4);
TASK_PP(16'h106B8,4);
TASK_PP(16'h106B9,4);
TASK_PP(16'h106BA,4);
TASK_PP(16'h106BB,4);
TASK_PP(16'h106BC,4);
TASK_PP(16'h106BD,4);
TASK_PP(16'h106BE,4);
TASK_PP(16'h106BF,4);
TASK_PP(16'h106C0,4);
TASK_PP(16'h106C1,4);
TASK_PP(16'h106C2,4);
TASK_PP(16'h106C3,4);
TASK_PP(16'h106C4,4);
TASK_PP(16'h106C5,4);
TASK_PP(16'h106C6,4);
TASK_PP(16'h106C7,4);
TASK_PP(16'h106C8,4);
TASK_PP(16'h106C9,4);
TASK_PP(16'h106CA,4);
TASK_PP(16'h106CB,4);
TASK_PP(16'h106CC,4);
TASK_PP(16'h106CD,4);
TASK_PP(16'h106CE,4);
TASK_PP(16'h106CF,4);
TASK_PP(16'h106D0,4);
TASK_PP(16'h106D1,4);
TASK_PP(16'h106D2,4);
TASK_PP(16'h106D3,4);
TASK_PP(16'h106D4,4);
TASK_PP(16'h106D5,4);
TASK_PP(16'h106D6,4);
TASK_PP(16'h106D7,4);
TASK_PP(16'h106D8,4);
TASK_PP(16'h106D9,4);
TASK_PP(16'h106DA,4);
TASK_PP(16'h106DB,4);
TASK_PP(16'h106DC,4);
TASK_PP(16'h106DD,4);
TASK_PP(16'h106DE,4);
TASK_PP(16'h106DF,4);
TASK_PP(16'h106E0,4);
TASK_PP(16'h106E1,4);
TASK_PP(16'h106E2,4);
TASK_PP(16'h106E3,4);
TASK_PP(16'h106E4,4);
TASK_PP(16'h106E5,4);
TASK_PP(16'h106E6,4);
TASK_PP(16'h106E7,4);
TASK_PP(16'h106E8,4);
TASK_PP(16'h106E9,4);
TASK_PP(16'h106EA,4);
TASK_PP(16'h106EB,4);
TASK_PP(16'h106EC,4);
TASK_PP(16'h106ED,4);
TASK_PP(16'h106EE,4);
TASK_PP(16'h106EF,4);
TASK_PP(16'h106F0,4);
TASK_PP(16'h106F1,4);
TASK_PP(16'h106F2,4);
TASK_PP(16'h106F3,4);
TASK_PP(16'h106F4,4);
TASK_PP(16'h106F5,4);
TASK_PP(16'h106F6,4);
TASK_PP(16'h106F7,4);
TASK_PP(16'h106F8,4);
TASK_PP(16'h106F9,4);
TASK_PP(16'h106FA,4);
TASK_PP(16'h106FB,4);
TASK_PP(16'h106FC,4);
TASK_PP(16'h106FD,4);
TASK_PP(16'h106FE,4);
TASK_PP(16'h106FF,4);
TASK_PP(16'h10700,4);
TASK_PP(16'h10701,4);
TASK_PP(16'h10702,4);
TASK_PP(16'h10703,4);
TASK_PP(16'h10704,4);
TASK_PP(16'h10705,4);
TASK_PP(16'h10706,4);
TASK_PP(16'h10707,4);
TASK_PP(16'h10708,4);
TASK_PP(16'h10709,4);
TASK_PP(16'h1070A,4);
TASK_PP(16'h1070B,4);
TASK_PP(16'h1070C,4);
TASK_PP(16'h1070D,4);
TASK_PP(16'h1070E,4);
TASK_PP(16'h1070F,4);
TASK_PP(16'h10710,4);
TASK_PP(16'h10711,4);
TASK_PP(16'h10712,4);
TASK_PP(16'h10713,4);
TASK_PP(16'h10714,4);
TASK_PP(16'h10715,4);
TASK_PP(16'h10716,4);
TASK_PP(16'h10717,4);
TASK_PP(16'h10718,4);
TASK_PP(16'h10719,4);
TASK_PP(16'h1071A,4);
TASK_PP(16'h1071B,4);
TASK_PP(16'h1071C,4);
TASK_PP(16'h1071D,4);
TASK_PP(16'h1071E,4);
TASK_PP(16'h1071F,4);
TASK_PP(16'h10720,4);
TASK_PP(16'h10721,4);
TASK_PP(16'h10722,4);
TASK_PP(16'h10723,4);
TASK_PP(16'h10724,4);
TASK_PP(16'h10725,4);
TASK_PP(16'h10726,4);
TASK_PP(16'h10727,4);
TASK_PP(16'h10728,4);
TASK_PP(16'h10729,4);
TASK_PP(16'h1072A,4);
TASK_PP(16'h1072B,4);
TASK_PP(16'h1072C,4);
TASK_PP(16'h1072D,4);
TASK_PP(16'h1072E,4);
TASK_PP(16'h1072F,4);
TASK_PP(16'h10730,4);
TASK_PP(16'h10731,4);
TASK_PP(16'h10732,4);
TASK_PP(16'h10733,4);
TASK_PP(16'h10734,4);
TASK_PP(16'h10735,4);
TASK_PP(16'h10736,4);
TASK_PP(16'h10737,4);
TASK_PP(16'h10738,4);
TASK_PP(16'h10739,4);
TASK_PP(16'h1073A,4);
TASK_PP(16'h1073B,4);
TASK_PP(16'h1073C,4);
TASK_PP(16'h1073D,4);
TASK_PP(16'h1073E,4);
TASK_PP(16'h1073F,4);
TASK_PP(16'h10740,4);
TASK_PP(16'h10741,4);
TASK_PP(16'h10742,4);
TASK_PP(16'h10743,4);
TASK_PP(16'h10744,4);
TASK_PP(16'h10745,4);
TASK_PP(16'h10746,4);
TASK_PP(16'h10747,4);
TASK_PP(16'h10748,4);
TASK_PP(16'h10749,4);
TASK_PP(16'h1074A,4);
TASK_PP(16'h1074B,4);
TASK_PP(16'h1074C,4);
TASK_PP(16'h1074D,4);
TASK_PP(16'h1074E,4);
TASK_PP(16'h1074F,4);
TASK_PP(16'h10750,4);
TASK_PP(16'h10751,4);
TASK_PP(16'h10752,4);
TASK_PP(16'h10753,4);
TASK_PP(16'h10754,4);
TASK_PP(16'h10755,4);
TASK_PP(16'h10756,4);
TASK_PP(16'h10757,4);
TASK_PP(16'h10758,4);
TASK_PP(16'h10759,4);
TASK_PP(16'h1075A,4);
TASK_PP(16'h1075B,4);
TASK_PP(16'h1075C,4);
TASK_PP(16'h1075D,4);
TASK_PP(16'h1075E,4);
TASK_PP(16'h1075F,4);
TASK_PP(16'h10760,4);
TASK_PP(16'h10761,4);
TASK_PP(16'h10762,4);
TASK_PP(16'h10763,4);
TASK_PP(16'h10764,4);
TASK_PP(16'h10765,4);
TASK_PP(16'h10766,4);
TASK_PP(16'h10767,4);
TASK_PP(16'h10768,4);
TASK_PP(16'h10769,4);
TASK_PP(16'h1076A,4);
TASK_PP(16'h1076B,4);
TASK_PP(16'h1076C,4);
TASK_PP(16'h1076D,4);
TASK_PP(16'h1076E,4);
TASK_PP(16'h1076F,4);
TASK_PP(16'h10770,4);
TASK_PP(16'h10771,4);
TASK_PP(16'h10772,4);
TASK_PP(16'h10773,4);
TASK_PP(16'h10774,4);
TASK_PP(16'h10775,4);
TASK_PP(16'h10776,4);
TASK_PP(16'h10777,4);
TASK_PP(16'h10778,4);
TASK_PP(16'h10779,4);
TASK_PP(16'h1077A,4);
TASK_PP(16'h1077B,4);
TASK_PP(16'h1077C,4);
TASK_PP(16'h1077D,4);
TASK_PP(16'h1077E,4);
TASK_PP(16'h1077F,4);
TASK_PP(16'h10780,4);
TASK_PP(16'h10781,4);
TASK_PP(16'h10782,4);
TASK_PP(16'h10783,4);
TASK_PP(16'h10784,4);
TASK_PP(16'h10785,4);
TASK_PP(16'h10786,4);
TASK_PP(16'h10787,4);
TASK_PP(16'h10788,4);
TASK_PP(16'h10789,4);
TASK_PP(16'h1078A,4);
TASK_PP(16'h1078B,4);
TASK_PP(16'h1078C,4);
TASK_PP(16'h1078D,4);
TASK_PP(16'h1078E,4);
TASK_PP(16'h1078F,4);
TASK_PP(16'h10790,4);
TASK_PP(16'h10791,4);
TASK_PP(16'h10792,4);
TASK_PP(16'h10793,4);
TASK_PP(16'h10794,4);
TASK_PP(16'h10795,4);
TASK_PP(16'h10796,4);
TASK_PP(16'h10797,4);
TASK_PP(16'h10798,4);
TASK_PP(16'h10799,4);
TASK_PP(16'h1079A,4);
TASK_PP(16'h1079B,4);
TASK_PP(16'h1079C,4);
TASK_PP(16'h1079D,4);
TASK_PP(16'h1079E,4);
TASK_PP(16'h1079F,4);
TASK_PP(16'h107A0,4);
TASK_PP(16'h107A1,4);
TASK_PP(16'h107A2,4);
TASK_PP(16'h107A3,4);
TASK_PP(16'h107A4,4);
TASK_PP(16'h107A5,4);
TASK_PP(16'h107A6,4);
TASK_PP(16'h107A7,4);
TASK_PP(16'h107A8,4);
TASK_PP(16'h107A9,4);
TASK_PP(16'h107AA,4);
TASK_PP(16'h107AB,4);
TASK_PP(16'h107AC,4);
TASK_PP(16'h107AD,4);
TASK_PP(16'h107AE,4);
TASK_PP(16'h107AF,4);
TASK_PP(16'h107B0,4);
TASK_PP(16'h107B1,4);
TASK_PP(16'h107B2,4);
TASK_PP(16'h107B3,4);
TASK_PP(16'h107B4,4);
TASK_PP(16'h107B5,4);
TASK_PP(16'h107B6,4);
TASK_PP(16'h107B7,4);
TASK_PP(16'h107B8,4);
TASK_PP(16'h107B9,4);
TASK_PP(16'h107BA,4);
TASK_PP(16'h107BB,4);
TASK_PP(16'h107BC,4);
TASK_PP(16'h107BD,4);
TASK_PP(16'h107BE,4);
TASK_PP(16'h107BF,4);
TASK_PP(16'h107C0,4);
TASK_PP(16'h107C1,4);
TASK_PP(16'h107C2,4);
TASK_PP(16'h107C3,4);
TASK_PP(16'h107C4,4);
TASK_PP(16'h107C5,4);
TASK_PP(16'h107C6,4);
TASK_PP(16'h107C7,4);
TASK_PP(16'h107C8,4);
TASK_PP(16'h107C9,4);
TASK_PP(16'h107CA,4);
TASK_PP(16'h107CB,4);
TASK_PP(16'h107CC,4);
TASK_PP(16'h107CD,4);
TASK_PP(16'h107CE,4);
TASK_PP(16'h107CF,4);
TASK_PP(16'h107D0,4);
TASK_PP(16'h107D1,4);
TASK_PP(16'h107D2,4);
TASK_PP(16'h107D3,4);
TASK_PP(16'h107D4,4);
TASK_PP(16'h107D5,4);
TASK_PP(16'h107D6,4);
TASK_PP(16'h107D7,4);
TASK_PP(16'h107D8,4);
TASK_PP(16'h107D9,4);
TASK_PP(16'h107DA,4);
TASK_PP(16'h107DB,4);
TASK_PP(16'h107DC,4);
TASK_PP(16'h107DD,4);
TASK_PP(16'h107DE,4);
TASK_PP(16'h107DF,4);
TASK_PP(16'h107E0,4);
TASK_PP(16'h107E1,4);
TASK_PP(16'h107E2,4);
TASK_PP(16'h107E3,4);
TASK_PP(16'h107E4,4);
TASK_PP(16'h107E5,4);
TASK_PP(16'h107E6,4);
TASK_PP(16'h107E7,4);
TASK_PP(16'h107E8,4);
TASK_PP(16'h107E9,4);
TASK_PP(16'h107EA,4);
TASK_PP(16'h107EB,4);
TASK_PP(16'h107EC,4);
TASK_PP(16'h107ED,4);
TASK_PP(16'h107EE,4);
TASK_PP(16'h107EF,4);
TASK_PP(16'h107F0,4);
TASK_PP(16'h107F1,4);
TASK_PP(16'h107F2,4);
TASK_PP(16'h107F3,4);
TASK_PP(16'h107F4,4);
TASK_PP(16'h107F5,4);
TASK_PP(16'h107F6,4);
TASK_PP(16'h107F7,4);
TASK_PP(16'h107F8,4);
TASK_PP(16'h107F9,4);
TASK_PP(16'h107FA,4);
TASK_PP(16'h107FB,4);
TASK_PP(16'h107FC,4);
TASK_PP(16'h107FD,4);
TASK_PP(16'h107FE,4);
TASK_PP(16'h107FF,4);
TASK_PP(16'h10800,4);
TASK_PP(16'h10801,4);
TASK_PP(16'h10802,4);
TASK_PP(16'h10803,4);
TASK_PP(16'h10804,4);
TASK_PP(16'h10805,4);
TASK_PP(16'h10806,4);
TASK_PP(16'h10807,4);
TASK_PP(16'h10808,4);
TASK_PP(16'h10809,4);
TASK_PP(16'h1080A,4);
TASK_PP(16'h1080B,4);
TASK_PP(16'h1080C,4);
TASK_PP(16'h1080D,4);
TASK_PP(16'h1080E,4);
TASK_PP(16'h1080F,4);
TASK_PP(16'h10810,4);
TASK_PP(16'h10811,4);
TASK_PP(16'h10812,4);
TASK_PP(16'h10813,4);
TASK_PP(16'h10814,4);
TASK_PP(16'h10815,4);
TASK_PP(16'h10816,4);
TASK_PP(16'h10817,4);
TASK_PP(16'h10818,4);
TASK_PP(16'h10819,4);
TASK_PP(16'h1081A,4);
TASK_PP(16'h1081B,4);
TASK_PP(16'h1081C,4);
TASK_PP(16'h1081D,4);
TASK_PP(16'h1081E,4);
TASK_PP(16'h1081F,4);
TASK_PP(16'h10820,4);
TASK_PP(16'h10821,4);
TASK_PP(16'h10822,4);
TASK_PP(16'h10823,4);
TASK_PP(16'h10824,4);
TASK_PP(16'h10825,4);
TASK_PP(16'h10826,4);
TASK_PP(16'h10827,4);
TASK_PP(16'h10828,4);
TASK_PP(16'h10829,4);
TASK_PP(16'h1082A,4);
TASK_PP(16'h1082B,4);
TASK_PP(16'h1082C,4);
TASK_PP(16'h1082D,4);
TASK_PP(16'h1082E,4);
TASK_PP(16'h1082F,4);
TASK_PP(16'h10830,4);
TASK_PP(16'h10831,4);
TASK_PP(16'h10832,4);
TASK_PP(16'h10833,4);
TASK_PP(16'h10834,4);
TASK_PP(16'h10835,4);
TASK_PP(16'h10836,4);
TASK_PP(16'h10837,4);
TASK_PP(16'h10838,4);
TASK_PP(16'h10839,4);
TASK_PP(16'h1083A,4);
TASK_PP(16'h1083B,4);
TASK_PP(16'h1083C,4);
TASK_PP(16'h1083D,4);
TASK_PP(16'h1083E,4);
TASK_PP(16'h1083F,4);
TASK_PP(16'h10840,4);
TASK_PP(16'h10841,4);
TASK_PP(16'h10842,4);
TASK_PP(16'h10843,4);
TASK_PP(16'h10844,4);
TASK_PP(16'h10845,4);
TASK_PP(16'h10846,4);
TASK_PP(16'h10847,4);
TASK_PP(16'h10848,4);
TASK_PP(16'h10849,4);
TASK_PP(16'h1084A,4);
TASK_PP(16'h1084B,4);
TASK_PP(16'h1084C,4);
TASK_PP(16'h1084D,4);
TASK_PP(16'h1084E,4);
TASK_PP(16'h1084F,4);
TASK_PP(16'h10850,4);
TASK_PP(16'h10851,4);
TASK_PP(16'h10852,4);
TASK_PP(16'h10853,4);
TASK_PP(16'h10854,4);
TASK_PP(16'h10855,4);
TASK_PP(16'h10856,4);
TASK_PP(16'h10857,4);
TASK_PP(16'h10858,4);
TASK_PP(16'h10859,4);
TASK_PP(16'h1085A,4);
TASK_PP(16'h1085B,4);
TASK_PP(16'h1085C,4);
TASK_PP(16'h1085D,4);
TASK_PP(16'h1085E,4);
TASK_PP(16'h1085F,4);
TASK_PP(16'h10860,4);
TASK_PP(16'h10861,4);
TASK_PP(16'h10862,4);
TASK_PP(16'h10863,4);
TASK_PP(16'h10864,4);
TASK_PP(16'h10865,4);
TASK_PP(16'h10866,4);
TASK_PP(16'h10867,4);
TASK_PP(16'h10868,4);
TASK_PP(16'h10869,4);
TASK_PP(16'h1086A,4);
TASK_PP(16'h1086B,4);
TASK_PP(16'h1086C,4);
TASK_PP(16'h1086D,4);
TASK_PP(16'h1086E,4);
TASK_PP(16'h1086F,4);
TASK_PP(16'h10870,4);
TASK_PP(16'h10871,4);
TASK_PP(16'h10872,4);
TASK_PP(16'h10873,4);
TASK_PP(16'h10874,4);
TASK_PP(16'h10875,4);
TASK_PP(16'h10876,4);
TASK_PP(16'h10877,4);
TASK_PP(16'h10878,4);
TASK_PP(16'h10879,4);
TASK_PP(16'h1087A,4);
TASK_PP(16'h1087B,4);
TASK_PP(16'h1087C,4);
TASK_PP(16'h1087D,4);
TASK_PP(16'h1087E,4);
TASK_PP(16'h1087F,4);
TASK_PP(16'h10880,4);
TASK_PP(16'h10881,4);
TASK_PP(16'h10882,4);
TASK_PP(16'h10883,4);
TASK_PP(16'h10884,4);
TASK_PP(16'h10885,4);
TASK_PP(16'h10886,4);
TASK_PP(16'h10887,4);
TASK_PP(16'h10888,4);
TASK_PP(16'h10889,4);
TASK_PP(16'h1088A,4);
TASK_PP(16'h1088B,4);
TASK_PP(16'h1088C,4);
TASK_PP(16'h1088D,4);
TASK_PP(16'h1088E,4);
TASK_PP(16'h1088F,4);
TASK_PP(16'h10890,4);
TASK_PP(16'h10891,4);
TASK_PP(16'h10892,4);
TASK_PP(16'h10893,4);
TASK_PP(16'h10894,4);
TASK_PP(16'h10895,4);
TASK_PP(16'h10896,4);
TASK_PP(16'h10897,4);
TASK_PP(16'h10898,4);
TASK_PP(16'h10899,4);
TASK_PP(16'h1089A,4);
TASK_PP(16'h1089B,4);
TASK_PP(16'h1089C,4);
TASK_PP(16'h1089D,4);
TASK_PP(16'h1089E,4);
TASK_PP(16'h1089F,4);
TASK_PP(16'h108A0,4);
TASK_PP(16'h108A1,4);
TASK_PP(16'h108A2,4);
TASK_PP(16'h108A3,4);
TASK_PP(16'h108A4,4);
TASK_PP(16'h108A5,4);
TASK_PP(16'h108A6,4);
TASK_PP(16'h108A7,4);
TASK_PP(16'h108A8,4);
TASK_PP(16'h108A9,4);
TASK_PP(16'h108AA,4);
TASK_PP(16'h108AB,4);
TASK_PP(16'h108AC,4);
TASK_PP(16'h108AD,4);
TASK_PP(16'h108AE,4);
TASK_PP(16'h108AF,4);
TASK_PP(16'h108B0,4);
TASK_PP(16'h108B1,4);
TASK_PP(16'h108B2,4);
TASK_PP(16'h108B3,4);
TASK_PP(16'h108B4,4);
TASK_PP(16'h108B5,4);
TASK_PP(16'h108B6,4);
TASK_PP(16'h108B7,4);
TASK_PP(16'h108B8,4);
TASK_PP(16'h108B9,4);
TASK_PP(16'h108BA,4);
TASK_PP(16'h108BB,4);
TASK_PP(16'h108BC,4);
TASK_PP(16'h108BD,4);
TASK_PP(16'h108BE,4);
TASK_PP(16'h108BF,4);
TASK_PP(16'h108C0,4);
TASK_PP(16'h108C1,4);
TASK_PP(16'h108C2,4);
TASK_PP(16'h108C3,4);
TASK_PP(16'h108C4,4);
TASK_PP(16'h108C5,4);
TASK_PP(16'h108C6,4);
TASK_PP(16'h108C7,4);
TASK_PP(16'h108C8,4);
TASK_PP(16'h108C9,4);
TASK_PP(16'h108CA,4);
TASK_PP(16'h108CB,4);
TASK_PP(16'h108CC,4);
TASK_PP(16'h108CD,4);
TASK_PP(16'h108CE,4);
TASK_PP(16'h108CF,4);
TASK_PP(16'h108D0,4);
TASK_PP(16'h108D1,4);
TASK_PP(16'h108D2,4);
TASK_PP(16'h108D3,4);
TASK_PP(16'h108D4,4);
TASK_PP(16'h108D5,4);
TASK_PP(16'h108D6,4);
TASK_PP(16'h108D7,4);
TASK_PP(16'h108D8,4);
TASK_PP(16'h108D9,4);
TASK_PP(16'h108DA,4);
TASK_PP(16'h108DB,4);
TASK_PP(16'h108DC,4);
TASK_PP(16'h108DD,4);
TASK_PP(16'h108DE,4);
TASK_PP(16'h108DF,4);
TASK_PP(16'h108E0,4);
TASK_PP(16'h108E1,4);
TASK_PP(16'h108E2,4);
TASK_PP(16'h108E3,4);
TASK_PP(16'h108E4,4);
TASK_PP(16'h108E5,4);
TASK_PP(16'h108E6,4);
TASK_PP(16'h108E7,4);
TASK_PP(16'h108E8,4);
TASK_PP(16'h108E9,4);
TASK_PP(16'h108EA,4);
TASK_PP(16'h108EB,4);
TASK_PP(16'h108EC,4);
TASK_PP(16'h108ED,4);
TASK_PP(16'h108EE,4);
TASK_PP(16'h108EF,4);
TASK_PP(16'h108F0,4);
TASK_PP(16'h108F1,4);
TASK_PP(16'h108F2,4);
TASK_PP(16'h108F3,4);
TASK_PP(16'h108F4,4);
TASK_PP(16'h108F5,4);
TASK_PP(16'h108F6,4);
TASK_PP(16'h108F7,4);
TASK_PP(16'h108F8,4);
TASK_PP(16'h108F9,4);
TASK_PP(16'h108FA,4);
TASK_PP(16'h108FB,4);
TASK_PP(16'h108FC,4);
TASK_PP(16'h108FD,4);
TASK_PP(16'h108FE,4);
TASK_PP(16'h108FF,4);
TASK_PP(16'h10900,4);
TASK_PP(16'h10901,4);
TASK_PP(16'h10902,4);
TASK_PP(16'h10903,4);
TASK_PP(16'h10904,4);
TASK_PP(16'h10905,4);
TASK_PP(16'h10906,4);
TASK_PP(16'h10907,4);
TASK_PP(16'h10908,4);
TASK_PP(16'h10909,4);
TASK_PP(16'h1090A,4);
TASK_PP(16'h1090B,4);
TASK_PP(16'h1090C,4);
TASK_PP(16'h1090D,4);
TASK_PP(16'h1090E,4);
TASK_PP(16'h1090F,4);
TASK_PP(16'h10910,4);
TASK_PP(16'h10911,4);
TASK_PP(16'h10912,4);
TASK_PP(16'h10913,4);
TASK_PP(16'h10914,4);
TASK_PP(16'h10915,4);
TASK_PP(16'h10916,4);
TASK_PP(16'h10917,4);
TASK_PP(16'h10918,4);
TASK_PP(16'h10919,4);
TASK_PP(16'h1091A,4);
TASK_PP(16'h1091B,4);
TASK_PP(16'h1091C,4);
TASK_PP(16'h1091D,4);
TASK_PP(16'h1091E,4);
TASK_PP(16'h1091F,4);
TASK_PP(16'h10920,4);
TASK_PP(16'h10921,4);
TASK_PP(16'h10922,4);
TASK_PP(16'h10923,4);
TASK_PP(16'h10924,4);
TASK_PP(16'h10925,4);
TASK_PP(16'h10926,4);
TASK_PP(16'h10927,4);
TASK_PP(16'h10928,4);
TASK_PP(16'h10929,4);
TASK_PP(16'h1092A,4);
TASK_PP(16'h1092B,4);
TASK_PP(16'h1092C,4);
TASK_PP(16'h1092D,4);
TASK_PP(16'h1092E,4);
TASK_PP(16'h1092F,4);
TASK_PP(16'h10930,4);
TASK_PP(16'h10931,4);
TASK_PP(16'h10932,4);
TASK_PP(16'h10933,4);
TASK_PP(16'h10934,4);
TASK_PP(16'h10935,4);
TASK_PP(16'h10936,4);
TASK_PP(16'h10937,4);
TASK_PP(16'h10938,4);
TASK_PP(16'h10939,4);
TASK_PP(16'h1093A,4);
TASK_PP(16'h1093B,4);
TASK_PP(16'h1093C,4);
TASK_PP(16'h1093D,4);
TASK_PP(16'h1093E,4);
TASK_PP(16'h1093F,4);
TASK_PP(16'h10940,4);
TASK_PP(16'h10941,4);
TASK_PP(16'h10942,4);
TASK_PP(16'h10943,4);
TASK_PP(16'h10944,4);
TASK_PP(16'h10945,4);
TASK_PP(16'h10946,4);
TASK_PP(16'h10947,4);
TASK_PP(16'h10948,4);
TASK_PP(16'h10949,4);
TASK_PP(16'h1094A,4);
TASK_PP(16'h1094B,4);
TASK_PP(16'h1094C,4);
TASK_PP(16'h1094D,4);
TASK_PP(16'h1094E,4);
TASK_PP(16'h1094F,4);
TASK_PP(16'h10950,4);
TASK_PP(16'h10951,4);
TASK_PP(16'h10952,4);
TASK_PP(16'h10953,4);
TASK_PP(16'h10954,4);
TASK_PP(16'h10955,4);
TASK_PP(16'h10956,4);
TASK_PP(16'h10957,4);
TASK_PP(16'h10958,4);
TASK_PP(16'h10959,4);
TASK_PP(16'h1095A,4);
TASK_PP(16'h1095B,4);
TASK_PP(16'h1095C,4);
TASK_PP(16'h1095D,4);
TASK_PP(16'h1095E,4);
TASK_PP(16'h1095F,4);
TASK_PP(16'h10960,4);
TASK_PP(16'h10961,4);
TASK_PP(16'h10962,4);
TASK_PP(16'h10963,4);
TASK_PP(16'h10964,4);
TASK_PP(16'h10965,4);
TASK_PP(16'h10966,4);
TASK_PP(16'h10967,4);
TASK_PP(16'h10968,4);
TASK_PP(16'h10969,4);
TASK_PP(16'h1096A,4);
TASK_PP(16'h1096B,4);
TASK_PP(16'h1096C,4);
TASK_PP(16'h1096D,4);
TASK_PP(16'h1096E,4);
TASK_PP(16'h1096F,4);
TASK_PP(16'h10970,4);
TASK_PP(16'h10971,4);
TASK_PP(16'h10972,4);
TASK_PP(16'h10973,4);
TASK_PP(16'h10974,4);
TASK_PP(16'h10975,4);
TASK_PP(16'h10976,4);
TASK_PP(16'h10977,4);
TASK_PP(16'h10978,4);
TASK_PP(16'h10979,4);
TASK_PP(16'h1097A,4);
TASK_PP(16'h1097B,4);
TASK_PP(16'h1097C,4);
TASK_PP(16'h1097D,4);
TASK_PP(16'h1097E,4);
TASK_PP(16'h1097F,4);
TASK_PP(16'h10980,4);
TASK_PP(16'h10981,4);
TASK_PP(16'h10982,4);
TASK_PP(16'h10983,4);
TASK_PP(16'h10984,4);
TASK_PP(16'h10985,4);
TASK_PP(16'h10986,4);
TASK_PP(16'h10987,4);
TASK_PP(16'h10988,4);
TASK_PP(16'h10989,4);
TASK_PP(16'h1098A,4);
TASK_PP(16'h1098B,4);
TASK_PP(16'h1098C,4);
TASK_PP(16'h1098D,4);
TASK_PP(16'h1098E,4);
TASK_PP(16'h1098F,4);
TASK_PP(16'h10990,4);
TASK_PP(16'h10991,4);
TASK_PP(16'h10992,4);
TASK_PP(16'h10993,4);
TASK_PP(16'h10994,4);
TASK_PP(16'h10995,4);
TASK_PP(16'h10996,4);
TASK_PP(16'h10997,4);
TASK_PP(16'h10998,4);
TASK_PP(16'h10999,4);
TASK_PP(16'h1099A,4);
TASK_PP(16'h1099B,4);
TASK_PP(16'h1099C,4);
TASK_PP(16'h1099D,4);
TASK_PP(16'h1099E,4);
TASK_PP(16'h1099F,4);
TASK_PP(16'h109A0,4);
TASK_PP(16'h109A1,4);
TASK_PP(16'h109A2,4);
TASK_PP(16'h109A3,4);
TASK_PP(16'h109A4,4);
TASK_PP(16'h109A5,4);
TASK_PP(16'h109A6,4);
TASK_PP(16'h109A7,4);
TASK_PP(16'h109A8,4);
TASK_PP(16'h109A9,4);
TASK_PP(16'h109AA,4);
TASK_PP(16'h109AB,4);
TASK_PP(16'h109AC,4);
TASK_PP(16'h109AD,4);
TASK_PP(16'h109AE,4);
TASK_PP(16'h109AF,4);
TASK_PP(16'h109B0,4);
TASK_PP(16'h109B1,4);
TASK_PP(16'h109B2,4);
TASK_PP(16'h109B3,4);
TASK_PP(16'h109B4,4);
TASK_PP(16'h109B5,4);
TASK_PP(16'h109B6,4);
TASK_PP(16'h109B7,4);
TASK_PP(16'h109B8,4);
TASK_PP(16'h109B9,4);
TASK_PP(16'h109BA,4);
TASK_PP(16'h109BB,4);
TASK_PP(16'h109BC,4);
TASK_PP(16'h109BD,4);
TASK_PP(16'h109BE,4);
TASK_PP(16'h109BF,4);
TASK_PP(16'h109C0,4);
TASK_PP(16'h109C1,4);
TASK_PP(16'h109C2,4);
TASK_PP(16'h109C3,4);
TASK_PP(16'h109C4,4);
TASK_PP(16'h109C5,4);
TASK_PP(16'h109C6,4);
TASK_PP(16'h109C7,4);
TASK_PP(16'h109C8,4);
TASK_PP(16'h109C9,4);
TASK_PP(16'h109CA,4);
TASK_PP(16'h109CB,4);
TASK_PP(16'h109CC,4);
TASK_PP(16'h109CD,4);
TASK_PP(16'h109CE,4);
TASK_PP(16'h109CF,4);
TASK_PP(16'h109D0,4);
TASK_PP(16'h109D1,4);
TASK_PP(16'h109D2,4);
TASK_PP(16'h109D3,4);
TASK_PP(16'h109D4,4);
TASK_PP(16'h109D5,4);
TASK_PP(16'h109D6,4);
TASK_PP(16'h109D7,4);
TASK_PP(16'h109D8,4);
TASK_PP(16'h109D9,4);
TASK_PP(16'h109DA,4);
TASK_PP(16'h109DB,4);
TASK_PP(16'h109DC,4);
TASK_PP(16'h109DD,4);
TASK_PP(16'h109DE,4);
TASK_PP(16'h109DF,4);
TASK_PP(16'h109E0,4);
TASK_PP(16'h109E1,4);
TASK_PP(16'h109E2,4);
TASK_PP(16'h109E3,4);
TASK_PP(16'h109E4,4);
TASK_PP(16'h109E5,4);
TASK_PP(16'h109E6,4);
TASK_PP(16'h109E7,4);
TASK_PP(16'h109E8,4);
TASK_PP(16'h109E9,4);
TASK_PP(16'h109EA,4);
TASK_PP(16'h109EB,4);
TASK_PP(16'h109EC,4);
TASK_PP(16'h109ED,4);
TASK_PP(16'h109EE,4);
TASK_PP(16'h109EF,4);
TASK_PP(16'h109F0,4);
TASK_PP(16'h109F1,4);
TASK_PP(16'h109F2,4);
TASK_PP(16'h109F3,4);
TASK_PP(16'h109F4,4);
TASK_PP(16'h109F5,4);
TASK_PP(16'h109F6,4);
TASK_PP(16'h109F7,4);
TASK_PP(16'h109F8,4);
TASK_PP(16'h109F9,4);
TASK_PP(16'h109FA,4);
TASK_PP(16'h109FB,4);
TASK_PP(16'h109FC,4);
TASK_PP(16'h109FD,4);
TASK_PP(16'h109FE,4);
TASK_PP(16'h109FF,4);
TASK_PP(16'h10A00,4);
TASK_PP(16'h10A01,4);
TASK_PP(16'h10A02,4);
TASK_PP(16'h10A03,4);
TASK_PP(16'h10A04,4);
TASK_PP(16'h10A05,4);
TASK_PP(16'h10A06,4);
TASK_PP(16'h10A07,4);
TASK_PP(16'h10A08,4);
TASK_PP(16'h10A09,4);
TASK_PP(16'h10A0A,4);
TASK_PP(16'h10A0B,4);
TASK_PP(16'h10A0C,4);
TASK_PP(16'h10A0D,4);
TASK_PP(16'h10A0E,4);
TASK_PP(16'h10A0F,4);
TASK_PP(16'h10A10,4);
TASK_PP(16'h10A11,4);
TASK_PP(16'h10A12,4);
TASK_PP(16'h10A13,4);
TASK_PP(16'h10A14,4);
TASK_PP(16'h10A15,4);
TASK_PP(16'h10A16,4);
TASK_PP(16'h10A17,4);
TASK_PP(16'h10A18,4);
TASK_PP(16'h10A19,4);
TASK_PP(16'h10A1A,4);
TASK_PP(16'h10A1B,4);
TASK_PP(16'h10A1C,4);
TASK_PP(16'h10A1D,4);
TASK_PP(16'h10A1E,4);
TASK_PP(16'h10A1F,4);
TASK_PP(16'h10A20,4);
TASK_PP(16'h10A21,4);
TASK_PP(16'h10A22,4);
TASK_PP(16'h10A23,4);
TASK_PP(16'h10A24,4);
TASK_PP(16'h10A25,4);
TASK_PP(16'h10A26,4);
TASK_PP(16'h10A27,4);
TASK_PP(16'h10A28,4);
TASK_PP(16'h10A29,4);
TASK_PP(16'h10A2A,4);
TASK_PP(16'h10A2B,4);
TASK_PP(16'h10A2C,4);
TASK_PP(16'h10A2D,4);
TASK_PP(16'h10A2E,4);
TASK_PP(16'h10A2F,4);
TASK_PP(16'h10A30,4);
TASK_PP(16'h10A31,4);
TASK_PP(16'h10A32,4);
TASK_PP(16'h10A33,4);
TASK_PP(16'h10A34,4);
TASK_PP(16'h10A35,4);
TASK_PP(16'h10A36,4);
TASK_PP(16'h10A37,4);
TASK_PP(16'h10A38,4);
TASK_PP(16'h10A39,4);
TASK_PP(16'h10A3A,4);
TASK_PP(16'h10A3B,4);
TASK_PP(16'h10A3C,4);
TASK_PP(16'h10A3D,4);
TASK_PP(16'h10A3E,4);
TASK_PP(16'h10A3F,4);
TASK_PP(16'h10A40,4);
TASK_PP(16'h10A41,4);
TASK_PP(16'h10A42,4);
TASK_PP(16'h10A43,4);
TASK_PP(16'h10A44,4);
TASK_PP(16'h10A45,4);
TASK_PP(16'h10A46,4);
TASK_PP(16'h10A47,4);
TASK_PP(16'h10A48,4);
TASK_PP(16'h10A49,4);
TASK_PP(16'h10A4A,4);
TASK_PP(16'h10A4B,4);
TASK_PP(16'h10A4C,4);
TASK_PP(16'h10A4D,4);
TASK_PP(16'h10A4E,4);
TASK_PP(16'h10A4F,4);
TASK_PP(16'h10A50,4);
TASK_PP(16'h10A51,4);
TASK_PP(16'h10A52,4);
TASK_PP(16'h10A53,4);
TASK_PP(16'h10A54,4);
TASK_PP(16'h10A55,4);
TASK_PP(16'h10A56,4);
TASK_PP(16'h10A57,4);
TASK_PP(16'h10A58,4);
TASK_PP(16'h10A59,4);
TASK_PP(16'h10A5A,4);
TASK_PP(16'h10A5B,4);
TASK_PP(16'h10A5C,4);
TASK_PP(16'h10A5D,4);
TASK_PP(16'h10A5E,4);
TASK_PP(16'h10A5F,4);
TASK_PP(16'h10A60,4);
TASK_PP(16'h10A61,4);
TASK_PP(16'h10A62,4);
TASK_PP(16'h10A63,4);
TASK_PP(16'h10A64,4);
TASK_PP(16'h10A65,4);
TASK_PP(16'h10A66,4);
TASK_PP(16'h10A67,4);
TASK_PP(16'h10A68,4);
TASK_PP(16'h10A69,4);
TASK_PP(16'h10A6A,4);
TASK_PP(16'h10A6B,4);
TASK_PP(16'h10A6C,4);
TASK_PP(16'h10A6D,4);
TASK_PP(16'h10A6E,4);
TASK_PP(16'h10A6F,4);
TASK_PP(16'h10A70,4);
TASK_PP(16'h10A71,4);
TASK_PP(16'h10A72,4);
TASK_PP(16'h10A73,4);
TASK_PP(16'h10A74,4);
TASK_PP(16'h10A75,4);
TASK_PP(16'h10A76,4);
TASK_PP(16'h10A77,4);
TASK_PP(16'h10A78,4);
TASK_PP(16'h10A79,4);
TASK_PP(16'h10A7A,4);
TASK_PP(16'h10A7B,4);
TASK_PP(16'h10A7C,4);
TASK_PP(16'h10A7D,4);
TASK_PP(16'h10A7E,4);
TASK_PP(16'h10A7F,4);
TASK_PP(16'h10A80,4);
TASK_PP(16'h10A81,4);
TASK_PP(16'h10A82,4);
TASK_PP(16'h10A83,4);
TASK_PP(16'h10A84,4);
TASK_PP(16'h10A85,4);
TASK_PP(16'h10A86,4);
TASK_PP(16'h10A87,4);
TASK_PP(16'h10A88,4);
TASK_PP(16'h10A89,4);
TASK_PP(16'h10A8A,4);
TASK_PP(16'h10A8B,4);
TASK_PP(16'h10A8C,4);
TASK_PP(16'h10A8D,4);
TASK_PP(16'h10A8E,4);
TASK_PP(16'h10A8F,4);
TASK_PP(16'h10A90,4);
TASK_PP(16'h10A91,4);
TASK_PP(16'h10A92,4);
TASK_PP(16'h10A93,4);
TASK_PP(16'h10A94,4);
TASK_PP(16'h10A95,4);
TASK_PP(16'h10A96,4);
TASK_PP(16'h10A97,4);
TASK_PP(16'h10A98,4);
TASK_PP(16'h10A99,4);
TASK_PP(16'h10A9A,4);
TASK_PP(16'h10A9B,4);
TASK_PP(16'h10A9C,4);
TASK_PP(16'h10A9D,4);
TASK_PP(16'h10A9E,4);
TASK_PP(16'h10A9F,4);
TASK_PP(16'h10AA0,4);
TASK_PP(16'h10AA1,4);
TASK_PP(16'h10AA2,4);
TASK_PP(16'h10AA3,4);
TASK_PP(16'h10AA4,4);
TASK_PP(16'h10AA5,4);
TASK_PP(16'h10AA6,4);
TASK_PP(16'h10AA7,4);
TASK_PP(16'h10AA8,4);
TASK_PP(16'h10AA9,4);
TASK_PP(16'h10AAA,4);
TASK_PP(16'h10AAB,4);
TASK_PP(16'h10AAC,4);
TASK_PP(16'h10AAD,4);
TASK_PP(16'h10AAE,4);
TASK_PP(16'h10AAF,4);
TASK_PP(16'h10AB0,4);
TASK_PP(16'h10AB1,4);
TASK_PP(16'h10AB2,4);
TASK_PP(16'h10AB3,4);
TASK_PP(16'h10AB4,4);
TASK_PP(16'h10AB5,4);
TASK_PP(16'h10AB6,4);
TASK_PP(16'h10AB7,4);
TASK_PP(16'h10AB8,4);
TASK_PP(16'h10AB9,4);
TASK_PP(16'h10ABA,4);
TASK_PP(16'h10ABB,4);
TASK_PP(16'h10ABC,4);
TASK_PP(16'h10ABD,4);
TASK_PP(16'h10ABE,4);
TASK_PP(16'h10ABF,4);
TASK_PP(16'h10AC0,4);
TASK_PP(16'h10AC1,4);
TASK_PP(16'h10AC2,4);
TASK_PP(16'h10AC3,4);
TASK_PP(16'h10AC4,4);
TASK_PP(16'h10AC5,4);
TASK_PP(16'h10AC6,4);
TASK_PP(16'h10AC7,4);
TASK_PP(16'h10AC8,4);
TASK_PP(16'h10AC9,4);
TASK_PP(16'h10ACA,4);
TASK_PP(16'h10ACB,4);
TASK_PP(16'h10ACC,4);
TASK_PP(16'h10ACD,4);
TASK_PP(16'h10ACE,4);
TASK_PP(16'h10ACF,4);
TASK_PP(16'h10AD0,4);
TASK_PP(16'h10AD1,4);
TASK_PP(16'h10AD2,4);
TASK_PP(16'h10AD3,4);
TASK_PP(16'h10AD4,4);
TASK_PP(16'h10AD5,4);
TASK_PP(16'h10AD6,4);
TASK_PP(16'h10AD7,4);
TASK_PP(16'h10AD8,4);
TASK_PP(16'h10AD9,4);
TASK_PP(16'h10ADA,4);
TASK_PP(16'h10ADB,4);
TASK_PP(16'h10ADC,4);
TASK_PP(16'h10ADD,4);
TASK_PP(16'h10ADE,4);
TASK_PP(16'h10ADF,4);
TASK_PP(16'h10AE0,4);
TASK_PP(16'h10AE1,4);
TASK_PP(16'h10AE2,4);
TASK_PP(16'h10AE3,4);
TASK_PP(16'h10AE4,4);
TASK_PP(16'h10AE5,4);
TASK_PP(16'h10AE6,4);
TASK_PP(16'h10AE7,4);
TASK_PP(16'h10AE8,4);
TASK_PP(16'h10AE9,4);
TASK_PP(16'h10AEA,4);
TASK_PP(16'h10AEB,4);
TASK_PP(16'h10AEC,4);
TASK_PP(16'h10AED,4);
TASK_PP(16'h10AEE,4);
TASK_PP(16'h10AEF,4);
TASK_PP(16'h10AF0,4);
TASK_PP(16'h10AF1,4);
TASK_PP(16'h10AF2,4);
TASK_PP(16'h10AF3,4);
TASK_PP(16'h10AF4,4);
TASK_PP(16'h10AF5,4);
TASK_PP(16'h10AF6,4);
TASK_PP(16'h10AF7,4);
TASK_PP(16'h10AF8,4);
TASK_PP(16'h10AF9,4);
TASK_PP(16'h10AFA,4);
TASK_PP(16'h10AFB,4);
TASK_PP(16'h10AFC,4);
TASK_PP(16'h10AFD,4);
TASK_PP(16'h10AFE,4);
TASK_PP(16'h10AFF,4);
TASK_PP(16'h10B00,4);
TASK_PP(16'h10B01,4);
TASK_PP(16'h10B02,4);
TASK_PP(16'h10B03,4);
TASK_PP(16'h10B04,4);
TASK_PP(16'h10B05,4);
TASK_PP(16'h10B06,4);
TASK_PP(16'h10B07,4);
TASK_PP(16'h10B08,4);
TASK_PP(16'h10B09,4);
TASK_PP(16'h10B0A,4);
TASK_PP(16'h10B0B,4);
TASK_PP(16'h10B0C,4);
TASK_PP(16'h10B0D,4);
TASK_PP(16'h10B0E,4);
TASK_PP(16'h10B0F,4);
TASK_PP(16'h10B10,4);
TASK_PP(16'h10B11,4);
TASK_PP(16'h10B12,4);
TASK_PP(16'h10B13,4);
TASK_PP(16'h10B14,4);
TASK_PP(16'h10B15,4);
TASK_PP(16'h10B16,4);
TASK_PP(16'h10B17,4);
TASK_PP(16'h10B18,4);
TASK_PP(16'h10B19,4);
TASK_PP(16'h10B1A,4);
TASK_PP(16'h10B1B,4);
TASK_PP(16'h10B1C,4);
TASK_PP(16'h10B1D,4);
TASK_PP(16'h10B1E,4);
TASK_PP(16'h10B1F,4);
TASK_PP(16'h10B20,4);
TASK_PP(16'h10B21,4);
TASK_PP(16'h10B22,4);
TASK_PP(16'h10B23,4);
TASK_PP(16'h10B24,4);
TASK_PP(16'h10B25,4);
TASK_PP(16'h10B26,4);
TASK_PP(16'h10B27,4);
TASK_PP(16'h10B28,4);
TASK_PP(16'h10B29,4);
TASK_PP(16'h10B2A,4);
TASK_PP(16'h10B2B,4);
TASK_PP(16'h10B2C,4);
TASK_PP(16'h10B2D,4);
TASK_PP(16'h10B2E,4);
TASK_PP(16'h10B2F,4);
TASK_PP(16'h10B30,4);
TASK_PP(16'h10B31,4);
TASK_PP(16'h10B32,4);
TASK_PP(16'h10B33,4);
TASK_PP(16'h10B34,4);
TASK_PP(16'h10B35,4);
TASK_PP(16'h10B36,4);
TASK_PP(16'h10B37,4);
TASK_PP(16'h10B38,4);
TASK_PP(16'h10B39,4);
TASK_PP(16'h10B3A,4);
TASK_PP(16'h10B3B,4);
TASK_PP(16'h10B3C,4);
TASK_PP(16'h10B3D,4);
TASK_PP(16'h10B3E,4);
TASK_PP(16'h10B3F,4);
TASK_PP(16'h10B40,4);
TASK_PP(16'h10B41,4);
TASK_PP(16'h10B42,4);
TASK_PP(16'h10B43,4);
TASK_PP(16'h10B44,4);
TASK_PP(16'h10B45,4);
TASK_PP(16'h10B46,4);
TASK_PP(16'h10B47,4);
TASK_PP(16'h10B48,4);
TASK_PP(16'h10B49,4);
TASK_PP(16'h10B4A,4);
TASK_PP(16'h10B4B,4);
TASK_PP(16'h10B4C,4);
TASK_PP(16'h10B4D,4);
TASK_PP(16'h10B4E,4);
TASK_PP(16'h10B4F,4);
TASK_PP(16'h10B50,4);
TASK_PP(16'h10B51,4);
TASK_PP(16'h10B52,4);
TASK_PP(16'h10B53,4);
TASK_PP(16'h10B54,4);
TASK_PP(16'h10B55,4);
TASK_PP(16'h10B56,4);
TASK_PP(16'h10B57,4);
TASK_PP(16'h10B58,4);
TASK_PP(16'h10B59,4);
TASK_PP(16'h10B5A,4);
TASK_PP(16'h10B5B,4);
TASK_PP(16'h10B5C,4);
TASK_PP(16'h10B5D,4);
TASK_PP(16'h10B5E,4);
TASK_PP(16'h10B5F,4);
TASK_PP(16'h10B60,4);
TASK_PP(16'h10B61,4);
TASK_PP(16'h10B62,4);
TASK_PP(16'h10B63,4);
TASK_PP(16'h10B64,4);
TASK_PP(16'h10B65,4);
TASK_PP(16'h10B66,4);
TASK_PP(16'h10B67,4);
TASK_PP(16'h10B68,4);
TASK_PP(16'h10B69,4);
TASK_PP(16'h10B6A,4);
TASK_PP(16'h10B6B,4);
TASK_PP(16'h10B6C,4);
TASK_PP(16'h10B6D,4);
TASK_PP(16'h10B6E,4);
TASK_PP(16'h10B6F,4);
TASK_PP(16'h10B70,4);
TASK_PP(16'h10B71,4);
TASK_PP(16'h10B72,4);
TASK_PP(16'h10B73,4);
TASK_PP(16'h10B74,4);
TASK_PP(16'h10B75,4);
TASK_PP(16'h10B76,4);
TASK_PP(16'h10B77,4);
TASK_PP(16'h10B78,4);
TASK_PP(16'h10B79,4);
TASK_PP(16'h10B7A,4);
TASK_PP(16'h10B7B,4);
TASK_PP(16'h10B7C,4);
TASK_PP(16'h10B7D,4);
TASK_PP(16'h10B7E,4);
TASK_PP(16'h10B7F,4);
TASK_PP(16'h10B80,4);
TASK_PP(16'h10B81,4);
TASK_PP(16'h10B82,4);
TASK_PP(16'h10B83,4);
TASK_PP(16'h10B84,4);
TASK_PP(16'h10B85,4);
TASK_PP(16'h10B86,4);
TASK_PP(16'h10B87,4);
TASK_PP(16'h10B88,4);
TASK_PP(16'h10B89,4);
TASK_PP(16'h10B8A,4);
TASK_PP(16'h10B8B,4);
TASK_PP(16'h10B8C,4);
TASK_PP(16'h10B8D,4);
TASK_PP(16'h10B8E,4);
TASK_PP(16'h10B8F,4);
TASK_PP(16'h10B90,4);
TASK_PP(16'h10B91,4);
TASK_PP(16'h10B92,4);
TASK_PP(16'h10B93,4);
TASK_PP(16'h10B94,4);
TASK_PP(16'h10B95,4);
TASK_PP(16'h10B96,4);
TASK_PP(16'h10B97,4);
TASK_PP(16'h10B98,4);
TASK_PP(16'h10B99,4);
TASK_PP(16'h10B9A,4);
TASK_PP(16'h10B9B,4);
TASK_PP(16'h10B9C,4);
TASK_PP(16'h10B9D,4);
TASK_PP(16'h10B9E,4);
TASK_PP(16'h10B9F,4);
TASK_PP(16'h10BA0,4);
TASK_PP(16'h10BA1,4);
TASK_PP(16'h10BA2,4);
TASK_PP(16'h10BA3,4);
TASK_PP(16'h10BA4,4);
TASK_PP(16'h10BA5,4);
TASK_PP(16'h10BA6,4);
TASK_PP(16'h10BA7,4);
TASK_PP(16'h10BA8,4);
TASK_PP(16'h10BA9,4);
TASK_PP(16'h10BAA,4);
TASK_PP(16'h10BAB,4);
TASK_PP(16'h10BAC,4);
TASK_PP(16'h10BAD,4);
TASK_PP(16'h10BAE,4);
TASK_PP(16'h10BAF,4);
TASK_PP(16'h10BB0,4);
TASK_PP(16'h10BB1,4);
TASK_PP(16'h10BB2,4);
TASK_PP(16'h10BB3,4);
TASK_PP(16'h10BB4,4);
TASK_PP(16'h10BB5,4);
TASK_PP(16'h10BB6,4);
TASK_PP(16'h10BB7,4);
TASK_PP(16'h10BB8,4);
TASK_PP(16'h10BB9,4);
TASK_PP(16'h10BBA,4);
TASK_PP(16'h10BBB,4);
TASK_PP(16'h10BBC,4);
TASK_PP(16'h10BBD,4);
TASK_PP(16'h10BBE,4);
TASK_PP(16'h10BBF,4);
TASK_PP(16'h10BC0,4);
TASK_PP(16'h10BC1,4);
TASK_PP(16'h10BC2,4);
TASK_PP(16'h10BC3,4);
TASK_PP(16'h10BC4,4);
TASK_PP(16'h10BC5,4);
TASK_PP(16'h10BC6,4);
TASK_PP(16'h10BC7,4);
TASK_PP(16'h10BC8,4);
TASK_PP(16'h10BC9,4);
TASK_PP(16'h10BCA,4);
TASK_PP(16'h10BCB,4);
TASK_PP(16'h10BCC,4);
TASK_PP(16'h10BCD,4);
TASK_PP(16'h10BCE,4);
TASK_PP(16'h10BCF,4);
TASK_PP(16'h10BD0,4);
TASK_PP(16'h10BD1,4);
TASK_PP(16'h10BD2,4);
TASK_PP(16'h10BD3,4);
TASK_PP(16'h10BD4,4);
TASK_PP(16'h10BD5,4);
TASK_PP(16'h10BD6,4);
TASK_PP(16'h10BD7,4);
TASK_PP(16'h10BD8,4);
TASK_PP(16'h10BD9,4);
TASK_PP(16'h10BDA,4);
TASK_PP(16'h10BDB,4);
TASK_PP(16'h10BDC,4);
TASK_PP(16'h10BDD,4);
TASK_PP(16'h10BDE,4);
TASK_PP(16'h10BDF,4);
TASK_PP(16'h10BE0,4);
TASK_PP(16'h10BE1,4);
TASK_PP(16'h10BE2,4);
TASK_PP(16'h10BE3,4);
TASK_PP(16'h10BE4,4);
TASK_PP(16'h10BE5,4);
TASK_PP(16'h10BE6,4);
TASK_PP(16'h10BE7,4);
TASK_PP(16'h10BE8,4);
TASK_PP(16'h10BE9,4);
TASK_PP(16'h10BEA,4);
TASK_PP(16'h10BEB,4);
TASK_PP(16'h10BEC,4);
TASK_PP(16'h10BED,4);
TASK_PP(16'h10BEE,4);
TASK_PP(16'h10BEF,4);
TASK_PP(16'h10BF0,4);
TASK_PP(16'h10BF1,4);
TASK_PP(16'h10BF2,4);
TASK_PP(16'h10BF3,4);
TASK_PP(16'h10BF4,4);
TASK_PP(16'h10BF5,4);
TASK_PP(16'h10BF6,4);
TASK_PP(16'h10BF7,4);
TASK_PP(16'h10BF8,4);
TASK_PP(16'h10BF9,4);
TASK_PP(16'h10BFA,4);
TASK_PP(16'h10BFB,4);
TASK_PP(16'h10BFC,4);
TASK_PP(16'h10BFD,4);
TASK_PP(16'h10BFE,4);
TASK_PP(16'h10BFF,4);
TASK_PP(16'h10C00,4);
TASK_PP(16'h10C01,4);
TASK_PP(16'h10C02,4);
TASK_PP(16'h10C03,4);
TASK_PP(16'h10C04,4);
TASK_PP(16'h10C05,4);
TASK_PP(16'h10C06,4);
TASK_PP(16'h10C07,4);
TASK_PP(16'h10C08,4);
TASK_PP(16'h10C09,4);
TASK_PP(16'h10C0A,4);
TASK_PP(16'h10C0B,4);
TASK_PP(16'h10C0C,4);
TASK_PP(16'h10C0D,4);
TASK_PP(16'h10C0E,4);
TASK_PP(16'h10C0F,4);
TASK_PP(16'h10C10,4);
TASK_PP(16'h10C11,4);
TASK_PP(16'h10C12,4);
TASK_PP(16'h10C13,4);
TASK_PP(16'h10C14,4);
TASK_PP(16'h10C15,4);
TASK_PP(16'h10C16,4);
TASK_PP(16'h10C17,4);
TASK_PP(16'h10C18,4);
TASK_PP(16'h10C19,4);
TASK_PP(16'h10C1A,4);
TASK_PP(16'h10C1B,4);
TASK_PP(16'h10C1C,4);
TASK_PP(16'h10C1D,4);
TASK_PP(16'h10C1E,4);
TASK_PP(16'h10C1F,4);
TASK_PP(16'h10C20,4);
TASK_PP(16'h10C21,4);
TASK_PP(16'h10C22,4);
TASK_PP(16'h10C23,4);
TASK_PP(16'h10C24,4);
TASK_PP(16'h10C25,4);
TASK_PP(16'h10C26,4);
TASK_PP(16'h10C27,4);
TASK_PP(16'h10C28,4);
TASK_PP(16'h10C29,4);
TASK_PP(16'h10C2A,4);
TASK_PP(16'h10C2B,4);
TASK_PP(16'h10C2C,4);
TASK_PP(16'h10C2D,4);
TASK_PP(16'h10C2E,4);
TASK_PP(16'h10C2F,4);
TASK_PP(16'h10C30,4);
TASK_PP(16'h10C31,4);
TASK_PP(16'h10C32,4);
TASK_PP(16'h10C33,4);
TASK_PP(16'h10C34,4);
TASK_PP(16'h10C35,4);
TASK_PP(16'h10C36,4);
TASK_PP(16'h10C37,4);
TASK_PP(16'h10C38,4);
TASK_PP(16'h10C39,4);
TASK_PP(16'h10C3A,4);
TASK_PP(16'h10C3B,4);
TASK_PP(16'h10C3C,4);
TASK_PP(16'h10C3D,4);
TASK_PP(16'h10C3E,4);
TASK_PP(16'h10C3F,4);
TASK_PP(16'h10C40,4);
TASK_PP(16'h10C41,4);
TASK_PP(16'h10C42,4);
TASK_PP(16'h10C43,4);
TASK_PP(16'h10C44,4);
TASK_PP(16'h10C45,4);
TASK_PP(16'h10C46,4);
TASK_PP(16'h10C47,4);
TASK_PP(16'h10C48,4);
TASK_PP(16'h10C49,4);
TASK_PP(16'h10C4A,4);
TASK_PP(16'h10C4B,4);
TASK_PP(16'h10C4C,4);
TASK_PP(16'h10C4D,4);
TASK_PP(16'h10C4E,4);
TASK_PP(16'h10C4F,4);
TASK_PP(16'h10C50,4);
TASK_PP(16'h10C51,4);
TASK_PP(16'h10C52,4);
TASK_PP(16'h10C53,4);
TASK_PP(16'h10C54,4);
TASK_PP(16'h10C55,4);
TASK_PP(16'h10C56,4);
TASK_PP(16'h10C57,4);
TASK_PP(16'h10C58,4);
TASK_PP(16'h10C59,4);
TASK_PP(16'h10C5A,4);
TASK_PP(16'h10C5B,4);
TASK_PP(16'h10C5C,4);
TASK_PP(16'h10C5D,4);
TASK_PP(16'h10C5E,4);
TASK_PP(16'h10C5F,4);
TASK_PP(16'h10C60,4);
TASK_PP(16'h10C61,4);
TASK_PP(16'h10C62,4);
TASK_PP(16'h10C63,4);
TASK_PP(16'h10C64,4);
TASK_PP(16'h10C65,4);
TASK_PP(16'h10C66,4);
TASK_PP(16'h10C67,4);
TASK_PP(16'h10C68,4);
TASK_PP(16'h10C69,4);
TASK_PP(16'h10C6A,4);
TASK_PP(16'h10C6B,4);
TASK_PP(16'h10C6C,4);
TASK_PP(16'h10C6D,4);
TASK_PP(16'h10C6E,4);
TASK_PP(16'h10C6F,4);
TASK_PP(16'h10C70,4);
TASK_PP(16'h10C71,4);
TASK_PP(16'h10C72,4);
TASK_PP(16'h10C73,4);
TASK_PP(16'h10C74,4);
TASK_PP(16'h10C75,4);
TASK_PP(16'h10C76,4);
TASK_PP(16'h10C77,4);
TASK_PP(16'h10C78,4);
TASK_PP(16'h10C79,4);
TASK_PP(16'h10C7A,4);
TASK_PP(16'h10C7B,4);
TASK_PP(16'h10C7C,4);
TASK_PP(16'h10C7D,4);
TASK_PP(16'h10C7E,4);
TASK_PP(16'h10C7F,4);
TASK_PP(16'h10C80,4);
TASK_PP(16'h10C81,4);
TASK_PP(16'h10C82,4);
TASK_PP(16'h10C83,4);
TASK_PP(16'h10C84,4);
TASK_PP(16'h10C85,4);
TASK_PP(16'h10C86,4);
TASK_PP(16'h10C87,4);
TASK_PP(16'h10C88,4);
TASK_PP(16'h10C89,4);
TASK_PP(16'h10C8A,4);
TASK_PP(16'h10C8B,4);
TASK_PP(16'h10C8C,4);
TASK_PP(16'h10C8D,4);
TASK_PP(16'h10C8E,4);
TASK_PP(16'h10C8F,4);
TASK_PP(16'h10C90,4);
TASK_PP(16'h10C91,4);
TASK_PP(16'h10C92,4);
TASK_PP(16'h10C93,4);
TASK_PP(16'h10C94,4);
TASK_PP(16'h10C95,4);
TASK_PP(16'h10C96,4);
TASK_PP(16'h10C97,4);
TASK_PP(16'h10C98,4);
TASK_PP(16'h10C99,4);
TASK_PP(16'h10C9A,4);
TASK_PP(16'h10C9B,4);
TASK_PP(16'h10C9C,4);
TASK_PP(16'h10C9D,4);
TASK_PP(16'h10C9E,4);
TASK_PP(16'h10C9F,4);
TASK_PP(16'h10CA0,4);
TASK_PP(16'h10CA1,4);
TASK_PP(16'h10CA2,4);
TASK_PP(16'h10CA3,4);
TASK_PP(16'h10CA4,4);
TASK_PP(16'h10CA5,4);
TASK_PP(16'h10CA6,4);
TASK_PP(16'h10CA7,4);
TASK_PP(16'h10CA8,4);
TASK_PP(16'h10CA9,4);
TASK_PP(16'h10CAA,4);
TASK_PP(16'h10CAB,4);
TASK_PP(16'h10CAC,4);
TASK_PP(16'h10CAD,4);
TASK_PP(16'h10CAE,4);
TASK_PP(16'h10CAF,4);
TASK_PP(16'h10CB0,4);
TASK_PP(16'h10CB1,4);
TASK_PP(16'h10CB2,4);
TASK_PP(16'h10CB3,4);
TASK_PP(16'h10CB4,4);
TASK_PP(16'h10CB5,4);
TASK_PP(16'h10CB6,4);
TASK_PP(16'h10CB7,4);
TASK_PP(16'h10CB8,4);
TASK_PP(16'h10CB9,4);
TASK_PP(16'h10CBA,4);
TASK_PP(16'h10CBB,4);
TASK_PP(16'h10CBC,4);
TASK_PP(16'h10CBD,4);
TASK_PP(16'h10CBE,4);
TASK_PP(16'h10CBF,4);
TASK_PP(16'h10CC0,4);
TASK_PP(16'h10CC1,4);
TASK_PP(16'h10CC2,4);
TASK_PP(16'h10CC3,4);
TASK_PP(16'h10CC4,4);
TASK_PP(16'h10CC5,4);
TASK_PP(16'h10CC6,4);
TASK_PP(16'h10CC7,4);
TASK_PP(16'h10CC8,4);
TASK_PP(16'h10CC9,4);
TASK_PP(16'h10CCA,4);
TASK_PP(16'h10CCB,4);
TASK_PP(16'h10CCC,4);
TASK_PP(16'h10CCD,4);
TASK_PP(16'h10CCE,4);
TASK_PP(16'h10CCF,4);
TASK_PP(16'h10CD0,4);
TASK_PP(16'h10CD1,4);
TASK_PP(16'h10CD2,4);
TASK_PP(16'h10CD3,4);
TASK_PP(16'h10CD4,4);
TASK_PP(16'h10CD5,4);
TASK_PP(16'h10CD6,4);
TASK_PP(16'h10CD7,4);
TASK_PP(16'h10CD8,4);
TASK_PP(16'h10CD9,4);
TASK_PP(16'h10CDA,4);
TASK_PP(16'h10CDB,4);
TASK_PP(16'h10CDC,4);
TASK_PP(16'h10CDD,4);
TASK_PP(16'h10CDE,4);
TASK_PP(16'h10CDF,4);
TASK_PP(16'h10CE0,4);
TASK_PP(16'h10CE1,4);
TASK_PP(16'h10CE2,4);
TASK_PP(16'h10CE3,4);
TASK_PP(16'h10CE4,4);
TASK_PP(16'h10CE5,4);
TASK_PP(16'h10CE6,4);
TASK_PP(16'h10CE7,4);
TASK_PP(16'h10CE8,4);
TASK_PP(16'h10CE9,4);
TASK_PP(16'h10CEA,4);
TASK_PP(16'h10CEB,4);
TASK_PP(16'h10CEC,4);
TASK_PP(16'h10CED,4);
TASK_PP(16'h10CEE,4);
TASK_PP(16'h10CEF,4);
TASK_PP(16'h10CF0,4);
TASK_PP(16'h10CF1,4);
TASK_PP(16'h10CF2,4);
TASK_PP(16'h10CF3,4);
TASK_PP(16'h10CF4,4);
TASK_PP(16'h10CF5,4);
TASK_PP(16'h10CF6,4);
TASK_PP(16'h10CF7,4);
TASK_PP(16'h10CF8,4);
TASK_PP(16'h10CF9,4);
TASK_PP(16'h10CFA,4);
TASK_PP(16'h10CFB,4);
TASK_PP(16'h10CFC,4);
TASK_PP(16'h10CFD,4);
TASK_PP(16'h10CFE,4);
TASK_PP(16'h10CFF,4);
TASK_PP(16'h10D00,4);
TASK_PP(16'h10D01,4);
TASK_PP(16'h10D02,4);
TASK_PP(16'h10D03,4);
TASK_PP(16'h10D04,4);
TASK_PP(16'h10D05,4);
TASK_PP(16'h10D06,4);
TASK_PP(16'h10D07,4);
TASK_PP(16'h10D08,4);
TASK_PP(16'h10D09,4);
TASK_PP(16'h10D0A,4);
TASK_PP(16'h10D0B,4);
TASK_PP(16'h10D0C,4);
TASK_PP(16'h10D0D,4);
TASK_PP(16'h10D0E,4);
TASK_PP(16'h10D0F,4);
TASK_PP(16'h10D10,4);
TASK_PP(16'h10D11,4);
TASK_PP(16'h10D12,4);
TASK_PP(16'h10D13,4);
TASK_PP(16'h10D14,4);
TASK_PP(16'h10D15,4);
TASK_PP(16'h10D16,4);
TASK_PP(16'h10D17,4);
TASK_PP(16'h10D18,4);
TASK_PP(16'h10D19,4);
TASK_PP(16'h10D1A,4);
TASK_PP(16'h10D1B,4);
TASK_PP(16'h10D1C,4);
TASK_PP(16'h10D1D,4);
TASK_PP(16'h10D1E,4);
TASK_PP(16'h10D1F,4);
TASK_PP(16'h10D20,4);
TASK_PP(16'h10D21,4);
TASK_PP(16'h10D22,4);
TASK_PP(16'h10D23,4);
TASK_PP(16'h10D24,4);
TASK_PP(16'h10D25,4);
TASK_PP(16'h10D26,4);
TASK_PP(16'h10D27,4);
TASK_PP(16'h10D28,4);
TASK_PP(16'h10D29,4);
TASK_PP(16'h10D2A,4);
TASK_PP(16'h10D2B,4);
TASK_PP(16'h10D2C,4);
TASK_PP(16'h10D2D,4);
TASK_PP(16'h10D2E,4);
TASK_PP(16'h10D2F,4);
TASK_PP(16'h10D30,4);
TASK_PP(16'h10D31,4);
TASK_PP(16'h10D32,4);
TASK_PP(16'h10D33,4);
TASK_PP(16'h10D34,4);
TASK_PP(16'h10D35,4);
TASK_PP(16'h10D36,4);
TASK_PP(16'h10D37,4);
TASK_PP(16'h10D38,4);
TASK_PP(16'h10D39,4);
TASK_PP(16'h10D3A,4);
TASK_PP(16'h10D3B,4);
TASK_PP(16'h10D3C,4);
TASK_PP(16'h10D3D,4);
TASK_PP(16'h10D3E,4);
TASK_PP(16'h10D3F,4);
TASK_PP(16'h10D40,4);
TASK_PP(16'h10D41,4);
TASK_PP(16'h10D42,4);
TASK_PP(16'h10D43,4);
TASK_PP(16'h10D44,4);
TASK_PP(16'h10D45,4);
TASK_PP(16'h10D46,4);
TASK_PP(16'h10D47,4);
TASK_PP(16'h10D48,4);
TASK_PP(16'h10D49,4);
TASK_PP(16'h10D4A,4);
TASK_PP(16'h10D4B,4);
TASK_PP(16'h10D4C,4);
TASK_PP(16'h10D4D,4);
TASK_PP(16'h10D4E,4);
TASK_PP(16'h10D4F,4);
TASK_PP(16'h10D50,4);
TASK_PP(16'h10D51,4);
TASK_PP(16'h10D52,4);
TASK_PP(16'h10D53,4);
TASK_PP(16'h10D54,4);
TASK_PP(16'h10D55,4);
TASK_PP(16'h10D56,4);
TASK_PP(16'h10D57,4);
TASK_PP(16'h10D58,4);
TASK_PP(16'h10D59,4);
TASK_PP(16'h10D5A,4);
TASK_PP(16'h10D5B,4);
TASK_PP(16'h10D5C,4);
TASK_PP(16'h10D5D,4);
TASK_PP(16'h10D5E,4);
TASK_PP(16'h10D5F,4);
TASK_PP(16'h10D60,4);
TASK_PP(16'h10D61,4);
TASK_PP(16'h10D62,4);
TASK_PP(16'h10D63,4);
TASK_PP(16'h10D64,4);
TASK_PP(16'h10D65,4);
TASK_PP(16'h10D66,4);
TASK_PP(16'h10D67,4);
TASK_PP(16'h10D68,4);
TASK_PP(16'h10D69,4);
TASK_PP(16'h10D6A,4);
TASK_PP(16'h10D6B,4);
TASK_PP(16'h10D6C,4);
TASK_PP(16'h10D6D,4);
TASK_PP(16'h10D6E,4);
TASK_PP(16'h10D6F,4);
TASK_PP(16'h10D70,4);
TASK_PP(16'h10D71,4);
TASK_PP(16'h10D72,4);
TASK_PP(16'h10D73,4);
TASK_PP(16'h10D74,4);
TASK_PP(16'h10D75,4);
TASK_PP(16'h10D76,4);
TASK_PP(16'h10D77,4);
TASK_PP(16'h10D78,4);
TASK_PP(16'h10D79,4);
TASK_PP(16'h10D7A,4);
TASK_PP(16'h10D7B,4);
TASK_PP(16'h10D7C,4);
TASK_PP(16'h10D7D,4);
TASK_PP(16'h10D7E,4);
TASK_PP(16'h10D7F,4);
TASK_PP(16'h10D80,4);
TASK_PP(16'h10D81,4);
TASK_PP(16'h10D82,4);
TASK_PP(16'h10D83,4);
TASK_PP(16'h10D84,4);
TASK_PP(16'h10D85,4);
TASK_PP(16'h10D86,4);
TASK_PP(16'h10D87,4);
TASK_PP(16'h10D88,4);
TASK_PP(16'h10D89,4);
TASK_PP(16'h10D8A,4);
TASK_PP(16'h10D8B,4);
TASK_PP(16'h10D8C,4);
TASK_PP(16'h10D8D,4);
TASK_PP(16'h10D8E,4);
TASK_PP(16'h10D8F,4);
TASK_PP(16'h10D90,4);
TASK_PP(16'h10D91,4);
TASK_PP(16'h10D92,4);
TASK_PP(16'h10D93,4);
TASK_PP(16'h10D94,4);
TASK_PP(16'h10D95,4);
TASK_PP(16'h10D96,4);
TASK_PP(16'h10D97,4);
TASK_PP(16'h10D98,4);
TASK_PP(16'h10D99,4);
TASK_PP(16'h10D9A,4);
TASK_PP(16'h10D9B,4);
TASK_PP(16'h10D9C,4);
TASK_PP(16'h10D9D,4);
TASK_PP(16'h10D9E,4);
TASK_PP(16'h10D9F,4);
TASK_PP(16'h10DA0,4);
TASK_PP(16'h10DA1,4);
TASK_PP(16'h10DA2,4);
TASK_PP(16'h10DA3,4);
TASK_PP(16'h10DA4,4);
TASK_PP(16'h10DA5,4);
TASK_PP(16'h10DA6,4);
TASK_PP(16'h10DA7,4);
TASK_PP(16'h10DA8,4);
TASK_PP(16'h10DA9,4);
TASK_PP(16'h10DAA,4);
TASK_PP(16'h10DAB,4);
TASK_PP(16'h10DAC,4);
TASK_PP(16'h10DAD,4);
TASK_PP(16'h10DAE,4);
TASK_PP(16'h10DAF,4);
TASK_PP(16'h10DB0,4);
TASK_PP(16'h10DB1,4);
TASK_PP(16'h10DB2,4);
TASK_PP(16'h10DB3,4);
TASK_PP(16'h10DB4,4);
TASK_PP(16'h10DB5,4);
TASK_PP(16'h10DB6,4);
TASK_PP(16'h10DB7,4);
TASK_PP(16'h10DB8,4);
TASK_PP(16'h10DB9,4);
TASK_PP(16'h10DBA,4);
TASK_PP(16'h10DBB,4);
TASK_PP(16'h10DBC,4);
TASK_PP(16'h10DBD,4);
TASK_PP(16'h10DBE,4);
TASK_PP(16'h10DBF,4);
TASK_PP(16'h10DC0,4);
TASK_PP(16'h10DC1,4);
TASK_PP(16'h10DC2,4);
TASK_PP(16'h10DC3,4);
TASK_PP(16'h10DC4,4);
TASK_PP(16'h10DC5,4);
TASK_PP(16'h10DC6,4);
TASK_PP(16'h10DC7,4);
TASK_PP(16'h10DC8,4);
TASK_PP(16'h10DC9,4);
TASK_PP(16'h10DCA,4);
TASK_PP(16'h10DCB,4);
TASK_PP(16'h10DCC,4);
TASK_PP(16'h10DCD,4);
TASK_PP(16'h10DCE,4);
TASK_PP(16'h10DCF,4);
TASK_PP(16'h10DD0,4);
TASK_PP(16'h10DD1,4);
TASK_PP(16'h10DD2,4);
TASK_PP(16'h10DD3,4);
TASK_PP(16'h10DD4,4);
TASK_PP(16'h10DD5,4);
TASK_PP(16'h10DD6,4);
TASK_PP(16'h10DD7,4);
TASK_PP(16'h10DD8,4);
TASK_PP(16'h10DD9,4);
TASK_PP(16'h10DDA,4);
TASK_PP(16'h10DDB,4);
TASK_PP(16'h10DDC,4);
TASK_PP(16'h10DDD,4);
TASK_PP(16'h10DDE,4);
TASK_PP(16'h10DDF,4);
TASK_PP(16'h10DE0,4);
TASK_PP(16'h10DE1,4);
TASK_PP(16'h10DE2,4);
TASK_PP(16'h10DE3,4);
TASK_PP(16'h10DE4,4);
TASK_PP(16'h10DE5,4);
TASK_PP(16'h10DE6,4);
TASK_PP(16'h10DE7,4);
TASK_PP(16'h10DE8,4);
TASK_PP(16'h10DE9,4);
TASK_PP(16'h10DEA,4);
TASK_PP(16'h10DEB,4);
TASK_PP(16'h10DEC,4);
TASK_PP(16'h10DED,4);
TASK_PP(16'h10DEE,4);
TASK_PP(16'h10DEF,4);
TASK_PP(16'h10DF0,4);
TASK_PP(16'h10DF1,4);
TASK_PP(16'h10DF2,4);
TASK_PP(16'h10DF3,4);
TASK_PP(16'h10DF4,4);
TASK_PP(16'h10DF5,4);
TASK_PP(16'h10DF6,4);
TASK_PP(16'h10DF7,4);
TASK_PP(16'h10DF8,4);
TASK_PP(16'h10DF9,4);
TASK_PP(16'h10DFA,4);
TASK_PP(16'h10DFB,4);
TASK_PP(16'h10DFC,4);
TASK_PP(16'h10DFD,4);
TASK_PP(16'h10DFE,4);
TASK_PP(16'h10DFF,4);
TASK_PP(16'h10E00,4);
TASK_PP(16'h10E01,4);
TASK_PP(16'h10E02,4);
TASK_PP(16'h10E03,4);
TASK_PP(16'h10E04,4);
TASK_PP(16'h10E05,4);
TASK_PP(16'h10E06,4);
TASK_PP(16'h10E07,4);
TASK_PP(16'h10E08,4);
TASK_PP(16'h10E09,4);
TASK_PP(16'h10E0A,4);
TASK_PP(16'h10E0B,4);
TASK_PP(16'h10E0C,4);
TASK_PP(16'h10E0D,4);
TASK_PP(16'h10E0E,4);
TASK_PP(16'h10E0F,4);
TASK_PP(16'h10E10,4);
TASK_PP(16'h10E11,4);
TASK_PP(16'h10E12,4);
TASK_PP(16'h10E13,4);
TASK_PP(16'h10E14,4);
TASK_PP(16'h10E15,4);
TASK_PP(16'h10E16,4);
TASK_PP(16'h10E17,4);
TASK_PP(16'h10E18,4);
TASK_PP(16'h10E19,4);
TASK_PP(16'h10E1A,4);
TASK_PP(16'h10E1B,4);
TASK_PP(16'h10E1C,4);
TASK_PP(16'h10E1D,4);
TASK_PP(16'h10E1E,4);
TASK_PP(16'h10E1F,4);
TASK_PP(16'h10E20,4);
TASK_PP(16'h10E21,4);
TASK_PP(16'h10E22,4);
TASK_PP(16'h10E23,4);
TASK_PP(16'h10E24,4);
TASK_PP(16'h10E25,4);
TASK_PP(16'h10E26,4);
TASK_PP(16'h10E27,4);
TASK_PP(16'h10E28,4);
TASK_PP(16'h10E29,4);
TASK_PP(16'h10E2A,4);
TASK_PP(16'h10E2B,4);
TASK_PP(16'h10E2C,4);
TASK_PP(16'h10E2D,4);
TASK_PP(16'h10E2E,4);
TASK_PP(16'h10E2F,4);
TASK_PP(16'h10E30,4);
TASK_PP(16'h10E31,4);
TASK_PP(16'h10E32,4);
TASK_PP(16'h10E33,4);
TASK_PP(16'h10E34,4);
TASK_PP(16'h10E35,4);
TASK_PP(16'h10E36,4);
TASK_PP(16'h10E37,4);
TASK_PP(16'h10E38,4);
TASK_PP(16'h10E39,4);
TASK_PP(16'h10E3A,4);
TASK_PP(16'h10E3B,4);
TASK_PP(16'h10E3C,4);
TASK_PP(16'h10E3D,4);
TASK_PP(16'h10E3E,4);
TASK_PP(16'h10E3F,4);
TASK_PP(16'h10E40,4);
TASK_PP(16'h10E41,4);
TASK_PP(16'h10E42,4);
TASK_PP(16'h10E43,4);
TASK_PP(16'h10E44,4);
TASK_PP(16'h10E45,4);
TASK_PP(16'h10E46,4);
TASK_PP(16'h10E47,4);
TASK_PP(16'h10E48,4);
TASK_PP(16'h10E49,4);
TASK_PP(16'h10E4A,4);
TASK_PP(16'h10E4B,4);
TASK_PP(16'h10E4C,4);
TASK_PP(16'h10E4D,4);
TASK_PP(16'h10E4E,4);
TASK_PP(16'h10E4F,4);
TASK_PP(16'h10E50,4);
TASK_PP(16'h10E51,4);
TASK_PP(16'h10E52,4);
TASK_PP(16'h10E53,4);
TASK_PP(16'h10E54,4);
TASK_PP(16'h10E55,4);
TASK_PP(16'h10E56,4);
TASK_PP(16'h10E57,4);
TASK_PP(16'h10E58,4);
TASK_PP(16'h10E59,4);
TASK_PP(16'h10E5A,4);
TASK_PP(16'h10E5B,4);
TASK_PP(16'h10E5C,4);
TASK_PP(16'h10E5D,4);
TASK_PP(16'h10E5E,4);
TASK_PP(16'h10E5F,4);
TASK_PP(16'h10E60,4);
TASK_PP(16'h10E61,4);
TASK_PP(16'h10E62,4);
TASK_PP(16'h10E63,4);
TASK_PP(16'h10E64,4);
TASK_PP(16'h10E65,4);
TASK_PP(16'h10E66,4);
TASK_PP(16'h10E67,4);
TASK_PP(16'h10E68,4);
TASK_PP(16'h10E69,4);
TASK_PP(16'h10E6A,4);
TASK_PP(16'h10E6B,4);
TASK_PP(16'h10E6C,4);
TASK_PP(16'h10E6D,4);
TASK_PP(16'h10E6E,4);
TASK_PP(16'h10E6F,4);
TASK_PP(16'h10E70,4);
TASK_PP(16'h10E71,4);
TASK_PP(16'h10E72,4);
TASK_PP(16'h10E73,4);
TASK_PP(16'h10E74,4);
TASK_PP(16'h10E75,4);
TASK_PP(16'h10E76,4);
TASK_PP(16'h10E77,4);
TASK_PP(16'h10E78,4);
TASK_PP(16'h10E79,4);
TASK_PP(16'h10E7A,4);
TASK_PP(16'h10E7B,4);
TASK_PP(16'h10E7C,4);
TASK_PP(16'h10E7D,4);
TASK_PP(16'h10E7E,4);
TASK_PP(16'h10E7F,4);
TASK_PP(16'h10E80,4);
TASK_PP(16'h10E81,4);
TASK_PP(16'h10E82,4);
TASK_PP(16'h10E83,4);
TASK_PP(16'h10E84,4);
TASK_PP(16'h10E85,4);
TASK_PP(16'h10E86,4);
TASK_PP(16'h10E87,4);
TASK_PP(16'h10E88,4);
TASK_PP(16'h10E89,4);
TASK_PP(16'h10E8A,4);
TASK_PP(16'h10E8B,4);
TASK_PP(16'h10E8C,4);
TASK_PP(16'h10E8D,4);
TASK_PP(16'h10E8E,4);
TASK_PP(16'h10E8F,4);
TASK_PP(16'h10E90,4);
TASK_PP(16'h10E91,4);
TASK_PP(16'h10E92,4);
TASK_PP(16'h10E93,4);
TASK_PP(16'h10E94,4);
TASK_PP(16'h10E95,4);
TASK_PP(16'h10E96,4);
TASK_PP(16'h10E97,4);
TASK_PP(16'h10E98,4);
TASK_PP(16'h10E99,4);
TASK_PP(16'h10E9A,4);
TASK_PP(16'h10E9B,4);
TASK_PP(16'h10E9C,4);
TASK_PP(16'h10E9D,4);
TASK_PP(16'h10E9E,4);
TASK_PP(16'h10E9F,4);
TASK_PP(16'h10EA0,4);
TASK_PP(16'h10EA1,4);
TASK_PP(16'h10EA2,4);
TASK_PP(16'h10EA3,4);
TASK_PP(16'h10EA4,4);
TASK_PP(16'h10EA5,4);
TASK_PP(16'h10EA6,4);
TASK_PP(16'h10EA7,4);
TASK_PP(16'h10EA8,4);
TASK_PP(16'h10EA9,4);
TASK_PP(16'h10EAA,4);
TASK_PP(16'h10EAB,4);
TASK_PP(16'h10EAC,4);
TASK_PP(16'h10EAD,4);
TASK_PP(16'h10EAE,4);
TASK_PP(16'h10EAF,4);
TASK_PP(16'h10EB0,4);
TASK_PP(16'h10EB1,4);
TASK_PP(16'h10EB2,4);
TASK_PP(16'h10EB3,4);
TASK_PP(16'h10EB4,4);
TASK_PP(16'h10EB5,4);
TASK_PP(16'h10EB6,4);
TASK_PP(16'h10EB7,4);
TASK_PP(16'h10EB8,4);
TASK_PP(16'h10EB9,4);
TASK_PP(16'h10EBA,4);
TASK_PP(16'h10EBB,4);
TASK_PP(16'h10EBC,4);
TASK_PP(16'h10EBD,4);
TASK_PP(16'h10EBE,4);
TASK_PP(16'h10EBF,4);
TASK_PP(16'h10EC0,4);
TASK_PP(16'h10EC1,4);
TASK_PP(16'h10EC2,4);
TASK_PP(16'h10EC3,4);
TASK_PP(16'h10EC4,4);
TASK_PP(16'h10EC5,4);
TASK_PP(16'h10EC6,4);
TASK_PP(16'h10EC7,4);
TASK_PP(16'h10EC8,4);
TASK_PP(16'h10EC9,4);
TASK_PP(16'h10ECA,4);
TASK_PP(16'h10ECB,4);
TASK_PP(16'h10ECC,4);
TASK_PP(16'h10ECD,4);
TASK_PP(16'h10ECE,4);
TASK_PP(16'h10ECF,4);
TASK_PP(16'h10ED0,4);
TASK_PP(16'h10ED1,4);
TASK_PP(16'h10ED2,4);
TASK_PP(16'h10ED3,4);
TASK_PP(16'h10ED4,4);
TASK_PP(16'h10ED5,4);
TASK_PP(16'h10ED6,4);
TASK_PP(16'h10ED7,4);
TASK_PP(16'h10ED8,4);
TASK_PP(16'h10ED9,4);
TASK_PP(16'h10EDA,4);
TASK_PP(16'h10EDB,4);
TASK_PP(16'h10EDC,4);
TASK_PP(16'h10EDD,4);
TASK_PP(16'h10EDE,4);
TASK_PP(16'h10EDF,4);
TASK_PP(16'h10EE0,4);
TASK_PP(16'h10EE1,4);
TASK_PP(16'h10EE2,4);
TASK_PP(16'h10EE3,4);
TASK_PP(16'h10EE4,4);
TASK_PP(16'h10EE5,4);
TASK_PP(16'h10EE6,4);
TASK_PP(16'h10EE7,4);
TASK_PP(16'h10EE8,4);
TASK_PP(16'h10EE9,4);
TASK_PP(16'h10EEA,4);
TASK_PP(16'h10EEB,4);
TASK_PP(16'h10EEC,4);
TASK_PP(16'h10EED,4);
TASK_PP(16'h10EEE,4);
TASK_PP(16'h10EEF,4);
TASK_PP(16'h10EF0,4);
TASK_PP(16'h10EF1,4);
TASK_PP(16'h10EF2,4);
TASK_PP(16'h10EF3,4);
TASK_PP(16'h10EF4,4);
TASK_PP(16'h10EF5,4);
TASK_PP(16'h10EF6,4);
TASK_PP(16'h10EF7,4);
TASK_PP(16'h10EF8,4);
TASK_PP(16'h10EF9,4);
TASK_PP(16'h10EFA,4);
TASK_PP(16'h10EFB,4);
TASK_PP(16'h10EFC,4);
TASK_PP(16'h10EFD,4);
TASK_PP(16'h10EFE,4);
TASK_PP(16'h10EFF,4);
TASK_PP(16'h10F00,4);
TASK_PP(16'h10F01,4);
TASK_PP(16'h10F02,4);
TASK_PP(16'h10F03,4);
TASK_PP(16'h10F04,4);
TASK_PP(16'h10F05,4);
TASK_PP(16'h10F06,4);
TASK_PP(16'h10F07,4);
TASK_PP(16'h10F08,4);
TASK_PP(16'h10F09,4);
TASK_PP(16'h10F0A,4);
TASK_PP(16'h10F0B,4);
TASK_PP(16'h10F0C,4);
TASK_PP(16'h10F0D,4);
TASK_PP(16'h10F0E,4);
TASK_PP(16'h10F0F,4);
TASK_PP(16'h10F10,4);
TASK_PP(16'h10F11,4);
TASK_PP(16'h10F12,4);
TASK_PP(16'h10F13,4);
TASK_PP(16'h10F14,4);
TASK_PP(16'h10F15,4);
TASK_PP(16'h10F16,4);
TASK_PP(16'h10F17,4);
TASK_PP(16'h10F18,4);
TASK_PP(16'h10F19,4);
TASK_PP(16'h10F1A,4);
TASK_PP(16'h10F1B,4);
TASK_PP(16'h10F1C,4);
TASK_PP(16'h10F1D,4);
TASK_PP(16'h10F1E,4);
TASK_PP(16'h10F1F,4);
TASK_PP(16'h10F20,4);
TASK_PP(16'h10F21,4);
TASK_PP(16'h10F22,4);
TASK_PP(16'h10F23,4);
TASK_PP(16'h10F24,4);
TASK_PP(16'h10F25,4);
TASK_PP(16'h10F26,4);
TASK_PP(16'h10F27,4);
TASK_PP(16'h10F28,4);
TASK_PP(16'h10F29,4);
TASK_PP(16'h10F2A,4);
TASK_PP(16'h10F2B,4);
TASK_PP(16'h10F2C,4);
TASK_PP(16'h10F2D,4);
TASK_PP(16'h10F2E,4);
TASK_PP(16'h10F2F,4);
TASK_PP(16'h10F30,4);
TASK_PP(16'h10F31,4);
TASK_PP(16'h10F32,4);
TASK_PP(16'h10F33,4);
TASK_PP(16'h10F34,4);
TASK_PP(16'h10F35,4);
TASK_PP(16'h10F36,4);
TASK_PP(16'h10F37,4);
TASK_PP(16'h10F38,4);
TASK_PP(16'h10F39,4);
TASK_PP(16'h10F3A,4);
TASK_PP(16'h10F3B,4);
TASK_PP(16'h10F3C,4);
TASK_PP(16'h10F3D,4);
TASK_PP(16'h10F3E,4);
TASK_PP(16'h10F3F,4);
TASK_PP(16'h10F40,4);
TASK_PP(16'h10F41,4);
TASK_PP(16'h10F42,4);
TASK_PP(16'h10F43,4);
TASK_PP(16'h10F44,4);
TASK_PP(16'h10F45,4);
TASK_PP(16'h10F46,4);
TASK_PP(16'h10F47,4);
TASK_PP(16'h10F48,4);
TASK_PP(16'h10F49,4);
TASK_PP(16'h10F4A,4);
TASK_PP(16'h10F4B,4);
TASK_PP(16'h10F4C,4);
TASK_PP(16'h10F4D,4);
TASK_PP(16'h10F4E,4);
TASK_PP(16'h10F4F,4);
TASK_PP(16'h10F50,4);
TASK_PP(16'h10F51,4);
TASK_PP(16'h10F52,4);
TASK_PP(16'h10F53,4);
TASK_PP(16'h10F54,4);
TASK_PP(16'h10F55,4);
TASK_PP(16'h10F56,4);
TASK_PP(16'h10F57,4);
TASK_PP(16'h10F58,4);
TASK_PP(16'h10F59,4);
TASK_PP(16'h10F5A,4);
TASK_PP(16'h10F5B,4);
TASK_PP(16'h10F5C,4);
TASK_PP(16'h10F5D,4);
TASK_PP(16'h10F5E,4);
TASK_PP(16'h10F5F,4);
TASK_PP(16'h10F60,4);
TASK_PP(16'h10F61,4);
TASK_PP(16'h10F62,4);
TASK_PP(16'h10F63,4);
TASK_PP(16'h10F64,4);
TASK_PP(16'h10F65,4);
TASK_PP(16'h10F66,4);
TASK_PP(16'h10F67,4);
TASK_PP(16'h10F68,4);
TASK_PP(16'h10F69,4);
TASK_PP(16'h10F6A,4);
TASK_PP(16'h10F6B,4);
TASK_PP(16'h10F6C,4);
TASK_PP(16'h10F6D,4);
TASK_PP(16'h10F6E,4);
TASK_PP(16'h10F6F,4);
TASK_PP(16'h10F70,4);
TASK_PP(16'h10F71,4);
TASK_PP(16'h10F72,4);
TASK_PP(16'h10F73,4);
TASK_PP(16'h10F74,4);
TASK_PP(16'h10F75,4);
TASK_PP(16'h10F76,4);
TASK_PP(16'h10F77,4);
TASK_PP(16'h10F78,4);
TASK_PP(16'h10F79,4);
TASK_PP(16'h10F7A,4);
TASK_PP(16'h10F7B,4);
TASK_PP(16'h10F7C,4);
TASK_PP(16'h10F7D,4);
TASK_PP(16'h10F7E,4);
TASK_PP(16'h10F7F,4);
TASK_PP(16'h10F80,4);
TASK_PP(16'h10F81,4);
TASK_PP(16'h10F82,4);
TASK_PP(16'h10F83,4);
TASK_PP(16'h10F84,4);
TASK_PP(16'h10F85,4);
TASK_PP(16'h10F86,4);
TASK_PP(16'h10F87,4);
TASK_PP(16'h10F88,4);
TASK_PP(16'h10F89,4);
TASK_PP(16'h10F8A,4);
TASK_PP(16'h10F8B,4);
TASK_PP(16'h10F8C,4);
TASK_PP(16'h10F8D,4);
TASK_PP(16'h10F8E,4);
TASK_PP(16'h10F8F,4);
TASK_PP(16'h10F90,4);
TASK_PP(16'h10F91,4);
TASK_PP(16'h10F92,4);
TASK_PP(16'h10F93,4);
TASK_PP(16'h10F94,4);
TASK_PP(16'h10F95,4);
TASK_PP(16'h10F96,4);
TASK_PP(16'h10F97,4);
TASK_PP(16'h10F98,4);
TASK_PP(16'h10F99,4);
TASK_PP(16'h10F9A,4);
TASK_PP(16'h10F9B,4);
TASK_PP(16'h10F9C,4);
TASK_PP(16'h10F9D,4);
TASK_PP(16'h10F9E,4);
TASK_PP(16'h10F9F,4);
TASK_PP(16'h10FA0,4);
TASK_PP(16'h10FA1,4);
TASK_PP(16'h10FA2,4);
TASK_PP(16'h10FA3,4);
TASK_PP(16'h10FA4,4);
TASK_PP(16'h10FA5,4);
TASK_PP(16'h10FA6,4);
TASK_PP(16'h10FA7,4);
TASK_PP(16'h10FA8,4);
TASK_PP(16'h10FA9,4);
TASK_PP(16'h10FAA,4);
TASK_PP(16'h10FAB,4);
TASK_PP(16'h10FAC,4);
TASK_PP(16'h10FAD,4);
TASK_PP(16'h10FAE,4);
TASK_PP(16'h10FAF,4);
TASK_PP(16'h10FB0,4);
TASK_PP(16'h10FB1,4);
TASK_PP(16'h10FB2,4);
TASK_PP(16'h10FB3,4);
TASK_PP(16'h10FB4,4);
TASK_PP(16'h10FB5,4);
TASK_PP(16'h10FB6,4);
TASK_PP(16'h10FB7,4);
TASK_PP(16'h10FB8,4);
TASK_PP(16'h10FB9,4);
TASK_PP(16'h10FBA,4);
TASK_PP(16'h10FBB,4);
TASK_PP(16'h10FBC,4);
TASK_PP(16'h10FBD,4);
TASK_PP(16'h10FBE,4);
TASK_PP(16'h10FBF,4);
TASK_PP(16'h10FC0,4);
TASK_PP(16'h10FC1,4);
TASK_PP(16'h10FC2,4);
TASK_PP(16'h10FC3,4);
TASK_PP(16'h10FC4,4);
TASK_PP(16'h10FC5,4);
TASK_PP(16'h10FC6,4);
TASK_PP(16'h10FC7,4);
TASK_PP(16'h10FC8,4);
TASK_PP(16'h10FC9,4);
TASK_PP(16'h10FCA,4);
TASK_PP(16'h10FCB,4);
TASK_PP(16'h10FCC,4);
TASK_PP(16'h10FCD,4);
TASK_PP(16'h10FCE,4);
TASK_PP(16'h10FCF,4);
TASK_PP(16'h10FD0,4);
TASK_PP(16'h10FD1,4);
TASK_PP(16'h10FD2,4);
TASK_PP(16'h10FD3,4);
TASK_PP(16'h10FD4,4);
TASK_PP(16'h10FD5,4);
TASK_PP(16'h10FD6,4);
TASK_PP(16'h10FD7,4);
TASK_PP(16'h10FD8,4);
TASK_PP(16'h10FD9,4);
TASK_PP(16'h10FDA,4);
TASK_PP(16'h10FDB,4);
TASK_PP(16'h10FDC,4);
TASK_PP(16'h10FDD,4);
TASK_PP(16'h10FDE,4);
TASK_PP(16'h10FDF,4);
TASK_PP(16'h10FE0,4);
TASK_PP(16'h10FE1,4);
TASK_PP(16'h10FE2,4);
TASK_PP(16'h10FE3,4);
TASK_PP(16'h10FE4,4);
TASK_PP(16'h10FE5,4);
TASK_PP(16'h10FE6,4);
TASK_PP(16'h10FE7,4);
TASK_PP(16'h10FE8,4);
TASK_PP(16'h10FE9,4);
TASK_PP(16'h10FEA,4);
TASK_PP(16'h10FEB,4);
TASK_PP(16'h10FEC,4);
TASK_PP(16'h10FED,4);
TASK_PP(16'h10FEE,4);
TASK_PP(16'h10FEF,4);
TASK_PP(16'h10FF0,4);
TASK_PP(16'h10FF1,4);
TASK_PP(16'h10FF2,4);
TASK_PP(16'h10FF3,4);
TASK_PP(16'h10FF4,4);
TASK_PP(16'h10FF5,4);
TASK_PP(16'h10FF6,4);
TASK_PP(16'h10FF7,4);
TASK_PP(16'h10FF8,4);
TASK_PP(16'h10FF9,4);
TASK_PP(16'h10FFA,4);
TASK_PP(16'h10FFB,4);
TASK_PP(16'h10FFC,4);
TASK_PP(16'h10FFD,4);
TASK_PP(16'h10FFE,4);
TASK_PP(16'h10FFF,4);
TASK_PP(16'h11000,4);
TASK_PP(16'h11001,4);
TASK_PP(16'h11002,4);
TASK_PP(16'h11003,4);
TASK_PP(16'h11004,4);
TASK_PP(16'h11005,4);
TASK_PP(16'h11006,4);
TASK_PP(16'h11007,4);
TASK_PP(16'h11008,4);
TASK_PP(16'h11009,4);
TASK_PP(16'h1100A,4);
TASK_PP(16'h1100B,4);
TASK_PP(16'h1100C,4);
TASK_PP(16'h1100D,4);
TASK_PP(16'h1100E,4);
TASK_PP(16'h1100F,4);
TASK_PP(16'h11010,4);
TASK_PP(16'h11011,4);
TASK_PP(16'h11012,4);
TASK_PP(16'h11013,4);
TASK_PP(16'h11014,4);
TASK_PP(16'h11015,4);
TASK_PP(16'h11016,4);
TASK_PP(16'h11017,4);
TASK_PP(16'h11018,4);
TASK_PP(16'h11019,4);
TASK_PP(16'h1101A,4);
TASK_PP(16'h1101B,4);
TASK_PP(16'h1101C,4);
TASK_PP(16'h1101D,4);
TASK_PP(16'h1101E,4);
TASK_PP(16'h1101F,4);
TASK_PP(16'h11020,4);
TASK_PP(16'h11021,4);
TASK_PP(16'h11022,4);
TASK_PP(16'h11023,4);
TASK_PP(16'h11024,4);
TASK_PP(16'h11025,4);
TASK_PP(16'h11026,4);
TASK_PP(16'h11027,4);
TASK_PP(16'h11028,4);
TASK_PP(16'h11029,4);
TASK_PP(16'h1102A,4);
TASK_PP(16'h1102B,4);
TASK_PP(16'h1102C,4);
TASK_PP(16'h1102D,4);
TASK_PP(16'h1102E,4);
TASK_PP(16'h1102F,4);
TASK_PP(16'h11030,4);
TASK_PP(16'h11031,4);
TASK_PP(16'h11032,4);
TASK_PP(16'h11033,4);
TASK_PP(16'h11034,4);
TASK_PP(16'h11035,4);
TASK_PP(16'h11036,4);
TASK_PP(16'h11037,4);
TASK_PP(16'h11038,4);
TASK_PP(16'h11039,4);
TASK_PP(16'h1103A,4);
TASK_PP(16'h1103B,4);
TASK_PP(16'h1103C,4);
TASK_PP(16'h1103D,4);
TASK_PP(16'h1103E,4);
TASK_PP(16'h1103F,4);
TASK_PP(16'h11040,4);
TASK_PP(16'h11041,4);
TASK_PP(16'h11042,4);
TASK_PP(16'h11043,4);
TASK_PP(16'h11044,4);
TASK_PP(16'h11045,4);
TASK_PP(16'h11046,4);
TASK_PP(16'h11047,4);
TASK_PP(16'h11048,4);
TASK_PP(16'h11049,4);
TASK_PP(16'h1104A,4);
TASK_PP(16'h1104B,4);
TASK_PP(16'h1104C,4);
TASK_PP(16'h1104D,4);
TASK_PP(16'h1104E,4);
TASK_PP(16'h1104F,4);
TASK_PP(16'h11050,4);
TASK_PP(16'h11051,4);
TASK_PP(16'h11052,4);
TASK_PP(16'h11053,4);
TASK_PP(16'h11054,4);
TASK_PP(16'h11055,4);
TASK_PP(16'h11056,4);
TASK_PP(16'h11057,4);
TASK_PP(16'h11058,4);
TASK_PP(16'h11059,4);
TASK_PP(16'h1105A,4);
TASK_PP(16'h1105B,4);
TASK_PP(16'h1105C,4);
TASK_PP(16'h1105D,4);
TASK_PP(16'h1105E,4);
TASK_PP(16'h1105F,4);
TASK_PP(16'h11060,4);
TASK_PP(16'h11061,4);
TASK_PP(16'h11062,4);
TASK_PP(16'h11063,4);
TASK_PP(16'h11064,4);
TASK_PP(16'h11065,4);
TASK_PP(16'h11066,4);
TASK_PP(16'h11067,4);
TASK_PP(16'h11068,4);
TASK_PP(16'h11069,4);
TASK_PP(16'h1106A,4);
TASK_PP(16'h1106B,4);
TASK_PP(16'h1106C,4);
TASK_PP(16'h1106D,4);
TASK_PP(16'h1106E,4);
TASK_PP(16'h1106F,4);
TASK_PP(16'h11070,4);
TASK_PP(16'h11071,4);
TASK_PP(16'h11072,4);
TASK_PP(16'h11073,4);
TASK_PP(16'h11074,4);
TASK_PP(16'h11075,4);
TASK_PP(16'h11076,4);
TASK_PP(16'h11077,4);
TASK_PP(16'h11078,4);
TASK_PP(16'h11079,4);
TASK_PP(16'h1107A,4);
TASK_PP(16'h1107B,4);
TASK_PP(16'h1107C,4);
TASK_PP(16'h1107D,4);
TASK_PP(16'h1107E,4);
TASK_PP(16'h1107F,4);
TASK_PP(16'h11080,4);
TASK_PP(16'h11081,4);
TASK_PP(16'h11082,4);
TASK_PP(16'h11083,4);
TASK_PP(16'h11084,4);
TASK_PP(16'h11085,4);
TASK_PP(16'h11086,4);
TASK_PP(16'h11087,4);
TASK_PP(16'h11088,4);
TASK_PP(16'h11089,4);
TASK_PP(16'h1108A,4);
TASK_PP(16'h1108B,4);
TASK_PP(16'h1108C,4);
TASK_PP(16'h1108D,4);
TASK_PP(16'h1108E,4);
TASK_PP(16'h1108F,4);
TASK_PP(16'h11090,4);
TASK_PP(16'h11091,4);
TASK_PP(16'h11092,4);
TASK_PP(16'h11093,4);
TASK_PP(16'h11094,4);
TASK_PP(16'h11095,4);
TASK_PP(16'h11096,4);
TASK_PP(16'h11097,4);
TASK_PP(16'h11098,4);
TASK_PP(16'h11099,4);
TASK_PP(16'h1109A,4);
TASK_PP(16'h1109B,4);
TASK_PP(16'h1109C,4);
TASK_PP(16'h1109D,4);
TASK_PP(16'h1109E,4);
TASK_PP(16'h1109F,4);
TASK_PP(16'h110A0,4);
TASK_PP(16'h110A1,4);
TASK_PP(16'h110A2,4);
TASK_PP(16'h110A3,4);
TASK_PP(16'h110A4,4);
TASK_PP(16'h110A5,4);
TASK_PP(16'h110A6,4);
TASK_PP(16'h110A7,4);
TASK_PP(16'h110A8,4);
TASK_PP(16'h110A9,4);
TASK_PP(16'h110AA,4);
TASK_PP(16'h110AB,4);
TASK_PP(16'h110AC,4);
TASK_PP(16'h110AD,4);
TASK_PP(16'h110AE,4);
TASK_PP(16'h110AF,4);
TASK_PP(16'h110B0,4);
TASK_PP(16'h110B1,4);
TASK_PP(16'h110B2,4);
TASK_PP(16'h110B3,4);
TASK_PP(16'h110B4,4);
TASK_PP(16'h110B5,4);
TASK_PP(16'h110B6,4);
TASK_PP(16'h110B7,4);
TASK_PP(16'h110B8,4);
TASK_PP(16'h110B9,4);
TASK_PP(16'h110BA,4);
TASK_PP(16'h110BB,4);
TASK_PP(16'h110BC,4);
TASK_PP(16'h110BD,4);
TASK_PP(16'h110BE,4);
TASK_PP(16'h110BF,4);
TASK_PP(16'h110C0,4);
TASK_PP(16'h110C1,4);
TASK_PP(16'h110C2,4);
TASK_PP(16'h110C3,4);
TASK_PP(16'h110C4,4);
TASK_PP(16'h110C5,4);
TASK_PP(16'h110C6,4);
TASK_PP(16'h110C7,4);
TASK_PP(16'h110C8,4);
TASK_PP(16'h110C9,4);
TASK_PP(16'h110CA,4);
TASK_PP(16'h110CB,4);
TASK_PP(16'h110CC,4);
TASK_PP(16'h110CD,4);
TASK_PP(16'h110CE,4);
TASK_PP(16'h110CF,4);
TASK_PP(16'h110D0,4);
TASK_PP(16'h110D1,4);
TASK_PP(16'h110D2,4);
TASK_PP(16'h110D3,4);
TASK_PP(16'h110D4,4);
TASK_PP(16'h110D5,4);
TASK_PP(16'h110D6,4);
TASK_PP(16'h110D7,4);
TASK_PP(16'h110D8,4);
TASK_PP(16'h110D9,4);
TASK_PP(16'h110DA,4);
TASK_PP(16'h110DB,4);
TASK_PP(16'h110DC,4);
TASK_PP(16'h110DD,4);
TASK_PP(16'h110DE,4);
TASK_PP(16'h110DF,4);
TASK_PP(16'h110E0,4);
TASK_PP(16'h110E1,4);
TASK_PP(16'h110E2,4);
TASK_PP(16'h110E3,4);
TASK_PP(16'h110E4,4);
TASK_PP(16'h110E5,4);
TASK_PP(16'h110E6,4);
TASK_PP(16'h110E7,4);
TASK_PP(16'h110E8,4);
TASK_PP(16'h110E9,4);
TASK_PP(16'h110EA,4);
TASK_PP(16'h110EB,4);
TASK_PP(16'h110EC,4);
TASK_PP(16'h110ED,4);
TASK_PP(16'h110EE,4);
TASK_PP(16'h110EF,4);
TASK_PP(16'h110F0,4);
TASK_PP(16'h110F1,4);
TASK_PP(16'h110F2,4);
TASK_PP(16'h110F3,4);
TASK_PP(16'h110F4,4);
TASK_PP(16'h110F5,4);
TASK_PP(16'h110F6,4);
TASK_PP(16'h110F7,4);
TASK_PP(16'h110F8,4);
TASK_PP(16'h110F9,4);
TASK_PP(16'h110FA,4);
TASK_PP(16'h110FB,4);
TASK_PP(16'h110FC,4);
TASK_PP(16'h110FD,4);
TASK_PP(16'h110FE,4);
TASK_PP(16'h110FF,4);
TASK_PP(16'h11100,4);
TASK_PP(16'h11101,4);
TASK_PP(16'h11102,4);
TASK_PP(16'h11103,4);
TASK_PP(16'h11104,4);
TASK_PP(16'h11105,4);
TASK_PP(16'h11106,4);
TASK_PP(16'h11107,4);
TASK_PP(16'h11108,4);
TASK_PP(16'h11109,4);
TASK_PP(16'h1110A,4);
TASK_PP(16'h1110B,4);
TASK_PP(16'h1110C,4);
TASK_PP(16'h1110D,4);
TASK_PP(16'h1110E,4);
TASK_PP(16'h1110F,4);
TASK_PP(16'h11110,4);
TASK_PP(16'h11111,4);
TASK_PP(16'h11112,4);
TASK_PP(16'h11113,4);
TASK_PP(16'h11114,4);
TASK_PP(16'h11115,4);
TASK_PP(16'h11116,4);
TASK_PP(16'h11117,4);
TASK_PP(16'h11118,4);
TASK_PP(16'h11119,4);
TASK_PP(16'h1111A,4);
TASK_PP(16'h1111B,4);
TASK_PP(16'h1111C,4);
TASK_PP(16'h1111D,4);
TASK_PP(16'h1111E,4);
TASK_PP(16'h1111F,4);
TASK_PP(16'h11120,4);
TASK_PP(16'h11121,4);
TASK_PP(16'h11122,4);
TASK_PP(16'h11123,4);
TASK_PP(16'h11124,4);
TASK_PP(16'h11125,4);
TASK_PP(16'h11126,4);
TASK_PP(16'h11127,4);
TASK_PP(16'h11128,4);
TASK_PP(16'h11129,4);
TASK_PP(16'h1112A,4);
TASK_PP(16'h1112B,4);
TASK_PP(16'h1112C,4);
TASK_PP(16'h1112D,4);
TASK_PP(16'h1112E,4);
TASK_PP(16'h1112F,4);
TASK_PP(16'h11130,4);
TASK_PP(16'h11131,4);
TASK_PP(16'h11132,4);
TASK_PP(16'h11133,4);
TASK_PP(16'h11134,4);
TASK_PP(16'h11135,4);
TASK_PP(16'h11136,4);
TASK_PP(16'h11137,4);
TASK_PP(16'h11138,4);
TASK_PP(16'h11139,4);
TASK_PP(16'h1113A,4);
TASK_PP(16'h1113B,4);
TASK_PP(16'h1113C,4);
TASK_PP(16'h1113D,4);
TASK_PP(16'h1113E,4);
TASK_PP(16'h1113F,4);
TASK_PP(16'h11140,4);
TASK_PP(16'h11141,4);
TASK_PP(16'h11142,4);
TASK_PP(16'h11143,4);
TASK_PP(16'h11144,4);
TASK_PP(16'h11145,4);
TASK_PP(16'h11146,4);
TASK_PP(16'h11147,4);
TASK_PP(16'h11148,4);
TASK_PP(16'h11149,4);
TASK_PP(16'h1114A,4);
TASK_PP(16'h1114B,4);
TASK_PP(16'h1114C,4);
TASK_PP(16'h1114D,4);
TASK_PP(16'h1114E,4);
TASK_PP(16'h1114F,4);
TASK_PP(16'h11150,4);
TASK_PP(16'h11151,4);
TASK_PP(16'h11152,4);
TASK_PP(16'h11153,4);
TASK_PP(16'h11154,4);
TASK_PP(16'h11155,4);
TASK_PP(16'h11156,4);
TASK_PP(16'h11157,4);
TASK_PP(16'h11158,4);
TASK_PP(16'h11159,4);
TASK_PP(16'h1115A,4);
TASK_PP(16'h1115B,4);
TASK_PP(16'h1115C,4);
TASK_PP(16'h1115D,4);
TASK_PP(16'h1115E,4);
TASK_PP(16'h1115F,4);
TASK_PP(16'h11160,4);
TASK_PP(16'h11161,4);
TASK_PP(16'h11162,4);
TASK_PP(16'h11163,4);
TASK_PP(16'h11164,4);
TASK_PP(16'h11165,4);
TASK_PP(16'h11166,4);
TASK_PP(16'h11167,4);
TASK_PP(16'h11168,4);
TASK_PP(16'h11169,4);
TASK_PP(16'h1116A,4);
TASK_PP(16'h1116B,4);
TASK_PP(16'h1116C,4);
TASK_PP(16'h1116D,4);
TASK_PP(16'h1116E,4);
TASK_PP(16'h1116F,4);
TASK_PP(16'h11170,4);
TASK_PP(16'h11171,4);
TASK_PP(16'h11172,4);
TASK_PP(16'h11173,4);
TASK_PP(16'h11174,4);
TASK_PP(16'h11175,4);
TASK_PP(16'h11176,4);
TASK_PP(16'h11177,4);
TASK_PP(16'h11178,4);
TASK_PP(16'h11179,4);
TASK_PP(16'h1117A,4);
TASK_PP(16'h1117B,4);
TASK_PP(16'h1117C,4);
TASK_PP(16'h1117D,4);
TASK_PP(16'h1117E,4);
TASK_PP(16'h1117F,4);
TASK_PP(16'h11180,4);
TASK_PP(16'h11181,4);
TASK_PP(16'h11182,4);
TASK_PP(16'h11183,4);
TASK_PP(16'h11184,4);
TASK_PP(16'h11185,4);
TASK_PP(16'h11186,4);
TASK_PP(16'h11187,4);
TASK_PP(16'h11188,4);
TASK_PP(16'h11189,4);
TASK_PP(16'h1118A,4);
TASK_PP(16'h1118B,4);
TASK_PP(16'h1118C,4);
TASK_PP(16'h1118D,4);
TASK_PP(16'h1118E,4);
TASK_PP(16'h1118F,4);
TASK_PP(16'h11190,4);
TASK_PP(16'h11191,4);
TASK_PP(16'h11192,4);
TASK_PP(16'h11193,4);
TASK_PP(16'h11194,4);
TASK_PP(16'h11195,4);
TASK_PP(16'h11196,4);
TASK_PP(16'h11197,4);
TASK_PP(16'h11198,4);
TASK_PP(16'h11199,4);
TASK_PP(16'h1119A,4);
TASK_PP(16'h1119B,4);
TASK_PP(16'h1119C,4);
TASK_PP(16'h1119D,4);
TASK_PP(16'h1119E,4);
TASK_PP(16'h1119F,4);
TASK_PP(16'h111A0,4);
TASK_PP(16'h111A1,4);
TASK_PP(16'h111A2,4);
TASK_PP(16'h111A3,4);
TASK_PP(16'h111A4,4);
TASK_PP(16'h111A5,4);
TASK_PP(16'h111A6,4);
TASK_PP(16'h111A7,4);
TASK_PP(16'h111A8,4);
TASK_PP(16'h111A9,4);
TASK_PP(16'h111AA,4);
TASK_PP(16'h111AB,4);
TASK_PP(16'h111AC,4);
TASK_PP(16'h111AD,4);
TASK_PP(16'h111AE,4);
TASK_PP(16'h111AF,4);
TASK_PP(16'h111B0,4);
TASK_PP(16'h111B1,4);
TASK_PP(16'h111B2,4);
TASK_PP(16'h111B3,4);
TASK_PP(16'h111B4,4);
TASK_PP(16'h111B5,4);
TASK_PP(16'h111B6,4);
TASK_PP(16'h111B7,4);
TASK_PP(16'h111B8,4);
TASK_PP(16'h111B9,4);
TASK_PP(16'h111BA,4);
TASK_PP(16'h111BB,4);
TASK_PP(16'h111BC,4);
TASK_PP(16'h111BD,4);
TASK_PP(16'h111BE,4);
TASK_PP(16'h111BF,4);
TASK_PP(16'h111C0,4);
TASK_PP(16'h111C1,4);
TASK_PP(16'h111C2,4);
TASK_PP(16'h111C3,4);
TASK_PP(16'h111C4,4);
TASK_PP(16'h111C5,4);
TASK_PP(16'h111C6,4);
TASK_PP(16'h111C7,4);
TASK_PP(16'h111C8,4);
TASK_PP(16'h111C9,4);
TASK_PP(16'h111CA,4);
TASK_PP(16'h111CB,4);
TASK_PP(16'h111CC,4);
TASK_PP(16'h111CD,4);
TASK_PP(16'h111CE,4);
TASK_PP(16'h111CF,4);
TASK_PP(16'h111D0,4);
TASK_PP(16'h111D1,4);
TASK_PP(16'h111D2,4);
TASK_PP(16'h111D3,4);
TASK_PP(16'h111D4,4);
TASK_PP(16'h111D5,4);
TASK_PP(16'h111D6,4);
TASK_PP(16'h111D7,4);
TASK_PP(16'h111D8,4);
TASK_PP(16'h111D9,4);
TASK_PP(16'h111DA,4);
TASK_PP(16'h111DB,4);
TASK_PP(16'h111DC,4);
TASK_PP(16'h111DD,4);
TASK_PP(16'h111DE,4);
TASK_PP(16'h111DF,4);
TASK_PP(16'h111E0,4);
TASK_PP(16'h111E1,4);
TASK_PP(16'h111E2,4);
TASK_PP(16'h111E3,4);
TASK_PP(16'h111E4,4);
TASK_PP(16'h111E5,4);
TASK_PP(16'h111E6,4);
TASK_PP(16'h111E7,4);
TASK_PP(16'h111E8,4);
TASK_PP(16'h111E9,4);
TASK_PP(16'h111EA,4);
TASK_PP(16'h111EB,4);
TASK_PP(16'h111EC,4);
TASK_PP(16'h111ED,4);
TASK_PP(16'h111EE,4);
TASK_PP(16'h111EF,4);
TASK_PP(16'h111F0,4);
TASK_PP(16'h111F1,4);
TASK_PP(16'h111F2,4);
TASK_PP(16'h111F3,4);
TASK_PP(16'h111F4,4);
TASK_PP(16'h111F5,4);
TASK_PP(16'h111F6,4);
TASK_PP(16'h111F7,4);
TASK_PP(16'h111F8,4);
TASK_PP(16'h111F9,4);
TASK_PP(16'h111FA,4);
TASK_PP(16'h111FB,4);
TASK_PP(16'h111FC,4);
TASK_PP(16'h111FD,4);
TASK_PP(16'h111FE,4);
TASK_PP(16'h111FF,4);
TASK_PP(16'h11200,4);
TASK_PP(16'h11201,4);
TASK_PP(16'h11202,4);
TASK_PP(16'h11203,4);
TASK_PP(16'h11204,4);
TASK_PP(16'h11205,4);
TASK_PP(16'h11206,4);
TASK_PP(16'h11207,4);
TASK_PP(16'h11208,4);
TASK_PP(16'h11209,4);
TASK_PP(16'h1120A,4);
TASK_PP(16'h1120B,4);
TASK_PP(16'h1120C,4);
TASK_PP(16'h1120D,4);
TASK_PP(16'h1120E,4);
TASK_PP(16'h1120F,4);
TASK_PP(16'h11210,4);
TASK_PP(16'h11211,4);
TASK_PP(16'h11212,4);
TASK_PP(16'h11213,4);
TASK_PP(16'h11214,4);
TASK_PP(16'h11215,4);
TASK_PP(16'h11216,4);
TASK_PP(16'h11217,4);
TASK_PP(16'h11218,4);
TASK_PP(16'h11219,4);
TASK_PP(16'h1121A,4);
TASK_PP(16'h1121B,4);
TASK_PP(16'h1121C,4);
TASK_PP(16'h1121D,4);
TASK_PP(16'h1121E,4);
TASK_PP(16'h1121F,4);
TASK_PP(16'h11220,4);
TASK_PP(16'h11221,4);
TASK_PP(16'h11222,4);
TASK_PP(16'h11223,4);
TASK_PP(16'h11224,4);
TASK_PP(16'h11225,4);
TASK_PP(16'h11226,4);
TASK_PP(16'h11227,4);
TASK_PP(16'h11228,4);
TASK_PP(16'h11229,4);
TASK_PP(16'h1122A,4);
TASK_PP(16'h1122B,4);
TASK_PP(16'h1122C,4);
TASK_PP(16'h1122D,4);
TASK_PP(16'h1122E,4);
TASK_PP(16'h1122F,4);
TASK_PP(16'h11230,4);
TASK_PP(16'h11231,4);
TASK_PP(16'h11232,4);
TASK_PP(16'h11233,4);
TASK_PP(16'h11234,4);
TASK_PP(16'h11235,4);
TASK_PP(16'h11236,4);
TASK_PP(16'h11237,4);
TASK_PP(16'h11238,4);
TASK_PP(16'h11239,4);
TASK_PP(16'h1123A,4);
TASK_PP(16'h1123B,4);
TASK_PP(16'h1123C,4);
TASK_PP(16'h1123D,4);
TASK_PP(16'h1123E,4);
TASK_PP(16'h1123F,4);
TASK_PP(16'h11240,4);
TASK_PP(16'h11241,4);
TASK_PP(16'h11242,4);
TASK_PP(16'h11243,4);
TASK_PP(16'h11244,4);
TASK_PP(16'h11245,4);
TASK_PP(16'h11246,4);
TASK_PP(16'h11247,4);
TASK_PP(16'h11248,4);
TASK_PP(16'h11249,4);
TASK_PP(16'h1124A,4);
TASK_PP(16'h1124B,4);
TASK_PP(16'h1124C,4);
TASK_PP(16'h1124D,4);
TASK_PP(16'h1124E,4);
TASK_PP(16'h1124F,4);
TASK_PP(16'h11250,4);
TASK_PP(16'h11251,4);
TASK_PP(16'h11252,4);
TASK_PP(16'h11253,4);
TASK_PP(16'h11254,4);
TASK_PP(16'h11255,4);
TASK_PP(16'h11256,4);
TASK_PP(16'h11257,4);
TASK_PP(16'h11258,4);
TASK_PP(16'h11259,4);
TASK_PP(16'h1125A,4);
TASK_PP(16'h1125B,4);
TASK_PP(16'h1125C,4);
TASK_PP(16'h1125D,4);
TASK_PP(16'h1125E,4);
TASK_PP(16'h1125F,4);
TASK_PP(16'h11260,4);
TASK_PP(16'h11261,4);
TASK_PP(16'h11262,4);
TASK_PP(16'h11263,4);
TASK_PP(16'h11264,4);
TASK_PP(16'h11265,4);
TASK_PP(16'h11266,4);
TASK_PP(16'h11267,4);
TASK_PP(16'h11268,4);
TASK_PP(16'h11269,4);
TASK_PP(16'h1126A,4);
TASK_PP(16'h1126B,4);
TASK_PP(16'h1126C,4);
TASK_PP(16'h1126D,4);
TASK_PP(16'h1126E,4);
TASK_PP(16'h1126F,4);
TASK_PP(16'h11270,4);
TASK_PP(16'h11271,4);
TASK_PP(16'h11272,4);
TASK_PP(16'h11273,4);
TASK_PP(16'h11274,4);
TASK_PP(16'h11275,4);
TASK_PP(16'h11276,4);
TASK_PP(16'h11277,4);
TASK_PP(16'h11278,4);
TASK_PP(16'h11279,4);
TASK_PP(16'h1127A,4);
TASK_PP(16'h1127B,4);
TASK_PP(16'h1127C,4);
TASK_PP(16'h1127D,4);
TASK_PP(16'h1127E,4);
TASK_PP(16'h1127F,4);
TASK_PP(16'h11280,4);
TASK_PP(16'h11281,4);
TASK_PP(16'h11282,4);
TASK_PP(16'h11283,4);
TASK_PP(16'h11284,4);
TASK_PP(16'h11285,4);
TASK_PP(16'h11286,4);
TASK_PP(16'h11287,4);
TASK_PP(16'h11288,4);
TASK_PP(16'h11289,4);
TASK_PP(16'h1128A,4);
TASK_PP(16'h1128B,4);
TASK_PP(16'h1128C,4);
TASK_PP(16'h1128D,4);
TASK_PP(16'h1128E,4);
TASK_PP(16'h1128F,4);
TASK_PP(16'h11290,4);
TASK_PP(16'h11291,4);
TASK_PP(16'h11292,4);
TASK_PP(16'h11293,4);
TASK_PP(16'h11294,4);
TASK_PP(16'h11295,4);
TASK_PP(16'h11296,4);
TASK_PP(16'h11297,4);
TASK_PP(16'h11298,4);
TASK_PP(16'h11299,4);
TASK_PP(16'h1129A,4);
TASK_PP(16'h1129B,4);
TASK_PP(16'h1129C,4);
TASK_PP(16'h1129D,4);
TASK_PP(16'h1129E,4);
TASK_PP(16'h1129F,4);
TASK_PP(16'h112A0,4);
TASK_PP(16'h112A1,4);
TASK_PP(16'h112A2,4);
TASK_PP(16'h112A3,4);
TASK_PP(16'h112A4,4);
TASK_PP(16'h112A5,4);
TASK_PP(16'h112A6,4);
TASK_PP(16'h112A7,4);
TASK_PP(16'h112A8,4);
TASK_PP(16'h112A9,4);
TASK_PP(16'h112AA,4);
TASK_PP(16'h112AB,4);
TASK_PP(16'h112AC,4);
TASK_PP(16'h112AD,4);
TASK_PP(16'h112AE,4);
TASK_PP(16'h112AF,4);
TASK_PP(16'h112B0,4);
TASK_PP(16'h112B1,4);
TASK_PP(16'h112B2,4);
TASK_PP(16'h112B3,4);
TASK_PP(16'h112B4,4);
TASK_PP(16'h112B5,4);
TASK_PP(16'h112B6,4);
TASK_PP(16'h112B7,4);
TASK_PP(16'h112B8,4);
TASK_PP(16'h112B9,4);
TASK_PP(16'h112BA,4);
TASK_PP(16'h112BB,4);
TASK_PP(16'h112BC,4);
TASK_PP(16'h112BD,4);
TASK_PP(16'h112BE,4);
TASK_PP(16'h112BF,4);
TASK_PP(16'h112C0,4);
TASK_PP(16'h112C1,4);
TASK_PP(16'h112C2,4);
TASK_PP(16'h112C3,4);
TASK_PP(16'h112C4,4);
TASK_PP(16'h112C5,4);
TASK_PP(16'h112C6,4);
TASK_PP(16'h112C7,4);
TASK_PP(16'h112C8,4);
TASK_PP(16'h112C9,4);
TASK_PP(16'h112CA,4);
TASK_PP(16'h112CB,4);
TASK_PP(16'h112CC,4);
TASK_PP(16'h112CD,4);
TASK_PP(16'h112CE,4);
TASK_PP(16'h112CF,4);
TASK_PP(16'h112D0,4);
TASK_PP(16'h112D1,4);
TASK_PP(16'h112D2,4);
TASK_PP(16'h112D3,4);
TASK_PP(16'h112D4,4);
TASK_PP(16'h112D5,4);
TASK_PP(16'h112D6,4);
TASK_PP(16'h112D7,4);
TASK_PP(16'h112D8,4);
TASK_PP(16'h112D9,4);
TASK_PP(16'h112DA,4);
TASK_PP(16'h112DB,4);
TASK_PP(16'h112DC,4);
TASK_PP(16'h112DD,4);
TASK_PP(16'h112DE,4);
TASK_PP(16'h112DF,4);
TASK_PP(16'h112E0,4);
TASK_PP(16'h112E1,4);
TASK_PP(16'h112E2,4);
TASK_PP(16'h112E3,4);
TASK_PP(16'h112E4,4);
TASK_PP(16'h112E5,4);
TASK_PP(16'h112E6,4);
TASK_PP(16'h112E7,4);
TASK_PP(16'h112E8,4);
TASK_PP(16'h112E9,4);
TASK_PP(16'h112EA,4);
TASK_PP(16'h112EB,4);
TASK_PP(16'h112EC,4);
TASK_PP(16'h112ED,4);
TASK_PP(16'h112EE,4);
TASK_PP(16'h112EF,4);
TASK_PP(16'h112F0,4);
TASK_PP(16'h112F1,4);
TASK_PP(16'h112F2,4);
TASK_PP(16'h112F3,4);
TASK_PP(16'h112F4,4);
TASK_PP(16'h112F5,4);
TASK_PP(16'h112F6,4);
TASK_PP(16'h112F7,4);
TASK_PP(16'h112F8,4);
TASK_PP(16'h112F9,4);
TASK_PP(16'h112FA,4);
TASK_PP(16'h112FB,4);
TASK_PP(16'h112FC,4);
TASK_PP(16'h112FD,4);
TASK_PP(16'h112FE,4);
TASK_PP(16'h112FF,4);
TASK_PP(16'h11300,4);
TASK_PP(16'h11301,4);
TASK_PP(16'h11302,4);
TASK_PP(16'h11303,4);
TASK_PP(16'h11304,4);
TASK_PP(16'h11305,4);
TASK_PP(16'h11306,4);
TASK_PP(16'h11307,4);
TASK_PP(16'h11308,4);
TASK_PP(16'h11309,4);
TASK_PP(16'h1130A,4);
TASK_PP(16'h1130B,4);
TASK_PP(16'h1130C,4);
TASK_PP(16'h1130D,4);
TASK_PP(16'h1130E,4);
TASK_PP(16'h1130F,4);
TASK_PP(16'h11310,4);
TASK_PP(16'h11311,4);
TASK_PP(16'h11312,4);
TASK_PP(16'h11313,4);
TASK_PP(16'h11314,4);
TASK_PP(16'h11315,4);
TASK_PP(16'h11316,4);
TASK_PP(16'h11317,4);
TASK_PP(16'h11318,4);
TASK_PP(16'h11319,4);
TASK_PP(16'h1131A,4);
TASK_PP(16'h1131B,4);
TASK_PP(16'h1131C,4);
TASK_PP(16'h1131D,4);
TASK_PP(16'h1131E,4);
TASK_PP(16'h1131F,4);
TASK_PP(16'h11320,4);
TASK_PP(16'h11321,4);
TASK_PP(16'h11322,4);
TASK_PP(16'h11323,4);
TASK_PP(16'h11324,4);
TASK_PP(16'h11325,4);
TASK_PP(16'h11326,4);
TASK_PP(16'h11327,4);
TASK_PP(16'h11328,4);
TASK_PP(16'h11329,4);
TASK_PP(16'h1132A,4);
TASK_PP(16'h1132B,4);
TASK_PP(16'h1132C,4);
TASK_PP(16'h1132D,4);
TASK_PP(16'h1132E,4);
TASK_PP(16'h1132F,4);
TASK_PP(16'h11330,4);
TASK_PP(16'h11331,4);
TASK_PP(16'h11332,4);
TASK_PP(16'h11333,4);
TASK_PP(16'h11334,4);
TASK_PP(16'h11335,4);
TASK_PP(16'h11336,4);
TASK_PP(16'h11337,4);
TASK_PP(16'h11338,4);
TASK_PP(16'h11339,4);
TASK_PP(16'h1133A,4);
TASK_PP(16'h1133B,4);
TASK_PP(16'h1133C,4);
TASK_PP(16'h1133D,4);
TASK_PP(16'h1133E,4);
TASK_PP(16'h1133F,4);
TASK_PP(16'h11340,4);
TASK_PP(16'h11341,4);
TASK_PP(16'h11342,4);
TASK_PP(16'h11343,4);
TASK_PP(16'h11344,4);
TASK_PP(16'h11345,4);
TASK_PP(16'h11346,4);
TASK_PP(16'h11347,4);
TASK_PP(16'h11348,4);
TASK_PP(16'h11349,4);
TASK_PP(16'h1134A,4);
TASK_PP(16'h1134B,4);
TASK_PP(16'h1134C,4);
TASK_PP(16'h1134D,4);
TASK_PP(16'h1134E,4);
TASK_PP(16'h1134F,4);
TASK_PP(16'h11350,4);
TASK_PP(16'h11351,4);
TASK_PP(16'h11352,4);
TASK_PP(16'h11353,4);
TASK_PP(16'h11354,4);
TASK_PP(16'h11355,4);
TASK_PP(16'h11356,4);
TASK_PP(16'h11357,4);
TASK_PP(16'h11358,4);
TASK_PP(16'h11359,4);
TASK_PP(16'h1135A,4);
TASK_PP(16'h1135B,4);
TASK_PP(16'h1135C,4);
TASK_PP(16'h1135D,4);
TASK_PP(16'h1135E,4);
TASK_PP(16'h1135F,4);
TASK_PP(16'h11360,4);
TASK_PP(16'h11361,4);
TASK_PP(16'h11362,4);
TASK_PP(16'h11363,4);
TASK_PP(16'h11364,4);
TASK_PP(16'h11365,4);
TASK_PP(16'h11366,4);
TASK_PP(16'h11367,4);
TASK_PP(16'h11368,4);
TASK_PP(16'h11369,4);
TASK_PP(16'h1136A,4);
TASK_PP(16'h1136B,4);
TASK_PP(16'h1136C,4);
TASK_PP(16'h1136D,4);
TASK_PP(16'h1136E,4);
TASK_PP(16'h1136F,4);
TASK_PP(16'h11370,4);
TASK_PP(16'h11371,4);
TASK_PP(16'h11372,4);
TASK_PP(16'h11373,4);
TASK_PP(16'h11374,4);
TASK_PP(16'h11375,4);
TASK_PP(16'h11376,4);
TASK_PP(16'h11377,4);
TASK_PP(16'h11378,4);
TASK_PP(16'h11379,4);
TASK_PP(16'h1137A,4);
TASK_PP(16'h1137B,4);
TASK_PP(16'h1137C,4);
TASK_PP(16'h1137D,4);
TASK_PP(16'h1137E,4);
TASK_PP(16'h1137F,4);
TASK_PP(16'h11380,4);
TASK_PP(16'h11381,4);
TASK_PP(16'h11382,4);
TASK_PP(16'h11383,4);
TASK_PP(16'h11384,4);
TASK_PP(16'h11385,4);
TASK_PP(16'h11386,4);
TASK_PP(16'h11387,4);
TASK_PP(16'h11388,4);
TASK_PP(16'h11389,4);
TASK_PP(16'h1138A,4);
TASK_PP(16'h1138B,4);
TASK_PP(16'h1138C,4);
TASK_PP(16'h1138D,4);
TASK_PP(16'h1138E,4);
TASK_PP(16'h1138F,4);
TASK_PP(16'h11390,4);
TASK_PP(16'h11391,4);
TASK_PP(16'h11392,4);
TASK_PP(16'h11393,4);
TASK_PP(16'h11394,4);
TASK_PP(16'h11395,4);
TASK_PP(16'h11396,4);
TASK_PP(16'h11397,4);
TASK_PP(16'h11398,4);
TASK_PP(16'h11399,4);
TASK_PP(16'h1139A,4);
TASK_PP(16'h1139B,4);
TASK_PP(16'h1139C,4);
TASK_PP(16'h1139D,4);
TASK_PP(16'h1139E,4);
TASK_PP(16'h1139F,4);
TASK_PP(16'h113A0,4);
TASK_PP(16'h113A1,4);
TASK_PP(16'h113A2,4);
TASK_PP(16'h113A3,4);
TASK_PP(16'h113A4,4);
TASK_PP(16'h113A5,4);
TASK_PP(16'h113A6,4);
TASK_PP(16'h113A7,4);
TASK_PP(16'h113A8,4);
TASK_PP(16'h113A9,4);
TASK_PP(16'h113AA,4);
TASK_PP(16'h113AB,4);
TASK_PP(16'h113AC,4);
TASK_PP(16'h113AD,4);
TASK_PP(16'h113AE,4);
TASK_PP(16'h113AF,4);
TASK_PP(16'h113B0,4);
TASK_PP(16'h113B1,4);
TASK_PP(16'h113B2,4);
TASK_PP(16'h113B3,4);
TASK_PP(16'h113B4,4);
TASK_PP(16'h113B5,4);
TASK_PP(16'h113B6,4);
TASK_PP(16'h113B7,4);
TASK_PP(16'h113B8,4);
TASK_PP(16'h113B9,4);
TASK_PP(16'h113BA,4);
TASK_PP(16'h113BB,4);
TASK_PP(16'h113BC,4);
TASK_PP(16'h113BD,4);
TASK_PP(16'h113BE,4);
TASK_PP(16'h113BF,4);
TASK_PP(16'h113C0,4);
TASK_PP(16'h113C1,4);
TASK_PP(16'h113C2,4);
TASK_PP(16'h113C3,4);
TASK_PP(16'h113C4,4);
TASK_PP(16'h113C5,4);
TASK_PP(16'h113C6,4);
TASK_PP(16'h113C7,4);
TASK_PP(16'h113C8,4);
TASK_PP(16'h113C9,4);
TASK_PP(16'h113CA,4);
TASK_PP(16'h113CB,4);
TASK_PP(16'h113CC,4);
TASK_PP(16'h113CD,4);
TASK_PP(16'h113CE,4);
TASK_PP(16'h113CF,4);
TASK_PP(16'h113D0,4);
TASK_PP(16'h113D1,4);
TASK_PP(16'h113D2,4);
TASK_PP(16'h113D3,4);
TASK_PP(16'h113D4,4);
TASK_PP(16'h113D5,4);
TASK_PP(16'h113D6,4);
TASK_PP(16'h113D7,4);
TASK_PP(16'h113D8,4);
TASK_PP(16'h113D9,4);
TASK_PP(16'h113DA,4);
TASK_PP(16'h113DB,4);
TASK_PP(16'h113DC,4);
TASK_PP(16'h113DD,4);
TASK_PP(16'h113DE,4);
TASK_PP(16'h113DF,4);
TASK_PP(16'h113E0,4);
TASK_PP(16'h113E1,4);
TASK_PP(16'h113E2,4);
TASK_PP(16'h113E3,4);
TASK_PP(16'h113E4,4);
TASK_PP(16'h113E5,4);
TASK_PP(16'h113E6,4);
TASK_PP(16'h113E7,4);
TASK_PP(16'h113E8,4);
TASK_PP(16'h113E9,4);
TASK_PP(16'h113EA,4);
TASK_PP(16'h113EB,4);
TASK_PP(16'h113EC,4);
TASK_PP(16'h113ED,4);
TASK_PP(16'h113EE,4);
TASK_PP(16'h113EF,4);
TASK_PP(16'h113F0,4);
TASK_PP(16'h113F1,4);
TASK_PP(16'h113F2,4);
TASK_PP(16'h113F3,4);
TASK_PP(16'h113F4,4);
TASK_PP(16'h113F5,4);
TASK_PP(16'h113F6,4);
TASK_PP(16'h113F7,4);
TASK_PP(16'h113F8,4);
TASK_PP(16'h113F9,4);
TASK_PP(16'h113FA,4);
TASK_PP(16'h113FB,4);
TASK_PP(16'h113FC,4);
TASK_PP(16'h113FD,4);
TASK_PP(16'h113FE,4);
TASK_PP(16'h113FF,4);
TASK_PP(16'h11400,4);
TASK_PP(16'h11401,4);
TASK_PP(16'h11402,4);
TASK_PP(16'h11403,4);
TASK_PP(16'h11404,4);
TASK_PP(16'h11405,4);
TASK_PP(16'h11406,4);
TASK_PP(16'h11407,4);
TASK_PP(16'h11408,4);
TASK_PP(16'h11409,4);
TASK_PP(16'h1140A,4);
TASK_PP(16'h1140B,4);
TASK_PP(16'h1140C,4);
TASK_PP(16'h1140D,4);
TASK_PP(16'h1140E,4);
TASK_PP(16'h1140F,4);
TASK_PP(16'h11410,4);
TASK_PP(16'h11411,4);
TASK_PP(16'h11412,4);
TASK_PP(16'h11413,4);
TASK_PP(16'h11414,4);
TASK_PP(16'h11415,4);
TASK_PP(16'h11416,4);
TASK_PP(16'h11417,4);
TASK_PP(16'h11418,4);
TASK_PP(16'h11419,4);
TASK_PP(16'h1141A,4);
TASK_PP(16'h1141B,4);
TASK_PP(16'h1141C,4);
TASK_PP(16'h1141D,4);
TASK_PP(16'h1141E,4);
TASK_PP(16'h1141F,4);
TASK_PP(16'h11420,4);
TASK_PP(16'h11421,4);
TASK_PP(16'h11422,4);
TASK_PP(16'h11423,4);
TASK_PP(16'h11424,4);
TASK_PP(16'h11425,4);
TASK_PP(16'h11426,4);
TASK_PP(16'h11427,4);
TASK_PP(16'h11428,4);
TASK_PP(16'h11429,4);
TASK_PP(16'h1142A,4);
TASK_PP(16'h1142B,4);
TASK_PP(16'h1142C,4);
TASK_PP(16'h1142D,4);
TASK_PP(16'h1142E,4);
TASK_PP(16'h1142F,4);
TASK_PP(16'h11430,4);
TASK_PP(16'h11431,4);
TASK_PP(16'h11432,4);
TASK_PP(16'h11433,4);
TASK_PP(16'h11434,4);
TASK_PP(16'h11435,4);
TASK_PP(16'h11436,4);
TASK_PP(16'h11437,4);
TASK_PP(16'h11438,4);
TASK_PP(16'h11439,4);
TASK_PP(16'h1143A,4);
TASK_PP(16'h1143B,4);
TASK_PP(16'h1143C,4);
TASK_PP(16'h1143D,4);
TASK_PP(16'h1143E,4);
TASK_PP(16'h1143F,4);
TASK_PP(16'h11440,4);
TASK_PP(16'h11441,4);
TASK_PP(16'h11442,4);
TASK_PP(16'h11443,4);
TASK_PP(16'h11444,4);
TASK_PP(16'h11445,4);
TASK_PP(16'h11446,4);
TASK_PP(16'h11447,4);
TASK_PP(16'h11448,4);
TASK_PP(16'h11449,4);
TASK_PP(16'h1144A,4);
TASK_PP(16'h1144B,4);
TASK_PP(16'h1144C,4);
TASK_PP(16'h1144D,4);
TASK_PP(16'h1144E,4);
TASK_PP(16'h1144F,4);
TASK_PP(16'h11450,4);
TASK_PP(16'h11451,4);
TASK_PP(16'h11452,4);
TASK_PP(16'h11453,4);
TASK_PP(16'h11454,4);
TASK_PP(16'h11455,4);
TASK_PP(16'h11456,4);
TASK_PP(16'h11457,4);
TASK_PP(16'h11458,4);
TASK_PP(16'h11459,4);
TASK_PP(16'h1145A,4);
TASK_PP(16'h1145B,4);
TASK_PP(16'h1145C,4);
TASK_PP(16'h1145D,4);
TASK_PP(16'h1145E,4);
TASK_PP(16'h1145F,4);
TASK_PP(16'h11460,4);
TASK_PP(16'h11461,4);
TASK_PP(16'h11462,4);
TASK_PP(16'h11463,4);
TASK_PP(16'h11464,4);
TASK_PP(16'h11465,4);
TASK_PP(16'h11466,4);
TASK_PP(16'h11467,4);
TASK_PP(16'h11468,4);
TASK_PP(16'h11469,4);
TASK_PP(16'h1146A,4);
TASK_PP(16'h1146B,4);
TASK_PP(16'h1146C,4);
TASK_PP(16'h1146D,4);
TASK_PP(16'h1146E,4);
TASK_PP(16'h1146F,4);
TASK_PP(16'h11470,4);
TASK_PP(16'h11471,4);
TASK_PP(16'h11472,4);
TASK_PP(16'h11473,4);
TASK_PP(16'h11474,4);
TASK_PP(16'h11475,4);
TASK_PP(16'h11476,4);
TASK_PP(16'h11477,4);
TASK_PP(16'h11478,4);
TASK_PP(16'h11479,4);
TASK_PP(16'h1147A,4);
TASK_PP(16'h1147B,4);
TASK_PP(16'h1147C,4);
TASK_PP(16'h1147D,4);
TASK_PP(16'h1147E,4);
TASK_PP(16'h1147F,4);
TASK_PP(16'h11480,4);
TASK_PP(16'h11481,4);
TASK_PP(16'h11482,4);
TASK_PP(16'h11483,4);
TASK_PP(16'h11484,4);
TASK_PP(16'h11485,4);
TASK_PP(16'h11486,4);
TASK_PP(16'h11487,4);
TASK_PP(16'h11488,4);
TASK_PP(16'h11489,4);
TASK_PP(16'h1148A,4);
TASK_PP(16'h1148B,4);
TASK_PP(16'h1148C,4);
TASK_PP(16'h1148D,4);
TASK_PP(16'h1148E,4);
TASK_PP(16'h1148F,4);
TASK_PP(16'h11490,4);
TASK_PP(16'h11491,4);
TASK_PP(16'h11492,4);
TASK_PP(16'h11493,4);
TASK_PP(16'h11494,4);
TASK_PP(16'h11495,4);
TASK_PP(16'h11496,4);
TASK_PP(16'h11497,4);
TASK_PP(16'h11498,4);
TASK_PP(16'h11499,4);
TASK_PP(16'h1149A,4);
TASK_PP(16'h1149B,4);
TASK_PP(16'h1149C,4);
TASK_PP(16'h1149D,4);
TASK_PP(16'h1149E,4);
TASK_PP(16'h1149F,4);
TASK_PP(16'h114A0,4);
TASK_PP(16'h114A1,4);
TASK_PP(16'h114A2,4);
TASK_PP(16'h114A3,4);
TASK_PP(16'h114A4,4);
TASK_PP(16'h114A5,4);
TASK_PP(16'h114A6,4);
TASK_PP(16'h114A7,4);
TASK_PP(16'h114A8,4);
TASK_PP(16'h114A9,4);
TASK_PP(16'h114AA,4);
TASK_PP(16'h114AB,4);
TASK_PP(16'h114AC,4);
TASK_PP(16'h114AD,4);
TASK_PP(16'h114AE,4);
TASK_PP(16'h114AF,4);
TASK_PP(16'h114B0,4);
TASK_PP(16'h114B1,4);
TASK_PP(16'h114B2,4);
TASK_PP(16'h114B3,4);
TASK_PP(16'h114B4,4);
TASK_PP(16'h114B5,4);
TASK_PP(16'h114B6,4);
TASK_PP(16'h114B7,4);
TASK_PP(16'h114B8,4);
TASK_PP(16'h114B9,4);
TASK_PP(16'h114BA,4);
TASK_PP(16'h114BB,4);
TASK_PP(16'h114BC,4);
TASK_PP(16'h114BD,4);
TASK_PP(16'h114BE,4);
TASK_PP(16'h114BF,4);
TASK_PP(16'h114C0,4);
TASK_PP(16'h114C1,4);
TASK_PP(16'h114C2,4);
TASK_PP(16'h114C3,4);
TASK_PP(16'h114C4,4);
TASK_PP(16'h114C5,4);
TASK_PP(16'h114C6,4);
TASK_PP(16'h114C7,4);
TASK_PP(16'h114C8,4);
TASK_PP(16'h114C9,4);
TASK_PP(16'h114CA,4);
TASK_PP(16'h114CB,4);
TASK_PP(16'h114CC,4);
TASK_PP(16'h114CD,4);
TASK_PP(16'h114CE,4);
TASK_PP(16'h114CF,4);
TASK_PP(16'h114D0,4);
TASK_PP(16'h114D1,4);
TASK_PP(16'h114D2,4);
TASK_PP(16'h114D3,4);
TASK_PP(16'h114D4,4);
TASK_PP(16'h114D5,4);
TASK_PP(16'h114D6,4);
TASK_PP(16'h114D7,4);
TASK_PP(16'h114D8,4);
TASK_PP(16'h114D9,4);
TASK_PP(16'h114DA,4);
TASK_PP(16'h114DB,4);
TASK_PP(16'h114DC,4);
TASK_PP(16'h114DD,4);
TASK_PP(16'h114DE,4);
TASK_PP(16'h114DF,4);
TASK_PP(16'h114E0,4);
TASK_PP(16'h114E1,4);
TASK_PP(16'h114E2,4);
TASK_PP(16'h114E3,4);
TASK_PP(16'h114E4,4);
TASK_PP(16'h114E5,4);
TASK_PP(16'h114E6,4);
TASK_PP(16'h114E7,4);
TASK_PP(16'h114E8,4);
TASK_PP(16'h114E9,4);
TASK_PP(16'h114EA,4);
TASK_PP(16'h114EB,4);
TASK_PP(16'h114EC,4);
TASK_PP(16'h114ED,4);
TASK_PP(16'h114EE,4);
TASK_PP(16'h114EF,4);
TASK_PP(16'h114F0,4);
TASK_PP(16'h114F1,4);
TASK_PP(16'h114F2,4);
TASK_PP(16'h114F3,4);
TASK_PP(16'h114F4,4);
TASK_PP(16'h114F5,4);
TASK_PP(16'h114F6,4);
TASK_PP(16'h114F7,4);
TASK_PP(16'h114F8,4);
TASK_PP(16'h114F9,4);
TASK_PP(16'h114FA,4);
TASK_PP(16'h114FB,4);
TASK_PP(16'h114FC,4);
TASK_PP(16'h114FD,4);
TASK_PP(16'h114FE,4);
TASK_PP(16'h114FF,4);
TASK_PP(16'h11500,4);
TASK_PP(16'h11501,4);
TASK_PP(16'h11502,4);
TASK_PP(16'h11503,4);
TASK_PP(16'h11504,4);
TASK_PP(16'h11505,4);
TASK_PP(16'h11506,4);
TASK_PP(16'h11507,4);
TASK_PP(16'h11508,4);
TASK_PP(16'h11509,4);
TASK_PP(16'h1150A,4);
TASK_PP(16'h1150B,4);
TASK_PP(16'h1150C,4);
TASK_PP(16'h1150D,4);
TASK_PP(16'h1150E,4);
TASK_PP(16'h1150F,4);
TASK_PP(16'h11510,4);
TASK_PP(16'h11511,4);
TASK_PP(16'h11512,4);
TASK_PP(16'h11513,4);
TASK_PP(16'h11514,4);
TASK_PP(16'h11515,4);
TASK_PP(16'h11516,4);
TASK_PP(16'h11517,4);
TASK_PP(16'h11518,4);
TASK_PP(16'h11519,4);
TASK_PP(16'h1151A,4);
TASK_PP(16'h1151B,4);
TASK_PP(16'h1151C,4);
TASK_PP(16'h1151D,4);
TASK_PP(16'h1151E,4);
TASK_PP(16'h1151F,4);
TASK_PP(16'h11520,4);
TASK_PP(16'h11521,4);
TASK_PP(16'h11522,4);
TASK_PP(16'h11523,4);
TASK_PP(16'h11524,4);
TASK_PP(16'h11525,4);
TASK_PP(16'h11526,4);
TASK_PP(16'h11527,4);
TASK_PP(16'h11528,4);
TASK_PP(16'h11529,4);
TASK_PP(16'h1152A,4);
TASK_PP(16'h1152B,4);
TASK_PP(16'h1152C,4);
TASK_PP(16'h1152D,4);
TASK_PP(16'h1152E,4);
TASK_PP(16'h1152F,4);
TASK_PP(16'h11530,4);
TASK_PP(16'h11531,4);
TASK_PP(16'h11532,4);
TASK_PP(16'h11533,4);
TASK_PP(16'h11534,4);
TASK_PP(16'h11535,4);
TASK_PP(16'h11536,4);
TASK_PP(16'h11537,4);
TASK_PP(16'h11538,4);
TASK_PP(16'h11539,4);
TASK_PP(16'h1153A,4);
TASK_PP(16'h1153B,4);
TASK_PP(16'h1153C,4);
TASK_PP(16'h1153D,4);
TASK_PP(16'h1153E,4);
TASK_PP(16'h1153F,4);
TASK_PP(16'h11540,4);
TASK_PP(16'h11541,4);
TASK_PP(16'h11542,4);
TASK_PP(16'h11543,4);
TASK_PP(16'h11544,4);
TASK_PP(16'h11545,4);
TASK_PP(16'h11546,4);
TASK_PP(16'h11547,4);
TASK_PP(16'h11548,4);
TASK_PP(16'h11549,4);
TASK_PP(16'h1154A,4);
TASK_PP(16'h1154B,4);
TASK_PP(16'h1154C,4);
TASK_PP(16'h1154D,4);
TASK_PP(16'h1154E,4);
TASK_PP(16'h1154F,4);
TASK_PP(16'h11550,4);
TASK_PP(16'h11551,4);
TASK_PP(16'h11552,4);
TASK_PP(16'h11553,4);
TASK_PP(16'h11554,4);
TASK_PP(16'h11555,4);
TASK_PP(16'h11556,4);
TASK_PP(16'h11557,4);
TASK_PP(16'h11558,4);
TASK_PP(16'h11559,4);
TASK_PP(16'h1155A,4);
TASK_PP(16'h1155B,4);
TASK_PP(16'h1155C,4);
TASK_PP(16'h1155D,4);
TASK_PP(16'h1155E,4);
TASK_PP(16'h1155F,4);
TASK_PP(16'h11560,4);
TASK_PP(16'h11561,4);
TASK_PP(16'h11562,4);
TASK_PP(16'h11563,4);
TASK_PP(16'h11564,4);
TASK_PP(16'h11565,4);
TASK_PP(16'h11566,4);
TASK_PP(16'h11567,4);
TASK_PP(16'h11568,4);
TASK_PP(16'h11569,4);
TASK_PP(16'h1156A,4);
TASK_PP(16'h1156B,4);
TASK_PP(16'h1156C,4);
TASK_PP(16'h1156D,4);
TASK_PP(16'h1156E,4);
TASK_PP(16'h1156F,4);
TASK_PP(16'h11570,4);
TASK_PP(16'h11571,4);
TASK_PP(16'h11572,4);
TASK_PP(16'h11573,4);
TASK_PP(16'h11574,4);
TASK_PP(16'h11575,4);
TASK_PP(16'h11576,4);
TASK_PP(16'h11577,4);
TASK_PP(16'h11578,4);
TASK_PP(16'h11579,4);
TASK_PP(16'h1157A,4);
TASK_PP(16'h1157B,4);
TASK_PP(16'h1157C,4);
TASK_PP(16'h1157D,4);
TASK_PP(16'h1157E,4);
TASK_PP(16'h1157F,4);
TASK_PP(16'h11580,4);
TASK_PP(16'h11581,4);
TASK_PP(16'h11582,4);
TASK_PP(16'h11583,4);
TASK_PP(16'h11584,4);
TASK_PP(16'h11585,4);
TASK_PP(16'h11586,4);
TASK_PP(16'h11587,4);
TASK_PP(16'h11588,4);
TASK_PP(16'h11589,4);
TASK_PP(16'h1158A,4);
TASK_PP(16'h1158B,4);
TASK_PP(16'h1158C,4);
TASK_PP(16'h1158D,4);
TASK_PP(16'h1158E,4);
TASK_PP(16'h1158F,4);
TASK_PP(16'h11590,4);
TASK_PP(16'h11591,4);
TASK_PP(16'h11592,4);
TASK_PP(16'h11593,4);
TASK_PP(16'h11594,4);
TASK_PP(16'h11595,4);
TASK_PP(16'h11596,4);
TASK_PP(16'h11597,4);
TASK_PP(16'h11598,4);
TASK_PP(16'h11599,4);
TASK_PP(16'h1159A,4);
TASK_PP(16'h1159B,4);
TASK_PP(16'h1159C,4);
TASK_PP(16'h1159D,4);
TASK_PP(16'h1159E,4);
TASK_PP(16'h1159F,4);
TASK_PP(16'h115A0,4);
TASK_PP(16'h115A1,4);
TASK_PP(16'h115A2,4);
TASK_PP(16'h115A3,4);
TASK_PP(16'h115A4,4);
TASK_PP(16'h115A5,4);
TASK_PP(16'h115A6,4);
TASK_PP(16'h115A7,4);
TASK_PP(16'h115A8,4);
TASK_PP(16'h115A9,4);
TASK_PP(16'h115AA,4);
TASK_PP(16'h115AB,4);
TASK_PP(16'h115AC,4);
TASK_PP(16'h115AD,4);
TASK_PP(16'h115AE,4);
TASK_PP(16'h115AF,4);
TASK_PP(16'h115B0,4);
TASK_PP(16'h115B1,4);
TASK_PP(16'h115B2,4);
TASK_PP(16'h115B3,4);
TASK_PP(16'h115B4,4);
TASK_PP(16'h115B5,4);
TASK_PP(16'h115B6,4);
TASK_PP(16'h115B7,4);
TASK_PP(16'h115B8,4);
TASK_PP(16'h115B9,4);
TASK_PP(16'h115BA,4);
TASK_PP(16'h115BB,4);
TASK_PP(16'h115BC,4);
TASK_PP(16'h115BD,4);
TASK_PP(16'h115BE,4);
TASK_PP(16'h115BF,4);
TASK_PP(16'h115C0,4);
TASK_PP(16'h115C1,4);
TASK_PP(16'h115C2,4);
TASK_PP(16'h115C3,4);
TASK_PP(16'h115C4,4);
TASK_PP(16'h115C5,4);
TASK_PP(16'h115C6,4);
TASK_PP(16'h115C7,4);
TASK_PP(16'h115C8,4);
TASK_PP(16'h115C9,4);
TASK_PP(16'h115CA,4);
TASK_PP(16'h115CB,4);
TASK_PP(16'h115CC,4);
TASK_PP(16'h115CD,4);
TASK_PP(16'h115CE,4);
TASK_PP(16'h115CF,4);
TASK_PP(16'h115D0,4);
TASK_PP(16'h115D1,4);
TASK_PP(16'h115D2,4);
TASK_PP(16'h115D3,4);
TASK_PP(16'h115D4,4);
TASK_PP(16'h115D5,4);
TASK_PP(16'h115D6,4);
TASK_PP(16'h115D7,4);
TASK_PP(16'h115D8,4);
TASK_PP(16'h115D9,4);
TASK_PP(16'h115DA,4);
TASK_PP(16'h115DB,4);
TASK_PP(16'h115DC,4);
TASK_PP(16'h115DD,4);
TASK_PP(16'h115DE,4);
TASK_PP(16'h115DF,4);
TASK_PP(16'h115E0,4);
TASK_PP(16'h115E1,4);
TASK_PP(16'h115E2,4);
TASK_PP(16'h115E3,4);
TASK_PP(16'h115E4,4);
TASK_PP(16'h115E5,4);
TASK_PP(16'h115E6,4);
TASK_PP(16'h115E7,4);
TASK_PP(16'h115E8,4);
TASK_PP(16'h115E9,4);
TASK_PP(16'h115EA,4);
TASK_PP(16'h115EB,4);
TASK_PP(16'h115EC,4);
TASK_PP(16'h115ED,4);
TASK_PP(16'h115EE,4);
TASK_PP(16'h115EF,4);
TASK_PP(16'h115F0,4);
TASK_PP(16'h115F1,4);
TASK_PP(16'h115F2,4);
TASK_PP(16'h115F3,4);
TASK_PP(16'h115F4,4);
TASK_PP(16'h115F5,4);
TASK_PP(16'h115F6,4);
TASK_PP(16'h115F7,4);
TASK_PP(16'h115F8,4);
TASK_PP(16'h115F9,4);
TASK_PP(16'h115FA,4);
TASK_PP(16'h115FB,4);
TASK_PP(16'h115FC,4);
TASK_PP(16'h115FD,4);
TASK_PP(16'h115FE,4);
TASK_PP(16'h115FF,4);
TASK_PP(16'h11600,4);
TASK_PP(16'h11601,4);
TASK_PP(16'h11602,4);
TASK_PP(16'h11603,4);
TASK_PP(16'h11604,4);
TASK_PP(16'h11605,4);
TASK_PP(16'h11606,4);
TASK_PP(16'h11607,4);
TASK_PP(16'h11608,4);
TASK_PP(16'h11609,4);
TASK_PP(16'h1160A,4);
TASK_PP(16'h1160B,4);
TASK_PP(16'h1160C,4);
TASK_PP(16'h1160D,4);
TASK_PP(16'h1160E,4);
TASK_PP(16'h1160F,4);
TASK_PP(16'h11610,4);
TASK_PP(16'h11611,4);
TASK_PP(16'h11612,4);
TASK_PP(16'h11613,4);
TASK_PP(16'h11614,4);
TASK_PP(16'h11615,4);
TASK_PP(16'h11616,4);
TASK_PP(16'h11617,4);
TASK_PP(16'h11618,4);
TASK_PP(16'h11619,4);
TASK_PP(16'h1161A,4);
TASK_PP(16'h1161B,4);
TASK_PP(16'h1161C,4);
TASK_PP(16'h1161D,4);
TASK_PP(16'h1161E,4);
TASK_PP(16'h1161F,4);
TASK_PP(16'h11620,4);
TASK_PP(16'h11621,4);
TASK_PP(16'h11622,4);
TASK_PP(16'h11623,4);
TASK_PP(16'h11624,4);
TASK_PP(16'h11625,4);
TASK_PP(16'h11626,4);
TASK_PP(16'h11627,4);
TASK_PP(16'h11628,4);
TASK_PP(16'h11629,4);
TASK_PP(16'h1162A,4);
TASK_PP(16'h1162B,4);
TASK_PP(16'h1162C,4);
TASK_PP(16'h1162D,4);
TASK_PP(16'h1162E,4);
TASK_PP(16'h1162F,4);
TASK_PP(16'h11630,4);
TASK_PP(16'h11631,4);
TASK_PP(16'h11632,4);
TASK_PP(16'h11633,4);
TASK_PP(16'h11634,4);
TASK_PP(16'h11635,4);
TASK_PP(16'h11636,4);
TASK_PP(16'h11637,4);
TASK_PP(16'h11638,4);
TASK_PP(16'h11639,4);
TASK_PP(16'h1163A,4);
TASK_PP(16'h1163B,4);
TASK_PP(16'h1163C,4);
TASK_PP(16'h1163D,4);
TASK_PP(16'h1163E,4);
TASK_PP(16'h1163F,4);
TASK_PP(16'h11640,4);
TASK_PP(16'h11641,4);
TASK_PP(16'h11642,4);
TASK_PP(16'h11643,4);
TASK_PP(16'h11644,4);
TASK_PP(16'h11645,4);
TASK_PP(16'h11646,4);
TASK_PP(16'h11647,4);
TASK_PP(16'h11648,4);
TASK_PP(16'h11649,4);
TASK_PP(16'h1164A,4);
TASK_PP(16'h1164B,4);
TASK_PP(16'h1164C,4);
TASK_PP(16'h1164D,4);
TASK_PP(16'h1164E,4);
TASK_PP(16'h1164F,4);
TASK_PP(16'h11650,4);
TASK_PP(16'h11651,4);
TASK_PP(16'h11652,4);
TASK_PP(16'h11653,4);
TASK_PP(16'h11654,4);
TASK_PP(16'h11655,4);
TASK_PP(16'h11656,4);
TASK_PP(16'h11657,4);
TASK_PP(16'h11658,4);
TASK_PP(16'h11659,4);
TASK_PP(16'h1165A,4);
TASK_PP(16'h1165B,4);
TASK_PP(16'h1165C,4);
TASK_PP(16'h1165D,4);
TASK_PP(16'h1165E,4);
TASK_PP(16'h1165F,4);
TASK_PP(16'h11660,4);
TASK_PP(16'h11661,4);
TASK_PP(16'h11662,4);
TASK_PP(16'h11663,4);
TASK_PP(16'h11664,4);
TASK_PP(16'h11665,4);
TASK_PP(16'h11666,4);
TASK_PP(16'h11667,4);
TASK_PP(16'h11668,4);
TASK_PP(16'h11669,4);
TASK_PP(16'h1166A,4);
TASK_PP(16'h1166B,4);
TASK_PP(16'h1166C,4);
TASK_PP(16'h1166D,4);
TASK_PP(16'h1166E,4);
TASK_PP(16'h1166F,4);
TASK_PP(16'h11670,4);
TASK_PP(16'h11671,4);
TASK_PP(16'h11672,4);
TASK_PP(16'h11673,4);
TASK_PP(16'h11674,4);
TASK_PP(16'h11675,4);
TASK_PP(16'h11676,4);
TASK_PP(16'h11677,4);
TASK_PP(16'h11678,4);
TASK_PP(16'h11679,4);
TASK_PP(16'h1167A,4);
TASK_PP(16'h1167B,4);
TASK_PP(16'h1167C,4);
TASK_PP(16'h1167D,4);
TASK_PP(16'h1167E,4);
TASK_PP(16'h1167F,4);
TASK_PP(16'h11680,4);
TASK_PP(16'h11681,4);
TASK_PP(16'h11682,4);
TASK_PP(16'h11683,4);
TASK_PP(16'h11684,4);
TASK_PP(16'h11685,4);
TASK_PP(16'h11686,4);
TASK_PP(16'h11687,4);
TASK_PP(16'h11688,4);
TASK_PP(16'h11689,4);
TASK_PP(16'h1168A,4);
TASK_PP(16'h1168B,4);
TASK_PP(16'h1168C,4);
TASK_PP(16'h1168D,4);
TASK_PP(16'h1168E,4);
TASK_PP(16'h1168F,4);
TASK_PP(16'h11690,4);
TASK_PP(16'h11691,4);
TASK_PP(16'h11692,4);
TASK_PP(16'h11693,4);
TASK_PP(16'h11694,4);
TASK_PP(16'h11695,4);
TASK_PP(16'h11696,4);
TASK_PP(16'h11697,4);
TASK_PP(16'h11698,4);
TASK_PP(16'h11699,4);
TASK_PP(16'h1169A,4);
TASK_PP(16'h1169B,4);
TASK_PP(16'h1169C,4);
TASK_PP(16'h1169D,4);
TASK_PP(16'h1169E,4);
TASK_PP(16'h1169F,4);
TASK_PP(16'h116A0,4);
TASK_PP(16'h116A1,4);
TASK_PP(16'h116A2,4);
TASK_PP(16'h116A3,4);
TASK_PP(16'h116A4,4);
TASK_PP(16'h116A5,4);
TASK_PP(16'h116A6,4);
TASK_PP(16'h116A7,4);
TASK_PP(16'h116A8,4);
TASK_PP(16'h116A9,4);
TASK_PP(16'h116AA,4);
TASK_PP(16'h116AB,4);
TASK_PP(16'h116AC,4);
TASK_PP(16'h116AD,4);
TASK_PP(16'h116AE,4);
TASK_PP(16'h116AF,4);
TASK_PP(16'h116B0,4);
TASK_PP(16'h116B1,4);
TASK_PP(16'h116B2,4);
TASK_PP(16'h116B3,4);
TASK_PP(16'h116B4,4);
TASK_PP(16'h116B5,4);
TASK_PP(16'h116B6,4);
TASK_PP(16'h116B7,4);
TASK_PP(16'h116B8,4);
TASK_PP(16'h116B9,4);
TASK_PP(16'h116BA,4);
TASK_PP(16'h116BB,4);
TASK_PP(16'h116BC,4);
TASK_PP(16'h116BD,4);
TASK_PP(16'h116BE,4);
TASK_PP(16'h116BF,4);
TASK_PP(16'h116C0,4);
TASK_PP(16'h116C1,4);
TASK_PP(16'h116C2,4);
TASK_PP(16'h116C3,4);
TASK_PP(16'h116C4,4);
TASK_PP(16'h116C5,4);
TASK_PP(16'h116C6,4);
TASK_PP(16'h116C7,4);
TASK_PP(16'h116C8,4);
TASK_PP(16'h116C9,4);
TASK_PP(16'h116CA,4);
TASK_PP(16'h116CB,4);
TASK_PP(16'h116CC,4);
TASK_PP(16'h116CD,4);
TASK_PP(16'h116CE,4);
TASK_PP(16'h116CF,4);
TASK_PP(16'h116D0,4);
TASK_PP(16'h116D1,4);
TASK_PP(16'h116D2,4);
TASK_PP(16'h116D3,4);
TASK_PP(16'h116D4,4);
TASK_PP(16'h116D5,4);
TASK_PP(16'h116D6,4);
TASK_PP(16'h116D7,4);
TASK_PP(16'h116D8,4);
TASK_PP(16'h116D9,4);
TASK_PP(16'h116DA,4);
TASK_PP(16'h116DB,4);
TASK_PP(16'h116DC,4);
TASK_PP(16'h116DD,4);
TASK_PP(16'h116DE,4);
TASK_PP(16'h116DF,4);
TASK_PP(16'h116E0,4);
TASK_PP(16'h116E1,4);
TASK_PP(16'h116E2,4);
TASK_PP(16'h116E3,4);
TASK_PP(16'h116E4,4);
TASK_PP(16'h116E5,4);
TASK_PP(16'h116E6,4);
TASK_PP(16'h116E7,4);
TASK_PP(16'h116E8,4);
TASK_PP(16'h116E9,4);
TASK_PP(16'h116EA,4);
TASK_PP(16'h116EB,4);
TASK_PP(16'h116EC,4);
TASK_PP(16'h116ED,4);
TASK_PP(16'h116EE,4);
TASK_PP(16'h116EF,4);
TASK_PP(16'h116F0,4);
TASK_PP(16'h116F1,4);
TASK_PP(16'h116F2,4);
TASK_PP(16'h116F3,4);
TASK_PP(16'h116F4,4);
TASK_PP(16'h116F5,4);
TASK_PP(16'h116F6,4);
TASK_PP(16'h116F7,4);
TASK_PP(16'h116F8,4);
TASK_PP(16'h116F9,4);
TASK_PP(16'h116FA,4);
TASK_PP(16'h116FB,4);
TASK_PP(16'h116FC,4);
TASK_PP(16'h116FD,4);
TASK_PP(16'h116FE,4);
TASK_PP(16'h116FF,4);
TASK_PP(16'h11700,4);
TASK_PP(16'h11701,4);
TASK_PP(16'h11702,4);
TASK_PP(16'h11703,4);
TASK_PP(16'h11704,4);
TASK_PP(16'h11705,4);
TASK_PP(16'h11706,4);
TASK_PP(16'h11707,4);
TASK_PP(16'h11708,4);
TASK_PP(16'h11709,4);
TASK_PP(16'h1170A,4);
TASK_PP(16'h1170B,4);
TASK_PP(16'h1170C,4);
TASK_PP(16'h1170D,4);
TASK_PP(16'h1170E,4);
TASK_PP(16'h1170F,4);
TASK_PP(16'h11710,4);
TASK_PP(16'h11711,4);
TASK_PP(16'h11712,4);
TASK_PP(16'h11713,4);
TASK_PP(16'h11714,4);
TASK_PP(16'h11715,4);
TASK_PP(16'h11716,4);
TASK_PP(16'h11717,4);
TASK_PP(16'h11718,4);
TASK_PP(16'h11719,4);
TASK_PP(16'h1171A,4);
TASK_PP(16'h1171B,4);
TASK_PP(16'h1171C,4);
TASK_PP(16'h1171D,4);
TASK_PP(16'h1171E,4);
TASK_PP(16'h1171F,4);
TASK_PP(16'h11720,4);
TASK_PP(16'h11721,4);
TASK_PP(16'h11722,4);
TASK_PP(16'h11723,4);
TASK_PP(16'h11724,4);
TASK_PP(16'h11725,4);
TASK_PP(16'h11726,4);
TASK_PP(16'h11727,4);
TASK_PP(16'h11728,4);
TASK_PP(16'h11729,4);
TASK_PP(16'h1172A,4);
TASK_PP(16'h1172B,4);
TASK_PP(16'h1172C,4);
TASK_PP(16'h1172D,4);
TASK_PP(16'h1172E,4);
TASK_PP(16'h1172F,4);
TASK_PP(16'h11730,4);
TASK_PP(16'h11731,4);
TASK_PP(16'h11732,4);
TASK_PP(16'h11733,4);
TASK_PP(16'h11734,4);
TASK_PP(16'h11735,4);
TASK_PP(16'h11736,4);
TASK_PP(16'h11737,4);
TASK_PP(16'h11738,4);
TASK_PP(16'h11739,4);
TASK_PP(16'h1173A,4);
TASK_PP(16'h1173B,4);
TASK_PP(16'h1173C,4);
TASK_PP(16'h1173D,4);
TASK_PP(16'h1173E,4);
TASK_PP(16'h1173F,4);
TASK_PP(16'h11740,4);
TASK_PP(16'h11741,4);
TASK_PP(16'h11742,4);
TASK_PP(16'h11743,4);
TASK_PP(16'h11744,4);
TASK_PP(16'h11745,4);
TASK_PP(16'h11746,4);
TASK_PP(16'h11747,4);
TASK_PP(16'h11748,4);
TASK_PP(16'h11749,4);
TASK_PP(16'h1174A,4);
TASK_PP(16'h1174B,4);
TASK_PP(16'h1174C,4);
TASK_PP(16'h1174D,4);
TASK_PP(16'h1174E,4);
TASK_PP(16'h1174F,4);
TASK_PP(16'h11750,4);
TASK_PP(16'h11751,4);
TASK_PP(16'h11752,4);
TASK_PP(16'h11753,4);
TASK_PP(16'h11754,4);
TASK_PP(16'h11755,4);
TASK_PP(16'h11756,4);
TASK_PP(16'h11757,4);
TASK_PP(16'h11758,4);
TASK_PP(16'h11759,4);
TASK_PP(16'h1175A,4);
TASK_PP(16'h1175B,4);
TASK_PP(16'h1175C,4);
TASK_PP(16'h1175D,4);
TASK_PP(16'h1175E,4);
TASK_PP(16'h1175F,4);
TASK_PP(16'h11760,4);
TASK_PP(16'h11761,4);
TASK_PP(16'h11762,4);
TASK_PP(16'h11763,4);
TASK_PP(16'h11764,4);
TASK_PP(16'h11765,4);
TASK_PP(16'h11766,4);
TASK_PP(16'h11767,4);
TASK_PP(16'h11768,4);
TASK_PP(16'h11769,4);
TASK_PP(16'h1176A,4);
TASK_PP(16'h1176B,4);
TASK_PP(16'h1176C,4);
TASK_PP(16'h1176D,4);
TASK_PP(16'h1176E,4);
TASK_PP(16'h1176F,4);
TASK_PP(16'h11770,4);
TASK_PP(16'h11771,4);
TASK_PP(16'h11772,4);
TASK_PP(16'h11773,4);
TASK_PP(16'h11774,4);
TASK_PP(16'h11775,4);
TASK_PP(16'h11776,4);
TASK_PP(16'h11777,4);
TASK_PP(16'h11778,4);
TASK_PP(16'h11779,4);
TASK_PP(16'h1177A,4);
TASK_PP(16'h1177B,4);
TASK_PP(16'h1177C,4);
TASK_PP(16'h1177D,4);
TASK_PP(16'h1177E,4);
TASK_PP(16'h1177F,4);
TASK_PP(16'h11780,4);
TASK_PP(16'h11781,4);
TASK_PP(16'h11782,4);
TASK_PP(16'h11783,4);
TASK_PP(16'h11784,4);
TASK_PP(16'h11785,4);
TASK_PP(16'h11786,4);
TASK_PP(16'h11787,4);
TASK_PP(16'h11788,4);
TASK_PP(16'h11789,4);
TASK_PP(16'h1178A,4);
TASK_PP(16'h1178B,4);
TASK_PP(16'h1178C,4);
TASK_PP(16'h1178D,4);
TASK_PP(16'h1178E,4);
TASK_PP(16'h1178F,4);
TASK_PP(16'h11790,4);
TASK_PP(16'h11791,4);
TASK_PP(16'h11792,4);
TASK_PP(16'h11793,4);
TASK_PP(16'h11794,4);
TASK_PP(16'h11795,4);
TASK_PP(16'h11796,4);
TASK_PP(16'h11797,4);
TASK_PP(16'h11798,4);
TASK_PP(16'h11799,4);
TASK_PP(16'h1179A,4);
TASK_PP(16'h1179B,4);
TASK_PP(16'h1179C,4);
TASK_PP(16'h1179D,4);
TASK_PP(16'h1179E,4);
TASK_PP(16'h1179F,4);
TASK_PP(16'h117A0,4);
TASK_PP(16'h117A1,4);
TASK_PP(16'h117A2,4);
TASK_PP(16'h117A3,4);
TASK_PP(16'h117A4,4);
TASK_PP(16'h117A5,4);
TASK_PP(16'h117A6,4);
TASK_PP(16'h117A7,4);
TASK_PP(16'h117A8,4);
TASK_PP(16'h117A9,4);
TASK_PP(16'h117AA,4);
TASK_PP(16'h117AB,4);
TASK_PP(16'h117AC,4);
TASK_PP(16'h117AD,4);
TASK_PP(16'h117AE,4);
TASK_PP(16'h117AF,4);
TASK_PP(16'h117B0,4);
TASK_PP(16'h117B1,4);
TASK_PP(16'h117B2,4);
TASK_PP(16'h117B3,4);
TASK_PP(16'h117B4,4);
TASK_PP(16'h117B5,4);
TASK_PP(16'h117B6,4);
TASK_PP(16'h117B7,4);
TASK_PP(16'h117B8,4);
TASK_PP(16'h117B9,4);
TASK_PP(16'h117BA,4);
TASK_PP(16'h117BB,4);
TASK_PP(16'h117BC,4);
TASK_PP(16'h117BD,4);
TASK_PP(16'h117BE,4);
TASK_PP(16'h117BF,4);
TASK_PP(16'h117C0,4);
TASK_PP(16'h117C1,4);
TASK_PP(16'h117C2,4);
TASK_PP(16'h117C3,4);
TASK_PP(16'h117C4,4);
TASK_PP(16'h117C5,4);
TASK_PP(16'h117C6,4);
TASK_PP(16'h117C7,4);
TASK_PP(16'h117C8,4);
TASK_PP(16'h117C9,4);
TASK_PP(16'h117CA,4);
TASK_PP(16'h117CB,4);
TASK_PP(16'h117CC,4);
TASK_PP(16'h117CD,4);
TASK_PP(16'h117CE,4);
TASK_PP(16'h117CF,4);
TASK_PP(16'h117D0,4);
TASK_PP(16'h117D1,4);
TASK_PP(16'h117D2,4);
TASK_PP(16'h117D3,4);
TASK_PP(16'h117D4,4);
TASK_PP(16'h117D5,4);
TASK_PP(16'h117D6,4);
TASK_PP(16'h117D7,4);
TASK_PP(16'h117D8,4);
TASK_PP(16'h117D9,4);
TASK_PP(16'h117DA,4);
TASK_PP(16'h117DB,4);
TASK_PP(16'h117DC,4);
TASK_PP(16'h117DD,4);
TASK_PP(16'h117DE,4);
TASK_PP(16'h117DF,4);
TASK_PP(16'h117E0,4);
TASK_PP(16'h117E1,4);
TASK_PP(16'h117E2,4);
TASK_PP(16'h117E3,4);
TASK_PP(16'h117E4,4);
TASK_PP(16'h117E5,4);
TASK_PP(16'h117E6,4);
TASK_PP(16'h117E7,4);
TASK_PP(16'h117E8,4);
TASK_PP(16'h117E9,4);
TASK_PP(16'h117EA,4);
TASK_PP(16'h117EB,4);
TASK_PP(16'h117EC,4);
TASK_PP(16'h117ED,4);
TASK_PP(16'h117EE,4);
TASK_PP(16'h117EF,4);
TASK_PP(16'h117F0,4);
TASK_PP(16'h117F1,4);
TASK_PP(16'h117F2,4);
TASK_PP(16'h117F3,4);
TASK_PP(16'h117F4,4);
TASK_PP(16'h117F5,4);
TASK_PP(16'h117F6,4);
TASK_PP(16'h117F7,4);
TASK_PP(16'h117F8,4);
TASK_PP(16'h117F9,4);
TASK_PP(16'h117FA,4);
TASK_PP(16'h117FB,4);
TASK_PP(16'h117FC,4);
TASK_PP(16'h117FD,4);
TASK_PP(16'h117FE,4);
TASK_PP(16'h117FF,4);
TASK_PP(16'h11800,4);
TASK_PP(16'h11801,4);
TASK_PP(16'h11802,4);
TASK_PP(16'h11803,4);
TASK_PP(16'h11804,4);
TASK_PP(16'h11805,4);
TASK_PP(16'h11806,4);
TASK_PP(16'h11807,4);
TASK_PP(16'h11808,4);
TASK_PP(16'h11809,4);
TASK_PP(16'h1180A,4);
TASK_PP(16'h1180B,4);
TASK_PP(16'h1180C,4);
TASK_PP(16'h1180D,4);
TASK_PP(16'h1180E,4);
TASK_PP(16'h1180F,4);
TASK_PP(16'h11810,4);
TASK_PP(16'h11811,4);
TASK_PP(16'h11812,4);
TASK_PP(16'h11813,4);
TASK_PP(16'h11814,4);
TASK_PP(16'h11815,4);
TASK_PP(16'h11816,4);
TASK_PP(16'h11817,4);
TASK_PP(16'h11818,4);
TASK_PP(16'h11819,4);
TASK_PP(16'h1181A,4);
TASK_PP(16'h1181B,4);
TASK_PP(16'h1181C,4);
TASK_PP(16'h1181D,4);
TASK_PP(16'h1181E,4);
TASK_PP(16'h1181F,4);
TASK_PP(16'h11820,4);
TASK_PP(16'h11821,4);
TASK_PP(16'h11822,4);
TASK_PP(16'h11823,4);
TASK_PP(16'h11824,4);
TASK_PP(16'h11825,4);
TASK_PP(16'h11826,4);
TASK_PP(16'h11827,4);
TASK_PP(16'h11828,4);
TASK_PP(16'h11829,4);
TASK_PP(16'h1182A,4);
TASK_PP(16'h1182B,4);
TASK_PP(16'h1182C,4);
TASK_PP(16'h1182D,4);
TASK_PP(16'h1182E,4);
TASK_PP(16'h1182F,4);
TASK_PP(16'h11830,4);
TASK_PP(16'h11831,4);
TASK_PP(16'h11832,4);
TASK_PP(16'h11833,4);
TASK_PP(16'h11834,4);
TASK_PP(16'h11835,4);
TASK_PP(16'h11836,4);
TASK_PP(16'h11837,4);
TASK_PP(16'h11838,4);
TASK_PP(16'h11839,4);
TASK_PP(16'h1183A,4);
TASK_PP(16'h1183B,4);
TASK_PP(16'h1183C,4);
TASK_PP(16'h1183D,4);
TASK_PP(16'h1183E,4);
TASK_PP(16'h1183F,4);
TASK_PP(16'h11840,4);
TASK_PP(16'h11841,4);
TASK_PP(16'h11842,4);
TASK_PP(16'h11843,4);
TASK_PP(16'h11844,4);
TASK_PP(16'h11845,4);
TASK_PP(16'h11846,4);
TASK_PP(16'h11847,4);
TASK_PP(16'h11848,4);
TASK_PP(16'h11849,4);
TASK_PP(16'h1184A,4);
TASK_PP(16'h1184B,4);
TASK_PP(16'h1184C,4);
TASK_PP(16'h1184D,4);
TASK_PP(16'h1184E,4);
TASK_PP(16'h1184F,4);
TASK_PP(16'h11850,4);
TASK_PP(16'h11851,4);
TASK_PP(16'h11852,4);
TASK_PP(16'h11853,4);
TASK_PP(16'h11854,4);
TASK_PP(16'h11855,4);
TASK_PP(16'h11856,4);
TASK_PP(16'h11857,4);
TASK_PP(16'h11858,4);
TASK_PP(16'h11859,4);
TASK_PP(16'h1185A,4);
TASK_PP(16'h1185B,4);
TASK_PP(16'h1185C,4);
TASK_PP(16'h1185D,4);
TASK_PP(16'h1185E,4);
TASK_PP(16'h1185F,4);
TASK_PP(16'h11860,4);
TASK_PP(16'h11861,4);
TASK_PP(16'h11862,4);
TASK_PP(16'h11863,4);
TASK_PP(16'h11864,4);
TASK_PP(16'h11865,4);
TASK_PP(16'h11866,4);
TASK_PP(16'h11867,4);
TASK_PP(16'h11868,4);
TASK_PP(16'h11869,4);
TASK_PP(16'h1186A,4);
TASK_PP(16'h1186B,4);
TASK_PP(16'h1186C,4);
TASK_PP(16'h1186D,4);
TASK_PP(16'h1186E,4);
TASK_PP(16'h1186F,4);
TASK_PP(16'h11870,4);
TASK_PP(16'h11871,4);
TASK_PP(16'h11872,4);
TASK_PP(16'h11873,4);
TASK_PP(16'h11874,4);
TASK_PP(16'h11875,4);
TASK_PP(16'h11876,4);
TASK_PP(16'h11877,4);
TASK_PP(16'h11878,4);
TASK_PP(16'h11879,4);
TASK_PP(16'h1187A,4);
TASK_PP(16'h1187B,4);
TASK_PP(16'h1187C,4);
TASK_PP(16'h1187D,4);
TASK_PP(16'h1187E,4);
TASK_PP(16'h1187F,4);
TASK_PP(16'h11880,4);
TASK_PP(16'h11881,4);
TASK_PP(16'h11882,4);
TASK_PP(16'h11883,4);
TASK_PP(16'h11884,4);
TASK_PP(16'h11885,4);
TASK_PP(16'h11886,4);
TASK_PP(16'h11887,4);
TASK_PP(16'h11888,4);
TASK_PP(16'h11889,4);
TASK_PP(16'h1188A,4);
TASK_PP(16'h1188B,4);
TASK_PP(16'h1188C,4);
TASK_PP(16'h1188D,4);
TASK_PP(16'h1188E,4);
TASK_PP(16'h1188F,4);
TASK_PP(16'h11890,4);
TASK_PP(16'h11891,4);
TASK_PP(16'h11892,4);
TASK_PP(16'h11893,4);
TASK_PP(16'h11894,4);
TASK_PP(16'h11895,4);
TASK_PP(16'h11896,4);
TASK_PP(16'h11897,4);
TASK_PP(16'h11898,4);
TASK_PP(16'h11899,4);
TASK_PP(16'h1189A,4);
TASK_PP(16'h1189B,4);
TASK_PP(16'h1189C,4);
TASK_PP(16'h1189D,4);
TASK_PP(16'h1189E,4);
TASK_PP(16'h1189F,4);
TASK_PP(16'h118A0,4);
TASK_PP(16'h118A1,4);
TASK_PP(16'h118A2,4);
TASK_PP(16'h118A3,4);
TASK_PP(16'h118A4,4);
TASK_PP(16'h118A5,4);
TASK_PP(16'h118A6,4);
TASK_PP(16'h118A7,4);
TASK_PP(16'h118A8,4);
TASK_PP(16'h118A9,4);
TASK_PP(16'h118AA,4);
TASK_PP(16'h118AB,4);
TASK_PP(16'h118AC,4);
TASK_PP(16'h118AD,4);
TASK_PP(16'h118AE,4);
TASK_PP(16'h118AF,4);
TASK_PP(16'h118B0,4);
TASK_PP(16'h118B1,4);
TASK_PP(16'h118B2,4);
TASK_PP(16'h118B3,4);
TASK_PP(16'h118B4,4);
TASK_PP(16'h118B5,4);
TASK_PP(16'h118B6,4);
TASK_PP(16'h118B7,4);
TASK_PP(16'h118B8,4);
TASK_PP(16'h118B9,4);
TASK_PP(16'h118BA,4);
TASK_PP(16'h118BB,4);
TASK_PP(16'h118BC,4);
TASK_PP(16'h118BD,4);
TASK_PP(16'h118BE,4);
TASK_PP(16'h118BF,4);
TASK_PP(16'h118C0,4);
TASK_PP(16'h118C1,4);
TASK_PP(16'h118C2,4);
TASK_PP(16'h118C3,4);
TASK_PP(16'h118C4,4);
TASK_PP(16'h118C5,4);
TASK_PP(16'h118C6,4);
TASK_PP(16'h118C7,4);
TASK_PP(16'h118C8,4);
TASK_PP(16'h118C9,4);
TASK_PP(16'h118CA,4);
TASK_PP(16'h118CB,4);
TASK_PP(16'h118CC,4);
TASK_PP(16'h118CD,4);
TASK_PP(16'h118CE,4);
TASK_PP(16'h118CF,4);
TASK_PP(16'h118D0,4);
TASK_PP(16'h118D1,4);
TASK_PP(16'h118D2,4);
TASK_PP(16'h118D3,4);
TASK_PP(16'h118D4,4);
TASK_PP(16'h118D5,4);
TASK_PP(16'h118D6,4);
TASK_PP(16'h118D7,4);
TASK_PP(16'h118D8,4);
TASK_PP(16'h118D9,4);
TASK_PP(16'h118DA,4);
TASK_PP(16'h118DB,4);
TASK_PP(16'h118DC,4);
TASK_PP(16'h118DD,4);
TASK_PP(16'h118DE,4);
TASK_PP(16'h118DF,4);
TASK_PP(16'h118E0,4);
TASK_PP(16'h118E1,4);
TASK_PP(16'h118E2,4);
TASK_PP(16'h118E3,4);
TASK_PP(16'h118E4,4);
TASK_PP(16'h118E5,4);
TASK_PP(16'h118E6,4);
TASK_PP(16'h118E7,4);
TASK_PP(16'h118E8,4);
TASK_PP(16'h118E9,4);
TASK_PP(16'h118EA,4);
TASK_PP(16'h118EB,4);
TASK_PP(16'h118EC,4);
TASK_PP(16'h118ED,4);
TASK_PP(16'h118EE,4);
TASK_PP(16'h118EF,4);
TASK_PP(16'h118F0,4);
TASK_PP(16'h118F1,4);
TASK_PP(16'h118F2,4);
TASK_PP(16'h118F3,4);
TASK_PP(16'h118F4,4);
TASK_PP(16'h118F5,4);
TASK_PP(16'h118F6,4);
TASK_PP(16'h118F7,4);
TASK_PP(16'h118F8,4);
TASK_PP(16'h118F9,4);
TASK_PP(16'h118FA,4);
TASK_PP(16'h118FB,4);
TASK_PP(16'h118FC,4);
TASK_PP(16'h118FD,4);
TASK_PP(16'h118FE,4);
TASK_PP(16'h118FF,4);
TASK_PP(16'h11900,4);
TASK_PP(16'h11901,4);
TASK_PP(16'h11902,4);
TASK_PP(16'h11903,4);
TASK_PP(16'h11904,4);
TASK_PP(16'h11905,4);
TASK_PP(16'h11906,4);
TASK_PP(16'h11907,4);
TASK_PP(16'h11908,4);
TASK_PP(16'h11909,4);
TASK_PP(16'h1190A,4);
TASK_PP(16'h1190B,4);
TASK_PP(16'h1190C,4);
TASK_PP(16'h1190D,4);
TASK_PP(16'h1190E,4);
TASK_PP(16'h1190F,4);
TASK_PP(16'h11910,4);
TASK_PP(16'h11911,4);
TASK_PP(16'h11912,4);
TASK_PP(16'h11913,4);
TASK_PP(16'h11914,4);
TASK_PP(16'h11915,4);
TASK_PP(16'h11916,4);
TASK_PP(16'h11917,4);
TASK_PP(16'h11918,4);
TASK_PP(16'h11919,4);
TASK_PP(16'h1191A,4);
TASK_PP(16'h1191B,4);
TASK_PP(16'h1191C,4);
TASK_PP(16'h1191D,4);
TASK_PP(16'h1191E,4);
TASK_PP(16'h1191F,4);
TASK_PP(16'h11920,4);
TASK_PP(16'h11921,4);
TASK_PP(16'h11922,4);
TASK_PP(16'h11923,4);
TASK_PP(16'h11924,4);
TASK_PP(16'h11925,4);
TASK_PP(16'h11926,4);
TASK_PP(16'h11927,4);
TASK_PP(16'h11928,4);
TASK_PP(16'h11929,4);
TASK_PP(16'h1192A,4);
TASK_PP(16'h1192B,4);
TASK_PP(16'h1192C,4);
TASK_PP(16'h1192D,4);
TASK_PP(16'h1192E,4);
TASK_PP(16'h1192F,4);
TASK_PP(16'h11930,4);
TASK_PP(16'h11931,4);
TASK_PP(16'h11932,4);
TASK_PP(16'h11933,4);
TASK_PP(16'h11934,4);
TASK_PP(16'h11935,4);
TASK_PP(16'h11936,4);
TASK_PP(16'h11937,4);
TASK_PP(16'h11938,4);
TASK_PP(16'h11939,4);
TASK_PP(16'h1193A,4);
TASK_PP(16'h1193B,4);
TASK_PP(16'h1193C,4);
TASK_PP(16'h1193D,4);
TASK_PP(16'h1193E,4);
TASK_PP(16'h1193F,4);
TASK_PP(16'h11940,4);
TASK_PP(16'h11941,4);
TASK_PP(16'h11942,4);
TASK_PP(16'h11943,4);
TASK_PP(16'h11944,4);
TASK_PP(16'h11945,4);
TASK_PP(16'h11946,4);
TASK_PP(16'h11947,4);
TASK_PP(16'h11948,4);
TASK_PP(16'h11949,4);
TASK_PP(16'h1194A,4);
TASK_PP(16'h1194B,4);
TASK_PP(16'h1194C,4);
TASK_PP(16'h1194D,4);
TASK_PP(16'h1194E,4);
TASK_PP(16'h1194F,4);
TASK_PP(16'h11950,4);
TASK_PP(16'h11951,4);
TASK_PP(16'h11952,4);
TASK_PP(16'h11953,4);
TASK_PP(16'h11954,4);
TASK_PP(16'h11955,4);
TASK_PP(16'h11956,4);
TASK_PP(16'h11957,4);
TASK_PP(16'h11958,4);
TASK_PP(16'h11959,4);
TASK_PP(16'h1195A,4);
TASK_PP(16'h1195B,4);
TASK_PP(16'h1195C,4);
TASK_PP(16'h1195D,4);
TASK_PP(16'h1195E,4);
TASK_PP(16'h1195F,4);
TASK_PP(16'h11960,4);
TASK_PP(16'h11961,4);
TASK_PP(16'h11962,4);
TASK_PP(16'h11963,4);
TASK_PP(16'h11964,4);
TASK_PP(16'h11965,4);
TASK_PP(16'h11966,4);
TASK_PP(16'h11967,4);
TASK_PP(16'h11968,4);
TASK_PP(16'h11969,4);
TASK_PP(16'h1196A,4);
TASK_PP(16'h1196B,4);
TASK_PP(16'h1196C,4);
TASK_PP(16'h1196D,4);
TASK_PP(16'h1196E,4);
TASK_PP(16'h1196F,4);
TASK_PP(16'h11970,4);
TASK_PP(16'h11971,4);
TASK_PP(16'h11972,4);
TASK_PP(16'h11973,4);
TASK_PP(16'h11974,4);
TASK_PP(16'h11975,4);
TASK_PP(16'h11976,4);
TASK_PP(16'h11977,4);
TASK_PP(16'h11978,4);
TASK_PP(16'h11979,4);
TASK_PP(16'h1197A,4);
TASK_PP(16'h1197B,4);
TASK_PP(16'h1197C,4);
TASK_PP(16'h1197D,4);
TASK_PP(16'h1197E,4);
TASK_PP(16'h1197F,4);
TASK_PP(16'h11980,4);
TASK_PP(16'h11981,4);
TASK_PP(16'h11982,4);
TASK_PP(16'h11983,4);
TASK_PP(16'h11984,4);
TASK_PP(16'h11985,4);
TASK_PP(16'h11986,4);
TASK_PP(16'h11987,4);
TASK_PP(16'h11988,4);
TASK_PP(16'h11989,4);
TASK_PP(16'h1198A,4);
TASK_PP(16'h1198B,4);
TASK_PP(16'h1198C,4);
TASK_PP(16'h1198D,4);
TASK_PP(16'h1198E,4);
TASK_PP(16'h1198F,4);
TASK_PP(16'h11990,4);
TASK_PP(16'h11991,4);
TASK_PP(16'h11992,4);
TASK_PP(16'h11993,4);
TASK_PP(16'h11994,4);
TASK_PP(16'h11995,4);
TASK_PP(16'h11996,4);
TASK_PP(16'h11997,4);
TASK_PP(16'h11998,4);
TASK_PP(16'h11999,4);
TASK_PP(16'h1199A,4);
TASK_PP(16'h1199B,4);
TASK_PP(16'h1199C,4);
TASK_PP(16'h1199D,4);
TASK_PP(16'h1199E,4);
TASK_PP(16'h1199F,4);
TASK_PP(16'h119A0,4);
TASK_PP(16'h119A1,4);
TASK_PP(16'h119A2,4);
TASK_PP(16'h119A3,4);
TASK_PP(16'h119A4,4);
TASK_PP(16'h119A5,4);
TASK_PP(16'h119A6,4);
TASK_PP(16'h119A7,4);
TASK_PP(16'h119A8,4);
TASK_PP(16'h119A9,4);
TASK_PP(16'h119AA,4);
TASK_PP(16'h119AB,4);
TASK_PP(16'h119AC,4);
TASK_PP(16'h119AD,4);
TASK_PP(16'h119AE,4);
TASK_PP(16'h119AF,4);
TASK_PP(16'h119B0,4);
TASK_PP(16'h119B1,4);
TASK_PP(16'h119B2,4);
TASK_PP(16'h119B3,4);
TASK_PP(16'h119B4,4);
TASK_PP(16'h119B5,4);
TASK_PP(16'h119B6,4);
TASK_PP(16'h119B7,4);
TASK_PP(16'h119B8,4);
TASK_PP(16'h119B9,4);
TASK_PP(16'h119BA,4);
TASK_PP(16'h119BB,4);
TASK_PP(16'h119BC,4);
TASK_PP(16'h119BD,4);
TASK_PP(16'h119BE,4);
TASK_PP(16'h119BF,4);
TASK_PP(16'h119C0,4);
TASK_PP(16'h119C1,4);
TASK_PP(16'h119C2,4);
TASK_PP(16'h119C3,4);
TASK_PP(16'h119C4,4);
TASK_PP(16'h119C5,4);
TASK_PP(16'h119C6,4);
TASK_PP(16'h119C7,4);
TASK_PP(16'h119C8,4);
TASK_PP(16'h119C9,4);
TASK_PP(16'h119CA,4);
TASK_PP(16'h119CB,4);
TASK_PP(16'h119CC,4);
TASK_PP(16'h119CD,4);
TASK_PP(16'h119CE,4);
TASK_PP(16'h119CF,4);
TASK_PP(16'h119D0,4);
TASK_PP(16'h119D1,4);
TASK_PP(16'h119D2,4);
TASK_PP(16'h119D3,4);
TASK_PP(16'h119D4,4);
TASK_PP(16'h119D5,4);
TASK_PP(16'h119D6,4);
TASK_PP(16'h119D7,4);
TASK_PP(16'h119D8,4);
TASK_PP(16'h119D9,4);
TASK_PP(16'h119DA,4);
TASK_PP(16'h119DB,4);
TASK_PP(16'h119DC,4);
TASK_PP(16'h119DD,4);
TASK_PP(16'h119DE,4);
TASK_PP(16'h119DF,4);
TASK_PP(16'h119E0,4);
TASK_PP(16'h119E1,4);
TASK_PP(16'h119E2,4);
TASK_PP(16'h119E3,4);
TASK_PP(16'h119E4,4);
TASK_PP(16'h119E5,4);
TASK_PP(16'h119E6,4);
TASK_PP(16'h119E7,4);
TASK_PP(16'h119E8,4);
TASK_PP(16'h119E9,4);
TASK_PP(16'h119EA,4);
TASK_PP(16'h119EB,4);
TASK_PP(16'h119EC,4);
TASK_PP(16'h119ED,4);
TASK_PP(16'h119EE,4);
TASK_PP(16'h119EF,4);
TASK_PP(16'h119F0,4);
TASK_PP(16'h119F1,4);
TASK_PP(16'h119F2,4);
TASK_PP(16'h119F3,4);
TASK_PP(16'h119F4,4);
TASK_PP(16'h119F5,4);
TASK_PP(16'h119F6,4);
TASK_PP(16'h119F7,4);
TASK_PP(16'h119F8,4);
TASK_PP(16'h119F9,4);
TASK_PP(16'h119FA,4);
TASK_PP(16'h119FB,4);
TASK_PP(16'h119FC,4);
TASK_PP(16'h119FD,4);
TASK_PP(16'h119FE,4);
TASK_PP(16'h119FF,4);
TASK_PP(16'h11A00,4);
TASK_PP(16'h11A01,4);
TASK_PP(16'h11A02,4);
TASK_PP(16'h11A03,4);
TASK_PP(16'h11A04,4);
TASK_PP(16'h11A05,4);
TASK_PP(16'h11A06,4);
TASK_PP(16'h11A07,4);
TASK_PP(16'h11A08,4);
TASK_PP(16'h11A09,4);
TASK_PP(16'h11A0A,4);
TASK_PP(16'h11A0B,4);
TASK_PP(16'h11A0C,4);
TASK_PP(16'h11A0D,4);
TASK_PP(16'h11A0E,4);
TASK_PP(16'h11A0F,4);
TASK_PP(16'h11A10,4);
TASK_PP(16'h11A11,4);
TASK_PP(16'h11A12,4);
TASK_PP(16'h11A13,4);
TASK_PP(16'h11A14,4);
TASK_PP(16'h11A15,4);
TASK_PP(16'h11A16,4);
TASK_PP(16'h11A17,4);
TASK_PP(16'h11A18,4);
TASK_PP(16'h11A19,4);
TASK_PP(16'h11A1A,4);
TASK_PP(16'h11A1B,4);
TASK_PP(16'h11A1C,4);
TASK_PP(16'h11A1D,4);
TASK_PP(16'h11A1E,4);
TASK_PP(16'h11A1F,4);
TASK_PP(16'h11A20,4);
TASK_PP(16'h11A21,4);
TASK_PP(16'h11A22,4);
TASK_PP(16'h11A23,4);
TASK_PP(16'h11A24,4);
TASK_PP(16'h11A25,4);
TASK_PP(16'h11A26,4);
TASK_PP(16'h11A27,4);
TASK_PP(16'h11A28,4);
TASK_PP(16'h11A29,4);
TASK_PP(16'h11A2A,4);
TASK_PP(16'h11A2B,4);
TASK_PP(16'h11A2C,4);
TASK_PP(16'h11A2D,4);
TASK_PP(16'h11A2E,4);
TASK_PP(16'h11A2F,4);
TASK_PP(16'h11A30,4);
TASK_PP(16'h11A31,4);
TASK_PP(16'h11A32,4);
TASK_PP(16'h11A33,4);
TASK_PP(16'h11A34,4);
TASK_PP(16'h11A35,4);
TASK_PP(16'h11A36,4);
TASK_PP(16'h11A37,4);
TASK_PP(16'h11A38,4);
TASK_PP(16'h11A39,4);
TASK_PP(16'h11A3A,4);
TASK_PP(16'h11A3B,4);
TASK_PP(16'h11A3C,4);
TASK_PP(16'h11A3D,4);
TASK_PP(16'h11A3E,4);
TASK_PP(16'h11A3F,4);
TASK_PP(16'h11A40,4);
TASK_PP(16'h11A41,4);
TASK_PP(16'h11A42,4);
TASK_PP(16'h11A43,4);
TASK_PP(16'h11A44,4);
TASK_PP(16'h11A45,4);
TASK_PP(16'h11A46,4);
TASK_PP(16'h11A47,4);
TASK_PP(16'h11A48,4);
TASK_PP(16'h11A49,4);
TASK_PP(16'h11A4A,4);
TASK_PP(16'h11A4B,4);
TASK_PP(16'h11A4C,4);
TASK_PP(16'h11A4D,4);
TASK_PP(16'h11A4E,4);
TASK_PP(16'h11A4F,4);
TASK_PP(16'h11A50,4);
TASK_PP(16'h11A51,4);
TASK_PP(16'h11A52,4);
TASK_PP(16'h11A53,4);
TASK_PP(16'h11A54,4);
TASK_PP(16'h11A55,4);
TASK_PP(16'h11A56,4);
TASK_PP(16'h11A57,4);
TASK_PP(16'h11A58,4);
TASK_PP(16'h11A59,4);
TASK_PP(16'h11A5A,4);
TASK_PP(16'h11A5B,4);
TASK_PP(16'h11A5C,4);
TASK_PP(16'h11A5D,4);
TASK_PP(16'h11A5E,4);
TASK_PP(16'h11A5F,4);
TASK_PP(16'h11A60,4);
TASK_PP(16'h11A61,4);
TASK_PP(16'h11A62,4);
TASK_PP(16'h11A63,4);
TASK_PP(16'h11A64,4);
TASK_PP(16'h11A65,4);
TASK_PP(16'h11A66,4);
TASK_PP(16'h11A67,4);
TASK_PP(16'h11A68,4);
TASK_PP(16'h11A69,4);
TASK_PP(16'h11A6A,4);
TASK_PP(16'h11A6B,4);
TASK_PP(16'h11A6C,4);
TASK_PP(16'h11A6D,4);
TASK_PP(16'h11A6E,4);
TASK_PP(16'h11A6F,4);
TASK_PP(16'h11A70,4);
TASK_PP(16'h11A71,4);
TASK_PP(16'h11A72,4);
TASK_PP(16'h11A73,4);
TASK_PP(16'h11A74,4);
TASK_PP(16'h11A75,4);
TASK_PP(16'h11A76,4);
TASK_PP(16'h11A77,4);
TASK_PP(16'h11A78,4);
TASK_PP(16'h11A79,4);
TASK_PP(16'h11A7A,4);
TASK_PP(16'h11A7B,4);
TASK_PP(16'h11A7C,4);
TASK_PP(16'h11A7D,4);
TASK_PP(16'h11A7E,4);
TASK_PP(16'h11A7F,4);
TASK_PP(16'h11A80,4);
TASK_PP(16'h11A81,4);
TASK_PP(16'h11A82,4);
TASK_PP(16'h11A83,4);
TASK_PP(16'h11A84,4);
TASK_PP(16'h11A85,4);
TASK_PP(16'h11A86,4);
TASK_PP(16'h11A87,4);
TASK_PP(16'h11A88,4);
TASK_PP(16'h11A89,4);
TASK_PP(16'h11A8A,4);
TASK_PP(16'h11A8B,4);
TASK_PP(16'h11A8C,4);
TASK_PP(16'h11A8D,4);
TASK_PP(16'h11A8E,4);
TASK_PP(16'h11A8F,4);
TASK_PP(16'h11A90,4);
TASK_PP(16'h11A91,4);
TASK_PP(16'h11A92,4);
TASK_PP(16'h11A93,4);
TASK_PP(16'h11A94,4);
TASK_PP(16'h11A95,4);
TASK_PP(16'h11A96,4);
TASK_PP(16'h11A97,4);
TASK_PP(16'h11A98,4);
TASK_PP(16'h11A99,4);
TASK_PP(16'h11A9A,4);
TASK_PP(16'h11A9B,4);
TASK_PP(16'h11A9C,4);
TASK_PP(16'h11A9D,4);
TASK_PP(16'h11A9E,4);
TASK_PP(16'h11A9F,4);
TASK_PP(16'h11AA0,4);
TASK_PP(16'h11AA1,4);
TASK_PP(16'h11AA2,4);
TASK_PP(16'h11AA3,4);
TASK_PP(16'h11AA4,4);
TASK_PP(16'h11AA5,4);
TASK_PP(16'h11AA6,4);
TASK_PP(16'h11AA7,4);
TASK_PP(16'h11AA8,4);
TASK_PP(16'h11AA9,4);
TASK_PP(16'h11AAA,4);
TASK_PP(16'h11AAB,4);
TASK_PP(16'h11AAC,4);
TASK_PP(16'h11AAD,4);
TASK_PP(16'h11AAE,4);
TASK_PP(16'h11AAF,4);
TASK_PP(16'h11AB0,4);
TASK_PP(16'h11AB1,4);
TASK_PP(16'h11AB2,4);
TASK_PP(16'h11AB3,4);
TASK_PP(16'h11AB4,4);
TASK_PP(16'h11AB5,4);
TASK_PP(16'h11AB6,4);
TASK_PP(16'h11AB7,4);
TASK_PP(16'h11AB8,4);
TASK_PP(16'h11AB9,4);
TASK_PP(16'h11ABA,4);
TASK_PP(16'h11ABB,4);
TASK_PP(16'h11ABC,4);
TASK_PP(16'h11ABD,4);
TASK_PP(16'h11ABE,4);
TASK_PP(16'h11ABF,4);
TASK_PP(16'h11AC0,4);
TASK_PP(16'h11AC1,4);
TASK_PP(16'h11AC2,4);
TASK_PP(16'h11AC3,4);
TASK_PP(16'h11AC4,4);
TASK_PP(16'h11AC5,4);
TASK_PP(16'h11AC6,4);
TASK_PP(16'h11AC7,4);
TASK_PP(16'h11AC8,4);
TASK_PP(16'h11AC9,4);
TASK_PP(16'h11ACA,4);
TASK_PP(16'h11ACB,4);
TASK_PP(16'h11ACC,4);
TASK_PP(16'h11ACD,4);
TASK_PP(16'h11ACE,4);
TASK_PP(16'h11ACF,4);
TASK_PP(16'h11AD0,4);
TASK_PP(16'h11AD1,4);
TASK_PP(16'h11AD2,4);
TASK_PP(16'h11AD3,4);
TASK_PP(16'h11AD4,4);
TASK_PP(16'h11AD5,4);
TASK_PP(16'h11AD6,4);
TASK_PP(16'h11AD7,4);
TASK_PP(16'h11AD8,4);
TASK_PP(16'h11AD9,4);
TASK_PP(16'h11ADA,4);
TASK_PP(16'h11ADB,4);
TASK_PP(16'h11ADC,4);
TASK_PP(16'h11ADD,4);
TASK_PP(16'h11ADE,4);
TASK_PP(16'h11ADF,4);
TASK_PP(16'h11AE0,4);
TASK_PP(16'h11AE1,4);
TASK_PP(16'h11AE2,4);
TASK_PP(16'h11AE3,4);
TASK_PP(16'h11AE4,4);
TASK_PP(16'h11AE5,4);
TASK_PP(16'h11AE6,4);
TASK_PP(16'h11AE7,4);
TASK_PP(16'h11AE8,4);
TASK_PP(16'h11AE9,4);
TASK_PP(16'h11AEA,4);
TASK_PP(16'h11AEB,4);
TASK_PP(16'h11AEC,4);
TASK_PP(16'h11AED,4);
TASK_PP(16'h11AEE,4);
TASK_PP(16'h11AEF,4);
TASK_PP(16'h11AF0,4);
TASK_PP(16'h11AF1,4);
TASK_PP(16'h11AF2,4);
TASK_PP(16'h11AF3,4);
TASK_PP(16'h11AF4,4);
TASK_PP(16'h11AF5,4);
TASK_PP(16'h11AF6,4);
TASK_PP(16'h11AF7,4);
TASK_PP(16'h11AF8,4);
TASK_PP(16'h11AF9,4);
TASK_PP(16'h11AFA,4);
TASK_PP(16'h11AFB,4);
TASK_PP(16'h11AFC,4);
TASK_PP(16'h11AFD,4);
TASK_PP(16'h11AFE,4);
TASK_PP(16'h11AFF,4);
TASK_PP(16'h11B00,4);
TASK_PP(16'h11B01,4);
TASK_PP(16'h11B02,4);
TASK_PP(16'h11B03,4);
TASK_PP(16'h11B04,4);
TASK_PP(16'h11B05,4);
TASK_PP(16'h11B06,4);
TASK_PP(16'h11B07,4);
TASK_PP(16'h11B08,4);
TASK_PP(16'h11B09,4);
TASK_PP(16'h11B0A,4);
TASK_PP(16'h11B0B,4);
TASK_PP(16'h11B0C,4);
TASK_PP(16'h11B0D,4);
TASK_PP(16'h11B0E,4);
TASK_PP(16'h11B0F,4);
TASK_PP(16'h11B10,4);
TASK_PP(16'h11B11,4);
TASK_PP(16'h11B12,4);
TASK_PP(16'h11B13,4);
TASK_PP(16'h11B14,4);
TASK_PP(16'h11B15,4);
TASK_PP(16'h11B16,4);
TASK_PP(16'h11B17,4);
TASK_PP(16'h11B18,4);
TASK_PP(16'h11B19,4);
TASK_PP(16'h11B1A,4);
TASK_PP(16'h11B1B,4);
TASK_PP(16'h11B1C,4);
TASK_PP(16'h11B1D,4);
TASK_PP(16'h11B1E,4);
TASK_PP(16'h11B1F,4);
TASK_PP(16'h11B20,4);
TASK_PP(16'h11B21,4);
TASK_PP(16'h11B22,4);
TASK_PP(16'h11B23,4);
TASK_PP(16'h11B24,4);
TASK_PP(16'h11B25,4);
TASK_PP(16'h11B26,4);
TASK_PP(16'h11B27,4);
TASK_PP(16'h11B28,4);
TASK_PP(16'h11B29,4);
TASK_PP(16'h11B2A,4);
TASK_PP(16'h11B2B,4);
TASK_PP(16'h11B2C,4);
TASK_PP(16'h11B2D,4);
TASK_PP(16'h11B2E,4);
TASK_PP(16'h11B2F,4);
TASK_PP(16'h11B30,4);
TASK_PP(16'h11B31,4);
TASK_PP(16'h11B32,4);
TASK_PP(16'h11B33,4);
TASK_PP(16'h11B34,4);
TASK_PP(16'h11B35,4);
TASK_PP(16'h11B36,4);
TASK_PP(16'h11B37,4);
TASK_PP(16'h11B38,4);
TASK_PP(16'h11B39,4);
TASK_PP(16'h11B3A,4);
TASK_PP(16'h11B3B,4);
TASK_PP(16'h11B3C,4);
TASK_PP(16'h11B3D,4);
TASK_PP(16'h11B3E,4);
TASK_PP(16'h11B3F,4);
TASK_PP(16'h11B40,4);
TASK_PP(16'h11B41,4);
TASK_PP(16'h11B42,4);
TASK_PP(16'h11B43,4);
TASK_PP(16'h11B44,4);
TASK_PP(16'h11B45,4);
TASK_PP(16'h11B46,4);
TASK_PP(16'h11B47,4);
TASK_PP(16'h11B48,4);
TASK_PP(16'h11B49,4);
TASK_PP(16'h11B4A,4);
TASK_PP(16'h11B4B,4);
TASK_PP(16'h11B4C,4);
TASK_PP(16'h11B4D,4);
TASK_PP(16'h11B4E,4);
TASK_PP(16'h11B4F,4);
TASK_PP(16'h11B50,4);
TASK_PP(16'h11B51,4);
TASK_PP(16'h11B52,4);
TASK_PP(16'h11B53,4);
TASK_PP(16'h11B54,4);
TASK_PP(16'h11B55,4);
TASK_PP(16'h11B56,4);
TASK_PP(16'h11B57,4);
TASK_PP(16'h11B58,4);
TASK_PP(16'h11B59,4);
TASK_PP(16'h11B5A,4);
TASK_PP(16'h11B5B,4);
TASK_PP(16'h11B5C,4);
TASK_PP(16'h11B5D,4);
TASK_PP(16'h11B5E,4);
TASK_PP(16'h11B5F,4);
TASK_PP(16'h11B60,4);
TASK_PP(16'h11B61,4);
TASK_PP(16'h11B62,4);
TASK_PP(16'h11B63,4);
TASK_PP(16'h11B64,4);
TASK_PP(16'h11B65,4);
TASK_PP(16'h11B66,4);
TASK_PP(16'h11B67,4);
TASK_PP(16'h11B68,4);
TASK_PP(16'h11B69,4);
TASK_PP(16'h11B6A,4);
TASK_PP(16'h11B6B,4);
TASK_PP(16'h11B6C,4);
TASK_PP(16'h11B6D,4);
TASK_PP(16'h11B6E,4);
TASK_PP(16'h11B6F,4);
TASK_PP(16'h11B70,4);
TASK_PP(16'h11B71,4);
TASK_PP(16'h11B72,4);
TASK_PP(16'h11B73,4);
TASK_PP(16'h11B74,4);
TASK_PP(16'h11B75,4);
TASK_PP(16'h11B76,4);
TASK_PP(16'h11B77,4);
TASK_PP(16'h11B78,4);
TASK_PP(16'h11B79,4);
TASK_PP(16'h11B7A,4);
TASK_PP(16'h11B7B,4);
TASK_PP(16'h11B7C,4);
TASK_PP(16'h11B7D,4);
TASK_PP(16'h11B7E,4);
TASK_PP(16'h11B7F,4);
TASK_PP(16'h11B80,4);
TASK_PP(16'h11B81,4);
TASK_PP(16'h11B82,4);
TASK_PP(16'h11B83,4);
TASK_PP(16'h11B84,4);
TASK_PP(16'h11B85,4);
TASK_PP(16'h11B86,4);
TASK_PP(16'h11B87,4);
TASK_PP(16'h11B88,4);
TASK_PP(16'h11B89,4);
TASK_PP(16'h11B8A,4);
TASK_PP(16'h11B8B,4);
TASK_PP(16'h11B8C,4);
TASK_PP(16'h11B8D,4);
TASK_PP(16'h11B8E,4);
TASK_PP(16'h11B8F,4);
TASK_PP(16'h11B90,4);
TASK_PP(16'h11B91,4);
TASK_PP(16'h11B92,4);
TASK_PP(16'h11B93,4);
TASK_PP(16'h11B94,4);
TASK_PP(16'h11B95,4);
TASK_PP(16'h11B96,4);
TASK_PP(16'h11B97,4);
TASK_PP(16'h11B98,4);
TASK_PP(16'h11B99,4);
TASK_PP(16'h11B9A,4);
TASK_PP(16'h11B9B,4);
TASK_PP(16'h11B9C,4);
TASK_PP(16'h11B9D,4);
TASK_PP(16'h11B9E,4);
TASK_PP(16'h11B9F,4);
TASK_PP(16'h11BA0,4);
TASK_PP(16'h11BA1,4);
TASK_PP(16'h11BA2,4);
TASK_PP(16'h11BA3,4);
TASK_PP(16'h11BA4,4);
TASK_PP(16'h11BA5,4);
TASK_PP(16'h11BA6,4);
TASK_PP(16'h11BA7,4);
TASK_PP(16'h11BA8,4);
TASK_PP(16'h11BA9,4);
TASK_PP(16'h11BAA,4);
TASK_PP(16'h11BAB,4);
TASK_PP(16'h11BAC,4);
TASK_PP(16'h11BAD,4);
TASK_PP(16'h11BAE,4);
TASK_PP(16'h11BAF,4);
TASK_PP(16'h11BB0,4);
TASK_PP(16'h11BB1,4);
TASK_PP(16'h11BB2,4);
TASK_PP(16'h11BB3,4);
TASK_PP(16'h11BB4,4);
TASK_PP(16'h11BB5,4);
TASK_PP(16'h11BB6,4);
TASK_PP(16'h11BB7,4);
TASK_PP(16'h11BB8,4);
TASK_PP(16'h11BB9,4);
TASK_PP(16'h11BBA,4);
TASK_PP(16'h11BBB,4);
TASK_PP(16'h11BBC,4);
TASK_PP(16'h11BBD,4);
TASK_PP(16'h11BBE,4);
TASK_PP(16'h11BBF,4);
TASK_PP(16'h11BC0,4);
TASK_PP(16'h11BC1,4);
TASK_PP(16'h11BC2,4);
TASK_PP(16'h11BC3,4);
TASK_PP(16'h11BC4,4);
TASK_PP(16'h11BC5,4);
TASK_PP(16'h11BC6,4);
TASK_PP(16'h11BC7,4);
TASK_PP(16'h11BC8,4);
TASK_PP(16'h11BC9,4);
TASK_PP(16'h11BCA,4);
TASK_PP(16'h11BCB,4);
TASK_PP(16'h11BCC,4);
TASK_PP(16'h11BCD,4);
TASK_PP(16'h11BCE,4);
TASK_PP(16'h11BCF,4);
TASK_PP(16'h11BD0,4);
TASK_PP(16'h11BD1,4);
TASK_PP(16'h11BD2,4);
TASK_PP(16'h11BD3,4);
TASK_PP(16'h11BD4,4);
TASK_PP(16'h11BD5,4);
TASK_PP(16'h11BD6,4);
TASK_PP(16'h11BD7,4);
TASK_PP(16'h11BD8,4);
TASK_PP(16'h11BD9,4);
TASK_PP(16'h11BDA,4);
TASK_PP(16'h11BDB,4);
TASK_PP(16'h11BDC,4);
TASK_PP(16'h11BDD,4);
TASK_PP(16'h11BDE,4);
TASK_PP(16'h11BDF,4);
TASK_PP(16'h11BE0,4);
TASK_PP(16'h11BE1,4);
TASK_PP(16'h11BE2,4);
TASK_PP(16'h11BE3,4);
TASK_PP(16'h11BE4,4);
TASK_PP(16'h11BE5,4);
TASK_PP(16'h11BE6,4);
TASK_PP(16'h11BE7,4);
TASK_PP(16'h11BE8,4);
TASK_PP(16'h11BE9,4);
TASK_PP(16'h11BEA,4);
TASK_PP(16'h11BEB,4);
TASK_PP(16'h11BEC,4);
TASK_PP(16'h11BED,4);
TASK_PP(16'h11BEE,4);
TASK_PP(16'h11BEF,4);
TASK_PP(16'h11BF0,4);
TASK_PP(16'h11BF1,4);
TASK_PP(16'h11BF2,4);
TASK_PP(16'h11BF3,4);
TASK_PP(16'h11BF4,4);
TASK_PP(16'h11BF5,4);
TASK_PP(16'h11BF6,4);
TASK_PP(16'h11BF7,4);
TASK_PP(16'h11BF8,4);
TASK_PP(16'h11BF9,4);
TASK_PP(16'h11BFA,4);
TASK_PP(16'h11BFB,4);
TASK_PP(16'h11BFC,4);
TASK_PP(16'h11BFD,4);
TASK_PP(16'h11BFE,4);
TASK_PP(16'h11BFF,4);
TASK_PP(16'h11C00,4);
TASK_PP(16'h11C01,4);
TASK_PP(16'h11C02,4);
TASK_PP(16'h11C03,4);
TASK_PP(16'h11C04,4);
TASK_PP(16'h11C05,4);
TASK_PP(16'h11C06,4);
TASK_PP(16'h11C07,4);
TASK_PP(16'h11C08,4);
TASK_PP(16'h11C09,4);
TASK_PP(16'h11C0A,4);
TASK_PP(16'h11C0B,4);
TASK_PP(16'h11C0C,4);
TASK_PP(16'h11C0D,4);
TASK_PP(16'h11C0E,4);
TASK_PP(16'h11C0F,4);
TASK_PP(16'h11C10,4);
TASK_PP(16'h11C11,4);
TASK_PP(16'h11C12,4);
TASK_PP(16'h11C13,4);
TASK_PP(16'h11C14,4);
TASK_PP(16'h11C15,4);
TASK_PP(16'h11C16,4);
TASK_PP(16'h11C17,4);
TASK_PP(16'h11C18,4);
TASK_PP(16'h11C19,4);
TASK_PP(16'h11C1A,4);
TASK_PP(16'h11C1B,4);
TASK_PP(16'h11C1C,4);
TASK_PP(16'h11C1D,4);
TASK_PP(16'h11C1E,4);
TASK_PP(16'h11C1F,4);
TASK_PP(16'h11C20,4);
TASK_PP(16'h11C21,4);
TASK_PP(16'h11C22,4);
TASK_PP(16'h11C23,4);
TASK_PP(16'h11C24,4);
TASK_PP(16'h11C25,4);
TASK_PP(16'h11C26,4);
TASK_PP(16'h11C27,4);
TASK_PP(16'h11C28,4);
TASK_PP(16'h11C29,4);
TASK_PP(16'h11C2A,4);
TASK_PP(16'h11C2B,4);
TASK_PP(16'h11C2C,4);
TASK_PP(16'h11C2D,4);
TASK_PP(16'h11C2E,4);
TASK_PP(16'h11C2F,4);
TASK_PP(16'h11C30,4);
TASK_PP(16'h11C31,4);
TASK_PP(16'h11C32,4);
TASK_PP(16'h11C33,4);
TASK_PP(16'h11C34,4);
TASK_PP(16'h11C35,4);
TASK_PP(16'h11C36,4);
TASK_PP(16'h11C37,4);
TASK_PP(16'h11C38,4);
TASK_PP(16'h11C39,4);
TASK_PP(16'h11C3A,4);
TASK_PP(16'h11C3B,4);
TASK_PP(16'h11C3C,4);
TASK_PP(16'h11C3D,4);
TASK_PP(16'h11C3E,4);
TASK_PP(16'h11C3F,4);
TASK_PP(16'h11C40,4);
TASK_PP(16'h11C41,4);
TASK_PP(16'h11C42,4);
TASK_PP(16'h11C43,4);
TASK_PP(16'h11C44,4);
TASK_PP(16'h11C45,4);
TASK_PP(16'h11C46,4);
TASK_PP(16'h11C47,4);
TASK_PP(16'h11C48,4);
TASK_PP(16'h11C49,4);
TASK_PP(16'h11C4A,4);
TASK_PP(16'h11C4B,4);
TASK_PP(16'h11C4C,4);
TASK_PP(16'h11C4D,4);
TASK_PP(16'h11C4E,4);
TASK_PP(16'h11C4F,4);
TASK_PP(16'h11C50,4);
TASK_PP(16'h11C51,4);
TASK_PP(16'h11C52,4);
TASK_PP(16'h11C53,4);
TASK_PP(16'h11C54,4);
TASK_PP(16'h11C55,4);
TASK_PP(16'h11C56,4);
TASK_PP(16'h11C57,4);
TASK_PP(16'h11C58,4);
TASK_PP(16'h11C59,4);
TASK_PP(16'h11C5A,4);
TASK_PP(16'h11C5B,4);
TASK_PP(16'h11C5C,4);
TASK_PP(16'h11C5D,4);
TASK_PP(16'h11C5E,4);
TASK_PP(16'h11C5F,4);
TASK_PP(16'h11C60,4);
TASK_PP(16'h11C61,4);
TASK_PP(16'h11C62,4);
TASK_PP(16'h11C63,4);
TASK_PP(16'h11C64,4);
TASK_PP(16'h11C65,4);
TASK_PP(16'h11C66,4);
TASK_PP(16'h11C67,4);
TASK_PP(16'h11C68,4);
TASK_PP(16'h11C69,4);
TASK_PP(16'h11C6A,4);
TASK_PP(16'h11C6B,4);
TASK_PP(16'h11C6C,4);
TASK_PP(16'h11C6D,4);
TASK_PP(16'h11C6E,4);
TASK_PP(16'h11C6F,4);
TASK_PP(16'h11C70,4);
TASK_PP(16'h11C71,4);
TASK_PP(16'h11C72,4);
TASK_PP(16'h11C73,4);
TASK_PP(16'h11C74,4);
TASK_PP(16'h11C75,4);
TASK_PP(16'h11C76,4);
TASK_PP(16'h11C77,4);
TASK_PP(16'h11C78,4);
TASK_PP(16'h11C79,4);
TASK_PP(16'h11C7A,4);
TASK_PP(16'h11C7B,4);
TASK_PP(16'h11C7C,4);
TASK_PP(16'h11C7D,4);
TASK_PP(16'h11C7E,4);
TASK_PP(16'h11C7F,4);
TASK_PP(16'h11C80,4);
TASK_PP(16'h11C81,4);
TASK_PP(16'h11C82,4);
TASK_PP(16'h11C83,4);
TASK_PP(16'h11C84,4);
TASK_PP(16'h11C85,4);
TASK_PP(16'h11C86,4);
TASK_PP(16'h11C87,4);
TASK_PP(16'h11C88,4);
TASK_PP(16'h11C89,4);
TASK_PP(16'h11C8A,4);
TASK_PP(16'h11C8B,4);
TASK_PP(16'h11C8C,4);
TASK_PP(16'h11C8D,4);
TASK_PP(16'h11C8E,4);
TASK_PP(16'h11C8F,4);
TASK_PP(16'h11C90,4);
TASK_PP(16'h11C91,4);
TASK_PP(16'h11C92,4);
TASK_PP(16'h11C93,4);
TASK_PP(16'h11C94,4);
TASK_PP(16'h11C95,4);
TASK_PP(16'h11C96,4);
TASK_PP(16'h11C97,4);
TASK_PP(16'h11C98,4);
TASK_PP(16'h11C99,4);
TASK_PP(16'h11C9A,4);
TASK_PP(16'h11C9B,4);
TASK_PP(16'h11C9C,4);
TASK_PP(16'h11C9D,4);
TASK_PP(16'h11C9E,4);
TASK_PP(16'h11C9F,4);
TASK_PP(16'h11CA0,4);
TASK_PP(16'h11CA1,4);
TASK_PP(16'h11CA2,4);
TASK_PP(16'h11CA3,4);
TASK_PP(16'h11CA4,4);
TASK_PP(16'h11CA5,4);
TASK_PP(16'h11CA6,4);
TASK_PP(16'h11CA7,4);
TASK_PP(16'h11CA8,4);
TASK_PP(16'h11CA9,4);
TASK_PP(16'h11CAA,4);
TASK_PP(16'h11CAB,4);
TASK_PP(16'h11CAC,4);
TASK_PP(16'h11CAD,4);
TASK_PP(16'h11CAE,4);
TASK_PP(16'h11CAF,4);
TASK_PP(16'h11CB0,4);
TASK_PP(16'h11CB1,4);
TASK_PP(16'h11CB2,4);
TASK_PP(16'h11CB3,4);
TASK_PP(16'h11CB4,4);
TASK_PP(16'h11CB5,4);
TASK_PP(16'h11CB6,4);
TASK_PP(16'h11CB7,4);
TASK_PP(16'h11CB8,4);
TASK_PP(16'h11CB9,4);
TASK_PP(16'h11CBA,4);
TASK_PP(16'h11CBB,4);
TASK_PP(16'h11CBC,4);
TASK_PP(16'h11CBD,4);
TASK_PP(16'h11CBE,4);
TASK_PP(16'h11CBF,4);
TASK_PP(16'h11CC0,4);
TASK_PP(16'h11CC1,4);
TASK_PP(16'h11CC2,4);
TASK_PP(16'h11CC3,4);
TASK_PP(16'h11CC4,4);
TASK_PP(16'h11CC5,4);
TASK_PP(16'h11CC6,4);
TASK_PP(16'h11CC7,4);
TASK_PP(16'h11CC8,4);
TASK_PP(16'h11CC9,4);
TASK_PP(16'h11CCA,4);
TASK_PP(16'h11CCB,4);
TASK_PP(16'h11CCC,4);
TASK_PP(16'h11CCD,4);
TASK_PP(16'h11CCE,4);
TASK_PP(16'h11CCF,4);
TASK_PP(16'h11CD0,4);
TASK_PP(16'h11CD1,4);
TASK_PP(16'h11CD2,4);
TASK_PP(16'h11CD3,4);
TASK_PP(16'h11CD4,4);
TASK_PP(16'h11CD5,4);
TASK_PP(16'h11CD6,4);
TASK_PP(16'h11CD7,4);
TASK_PP(16'h11CD8,4);
TASK_PP(16'h11CD9,4);
TASK_PP(16'h11CDA,4);
TASK_PP(16'h11CDB,4);
TASK_PP(16'h11CDC,4);
TASK_PP(16'h11CDD,4);
TASK_PP(16'h11CDE,4);
TASK_PP(16'h11CDF,4);
TASK_PP(16'h11CE0,4);
TASK_PP(16'h11CE1,4);
TASK_PP(16'h11CE2,4);
TASK_PP(16'h11CE3,4);
TASK_PP(16'h11CE4,4);
TASK_PP(16'h11CE5,4);
TASK_PP(16'h11CE6,4);
TASK_PP(16'h11CE7,4);
TASK_PP(16'h11CE8,4);
TASK_PP(16'h11CE9,4);
TASK_PP(16'h11CEA,4);
TASK_PP(16'h11CEB,4);
TASK_PP(16'h11CEC,4);
TASK_PP(16'h11CED,4);
TASK_PP(16'h11CEE,4);
TASK_PP(16'h11CEF,4);
TASK_PP(16'h11CF0,4);
TASK_PP(16'h11CF1,4);
TASK_PP(16'h11CF2,4);
TASK_PP(16'h11CF3,4);
TASK_PP(16'h11CF4,4);
TASK_PP(16'h11CF5,4);
TASK_PP(16'h11CF6,4);
TASK_PP(16'h11CF7,4);
TASK_PP(16'h11CF8,4);
TASK_PP(16'h11CF9,4);
TASK_PP(16'h11CFA,4);
TASK_PP(16'h11CFB,4);
TASK_PP(16'h11CFC,4);
TASK_PP(16'h11CFD,4);
TASK_PP(16'h11CFE,4);
TASK_PP(16'h11CFF,4);
TASK_PP(16'h11D00,4);
TASK_PP(16'h11D01,4);
TASK_PP(16'h11D02,4);
TASK_PP(16'h11D03,4);
TASK_PP(16'h11D04,4);
TASK_PP(16'h11D05,4);
TASK_PP(16'h11D06,4);
TASK_PP(16'h11D07,4);
TASK_PP(16'h11D08,4);
TASK_PP(16'h11D09,4);
TASK_PP(16'h11D0A,4);
TASK_PP(16'h11D0B,4);
TASK_PP(16'h11D0C,4);
TASK_PP(16'h11D0D,4);
TASK_PP(16'h11D0E,4);
TASK_PP(16'h11D0F,4);
TASK_PP(16'h11D10,4);
TASK_PP(16'h11D11,4);
TASK_PP(16'h11D12,4);
TASK_PP(16'h11D13,4);
TASK_PP(16'h11D14,4);
TASK_PP(16'h11D15,4);
TASK_PP(16'h11D16,4);
TASK_PP(16'h11D17,4);
TASK_PP(16'h11D18,4);
TASK_PP(16'h11D19,4);
TASK_PP(16'h11D1A,4);
TASK_PP(16'h11D1B,4);
TASK_PP(16'h11D1C,4);
TASK_PP(16'h11D1D,4);
TASK_PP(16'h11D1E,4);
TASK_PP(16'h11D1F,4);
TASK_PP(16'h11D20,4);
TASK_PP(16'h11D21,4);
TASK_PP(16'h11D22,4);
TASK_PP(16'h11D23,4);
TASK_PP(16'h11D24,4);
TASK_PP(16'h11D25,4);
TASK_PP(16'h11D26,4);
TASK_PP(16'h11D27,4);
TASK_PP(16'h11D28,4);
TASK_PP(16'h11D29,4);
TASK_PP(16'h11D2A,4);
TASK_PP(16'h11D2B,4);
TASK_PP(16'h11D2C,4);
TASK_PP(16'h11D2D,4);
TASK_PP(16'h11D2E,4);
TASK_PP(16'h11D2F,4);
TASK_PP(16'h11D30,4);
TASK_PP(16'h11D31,4);
TASK_PP(16'h11D32,4);
TASK_PP(16'h11D33,4);
TASK_PP(16'h11D34,4);
TASK_PP(16'h11D35,4);
TASK_PP(16'h11D36,4);
TASK_PP(16'h11D37,4);
TASK_PP(16'h11D38,4);
TASK_PP(16'h11D39,4);
TASK_PP(16'h11D3A,4);
TASK_PP(16'h11D3B,4);
TASK_PP(16'h11D3C,4);
TASK_PP(16'h11D3D,4);
TASK_PP(16'h11D3E,4);
TASK_PP(16'h11D3F,4);
TASK_PP(16'h11D40,4);
TASK_PP(16'h11D41,4);
TASK_PP(16'h11D42,4);
TASK_PP(16'h11D43,4);
TASK_PP(16'h11D44,4);
TASK_PP(16'h11D45,4);
TASK_PP(16'h11D46,4);
TASK_PP(16'h11D47,4);
TASK_PP(16'h11D48,4);
TASK_PP(16'h11D49,4);
TASK_PP(16'h11D4A,4);
TASK_PP(16'h11D4B,4);
TASK_PP(16'h11D4C,4);
TASK_PP(16'h11D4D,4);
TASK_PP(16'h11D4E,4);
TASK_PP(16'h11D4F,4);
TASK_PP(16'h11D50,4);
TASK_PP(16'h11D51,4);
TASK_PP(16'h11D52,4);
TASK_PP(16'h11D53,4);
TASK_PP(16'h11D54,4);
TASK_PP(16'h11D55,4);
TASK_PP(16'h11D56,4);
TASK_PP(16'h11D57,4);
TASK_PP(16'h11D58,4);
TASK_PP(16'h11D59,4);
TASK_PP(16'h11D5A,4);
TASK_PP(16'h11D5B,4);
TASK_PP(16'h11D5C,4);
TASK_PP(16'h11D5D,4);
TASK_PP(16'h11D5E,4);
TASK_PP(16'h11D5F,4);
TASK_PP(16'h11D60,4);
TASK_PP(16'h11D61,4);
TASK_PP(16'h11D62,4);
TASK_PP(16'h11D63,4);
TASK_PP(16'h11D64,4);
TASK_PP(16'h11D65,4);
TASK_PP(16'h11D66,4);
TASK_PP(16'h11D67,4);
TASK_PP(16'h11D68,4);
TASK_PP(16'h11D69,4);
TASK_PP(16'h11D6A,4);
TASK_PP(16'h11D6B,4);
TASK_PP(16'h11D6C,4);
TASK_PP(16'h11D6D,4);
TASK_PP(16'h11D6E,4);
TASK_PP(16'h11D6F,4);
TASK_PP(16'h11D70,4);
TASK_PP(16'h11D71,4);
TASK_PP(16'h11D72,4);
TASK_PP(16'h11D73,4);
TASK_PP(16'h11D74,4);
TASK_PP(16'h11D75,4);
TASK_PP(16'h11D76,4);
TASK_PP(16'h11D77,4);
TASK_PP(16'h11D78,4);
TASK_PP(16'h11D79,4);
TASK_PP(16'h11D7A,4);
TASK_PP(16'h11D7B,4);
TASK_PP(16'h11D7C,4);
TASK_PP(16'h11D7D,4);
TASK_PP(16'h11D7E,4);
TASK_PP(16'h11D7F,4);
TASK_PP(16'h11D80,4);
TASK_PP(16'h11D81,4);
TASK_PP(16'h11D82,4);
TASK_PP(16'h11D83,4);
TASK_PP(16'h11D84,4);
TASK_PP(16'h11D85,4);
TASK_PP(16'h11D86,4);
TASK_PP(16'h11D87,4);
TASK_PP(16'h11D88,4);
TASK_PP(16'h11D89,4);
TASK_PP(16'h11D8A,4);
TASK_PP(16'h11D8B,4);
TASK_PP(16'h11D8C,4);
TASK_PP(16'h11D8D,4);
TASK_PP(16'h11D8E,4);
TASK_PP(16'h11D8F,4);
TASK_PP(16'h11D90,4);
TASK_PP(16'h11D91,4);
TASK_PP(16'h11D92,4);
TASK_PP(16'h11D93,4);
TASK_PP(16'h11D94,4);
TASK_PP(16'h11D95,4);
TASK_PP(16'h11D96,4);
TASK_PP(16'h11D97,4);
TASK_PP(16'h11D98,4);
TASK_PP(16'h11D99,4);
TASK_PP(16'h11D9A,4);
TASK_PP(16'h11D9B,4);
TASK_PP(16'h11D9C,4);
TASK_PP(16'h11D9D,4);
TASK_PP(16'h11D9E,4);
TASK_PP(16'h11D9F,4);
TASK_PP(16'h11DA0,4);
TASK_PP(16'h11DA1,4);
TASK_PP(16'h11DA2,4);
TASK_PP(16'h11DA3,4);
TASK_PP(16'h11DA4,4);
TASK_PP(16'h11DA5,4);
TASK_PP(16'h11DA6,4);
TASK_PP(16'h11DA7,4);
TASK_PP(16'h11DA8,4);
TASK_PP(16'h11DA9,4);
TASK_PP(16'h11DAA,4);
TASK_PP(16'h11DAB,4);
TASK_PP(16'h11DAC,4);
TASK_PP(16'h11DAD,4);
TASK_PP(16'h11DAE,4);
TASK_PP(16'h11DAF,4);
TASK_PP(16'h11DB0,4);
TASK_PP(16'h11DB1,4);
TASK_PP(16'h11DB2,4);
TASK_PP(16'h11DB3,4);
TASK_PP(16'h11DB4,4);
TASK_PP(16'h11DB5,4);
TASK_PP(16'h11DB6,4);
TASK_PP(16'h11DB7,4);
TASK_PP(16'h11DB8,4);
TASK_PP(16'h11DB9,4);
TASK_PP(16'h11DBA,4);
TASK_PP(16'h11DBB,4);
TASK_PP(16'h11DBC,4);
TASK_PP(16'h11DBD,4);
TASK_PP(16'h11DBE,4);
TASK_PP(16'h11DBF,4);
TASK_PP(16'h11DC0,4);
TASK_PP(16'h11DC1,4);
TASK_PP(16'h11DC2,4);
TASK_PP(16'h11DC3,4);
TASK_PP(16'h11DC4,4);
TASK_PP(16'h11DC5,4);
TASK_PP(16'h11DC6,4);
TASK_PP(16'h11DC7,4);
TASK_PP(16'h11DC8,4);
TASK_PP(16'h11DC9,4);
TASK_PP(16'h11DCA,4);
TASK_PP(16'h11DCB,4);
TASK_PP(16'h11DCC,4);
TASK_PP(16'h11DCD,4);
TASK_PP(16'h11DCE,4);
TASK_PP(16'h11DCF,4);
TASK_PP(16'h11DD0,4);
TASK_PP(16'h11DD1,4);
TASK_PP(16'h11DD2,4);
TASK_PP(16'h11DD3,4);
TASK_PP(16'h11DD4,4);
TASK_PP(16'h11DD5,4);
TASK_PP(16'h11DD6,4);
TASK_PP(16'h11DD7,4);
TASK_PP(16'h11DD8,4);
TASK_PP(16'h11DD9,4);
TASK_PP(16'h11DDA,4);
TASK_PP(16'h11DDB,4);
TASK_PP(16'h11DDC,4);
TASK_PP(16'h11DDD,4);
TASK_PP(16'h11DDE,4);
TASK_PP(16'h11DDF,4);
TASK_PP(16'h11DE0,4);
TASK_PP(16'h11DE1,4);
TASK_PP(16'h11DE2,4);
TASK_PP(16'h11DE3,4);
TASK_PP(16'h11DE4,4);
TASK_PP(16'h11DE5,4);
TASK_PP(16'h11DE6,4);
TASK_PP(16'h11DE7,4);
TASK_PP(16'h11DE8,4);
TASK_PP(16'h11DE9,4);
TASK_PP(16'h11DEA,4);
TASK_PP(16'h11DEB,4);
TASK_PP(16'h11DEC,4);
TASK_PP(16'h11DED,4);
TASK_PP(16'h11DEE,4);
TASK_PP(16'h11DEF,4);
TASK_PP(16'h11DF0,4);
TASK_PP(16'h11DF1,4);
TASK_PP(16'h11DF2,4);
TASK_PP(16'h11DF3,4);
TASK_PP(16'h11DF4,4);
TASK_PP(16'h11DF5,4);
TASK_PP(16'h11DF6,4);
TASK_PP(16'h11DF7,4);
TASK_PP(16'h11DF8,4);
TASK_PP(16'h11DF9,4);
TASK_PP(16'h11DFA,4);
TASK_PP(16'h11DFB,4);
TASK_PP(16'h11DFC,4);
TASK_PP(16'h11DFD,4);
TASK_PP(16'h11DFE,4);
TASK_PP(16'h11DFF,4);
TASK_PP(16'h11E00,4);
TASK_PP(16'h11E01,4);
TASK_PP(16'h11E02,4);
TASK_PP(16'h11E03,4);
TASK_PP(16'h11E04,4);
TASK_PP(16'h11E05,4);
TASK_PP(16'h11E06,4);
TASK_PP(16'h11E07,4);
TASK_PP(16'h11E08,4);
TASK_PP(16'h11E09,4);
TASK_PP(16'h11E0A,4);
TASK_PP(16'h11E0B,4);
TASK_PP(16'h11E0C,4);
TASK_PP(16'h11E0D,4);
TASK_PP(16'h11E0E,4);
TASK_PP(16'h11E0F,4);
TASK_PP(16'h11E10,4);
TASK_PP(16'h11E11,4);
TASK_PP(16'h11E12,4);
TASK_PP(16'h11E13,4);
TASK_PP(16'h11E14,4);
TASK_PP(16'h11E15,4);
TASK_PP(16'h11E16,4);
TASK_PP(16'h11E17,4);
TASK_PP(16'h11E18,4);
TASK_PP(16'h11E19,4);
TASK_PP(16'h11E1A,4);
TASK_PP(16'h11E1B,4);
TASK_PP(16'h11E1C,4);
TASK_PP(16'h11E1D,4);
TASK_PP(16'h11E1E,4);
TASK_PP(16'h11E1F,4);
TASK_PP(16'h11E20,4);
TASK_PP(16'h11E21,4);
TASK_PP(16'h11E22,4);
TASK_PP(16'h11E23,4);
TASK_PP(16'h11E24,4);
TASK_PP(16'h11E25,4);
TASK_PP(16'h11E26,4);
TASK_PP(16'h11E27,4);
TASK_PP(16'h11E28,4);
TASK_PP(16'h11E29,4);
TASK_PP(16'h11E2A,4);
TASK_PP(16'h11E2B,4);
TASK_PP(16'h11E2C,4);
TASK_PP(16'h11E2D,4);
TASK_PP(16'h11E2E,4);
TASK_PP(16'h11E2F,4);
TASK_PP(16'h11E30,4);
TASK_PP(16'h11E31,4);
TASK_PP(16'h11E32,4);
TASK_PP(16'h11E33,4);
TASK_PP(16'h11E34,4);
TASK_PP(16'h11E35,4);
TASK_PP(16'h11E36,4);
TASK_PP(16'h11E37,4);
TASK_PP(16'h11E38,4);
TASK_PP(16'h11E39,4);
TASK_PP(16'h11E3A,4);
TASK_PP(16'h11E3B,4);
TASK_PP(16'h11E3C,4);
TASK_PP(16'h11E3D,4);
TASK_PP(16'h11E3E,4);
TASK_PP(16'h11E3F,4);
TASK_PP(16'h11E40,4);
TASK_PP(16'h11E41,4);
TASK_PP(16'h11E42,4);
TASK_PP(16'h11E43,4);
TASK_PP(16'h11E44,4);
TASK_PP(16'h11E45,4);
TASK_PP(16'h11E46,4);
TASK_PP(16'h11E47,4);
TASK_PP(16'h11E48,4);
TASK_PP(16'h11E49,4);
TASK_PP(16'h11E4A,4);
TASK_PP(16'h11E4B,4);
TASK_PP(16'h11E4C,4);
TASK_PP(16'h11E4D,4);
TASK_PP(16'h11E4E,4);
TASK_PP(16'h11E4F,4);
TASK_PP(16'h11E50,4);
TASK_PP(16'h11E51,4);
TASK_PP(16'h11E52,4);
TASK_PP(16'h11E53,4);
TASK_PP(16'h11E54,4);
TASK_PP(16'h11E55,4);
TASK_PP(16'h11E56,4);
TASK_PP(16'h11E57,4);
TASK_PP(16'h11E58,4);
TASK_PP(16'h11E59,4);
TASK_PP(16'h11E5A,4);
TASK_PP(16'h11E5B,4);
TASK_PP(16'h11E5C,4);
TASK_PP(16'h11E5D,4);
TASK_PP(16'h11E5E,4);
TASK_PP(16'h11E5F,4);
TASK_PP(16'h11E60,4);
TASK_PP(16'h11E61,4);
TASK_PP(16'h11E62,4);
TASK_PP(16'h11E63,4);
TASK_PP(16'h11E64,4);
TASK_PP(16'h11E65,4);
TASK_PP(16'h11E66,4);
TASK_PP(16'h11E67,4);
TASK_PP(16'h11E68,4);
TASK_PP(16'h11E69,4);
TASK_PP(16'h11E6A,4);
TASK_PP(16'h11E6B,4);
TASK_PP(16'h11E6C,4);
TASK_PP(16'h11E6D,4);
TASK_PP(16'h11E6E,4);
TASK_PP(16'h11E6F,4);
TASK_PP(16'h11E70,4);
TASK_PP(16'h11E71,4);
TASK_PP(16'h11E72,4);
TASK_PP(16'h11E73,4);
TASK_PP(16'h11E74,4);
TASK_PP(16'h11E75,4);
TASK_PP(16'h11E76,4);
TASK_PP(16'h11E77,4);
TASK_PP(16'h11E78,4);
TASK_PP(16'h11E79,4);
TASK_PP(16'h11E7A,4);
TASK_PP(16'h11E7B,4);
TASK_PP(16'h11E7C,4);
TASK_PP(16'h11E7D,4);
TASK_PP(16'h11E7E,4);
TASK_PP(16'h11E7F,4);
TASK_PP(16'h11E80,4);
TASK_PP(16'h11E81,4);
TASK_PP(16'h11E82,4);
TASK_PP(16'h11E83,4);
TASK_PP(16'h11E84,4);
TASK_PP(16'h11E85,4);
TASK_PP(16'h11E86,4);
TASK_PP(16'h11E87,4);
TASK_PP(16'h11E88,4);
TASK_PP(16'h11E89,4);
TASK_PP(16'h11E8A,4);
TASK_PP(16'h11E8B,4);
TASK_PP(16'h11E8C,4);
TASK_PP(16'h11E8D,4);
TASK_PP(16'h11E8E,4);
TASK_PP(16'h11E8F,4);
TASK_PP(16'h11E90,4);
TASK_PP(16'h11E91,4);
TASK_PP(16'h11E92,4);
TASK_PP(16'h11E93,4);
TASK_PP(16'h11E94,4);
TASK_PP(16'h11E95,4);
TASK_PP(16'h11E96,4);
TASK_PP(16'h11E97,4);
TASK_PP(16'h11E98,4);
TASK_PP(16'h11E99,4);
TASK_PP(16'h11E9A,4);
TASK_PP(16'h11E9B,4);
TASK_PP(16'h11E9C,4);
TASK_PP(16'h11E9D,4);
TASK_PP(16'h11E9E,4);
TASK_PP(16'h11E9F,4);
TASK_PP(16'h11EA0,4);
TASK_PP(16'h11EA1,4);
TASK_PP(16'h11EA2,4);
TASK_PP(16'h11EA3,4);
TASK_PP(16'h11EA4,4);
TASK_PP(16'h11EA5,4);
TASK_PP(16'h11EA6,4);
TASK_PP(16'h11EA7,4);
TASK_PP(16'h11EA8,4);
TASK_PP(16'h11EA9,4);
TASK_PP(16'h11EAA,4);
TASK_PP(16'h11EAB,4);
TASK_PP(16'h11EAC,4);
TASK_PP(16'h11EAD,4);
TASK_PP(16'h11EAE,4);
TASK_PP(16'h11EAF,4);
TASK_PP(16'h11EB0,4);
TASK_PP(16'h11EB1,4);
TASK_PP(16'h11EB2,4);
TASK_PP(16'h11EB3,4);
TASK_PP(16'h11EB4,4);
TASK_PP(16'h11EB5,4);
TASK_PP(16'h11EB6,4);
TASK_PP(16'h11EB7,4);
TASK_PP(16'h11EB8,4);
TASK_PP(16'h11EB9,4);
TASK_PP(16'h11EBA,4);
TASK_PP(16'h11EBB,4);
TASK_PP(16'h11EBC,4);
TASK_PP(16'h11EBD,4);
TASK_PP(16'h11EBE,4);
TASK_PP(16'h11EBF,4);
TASK_PP(16'h11EC0,4);
TASK_PP(16'h11EC1,4);
TASK_PP(16'h11EC2,4);
TASK_PP(16'h11EC3,4);
TASK_PP(16'h11EC4,4);
TASK_PP(16'h11EC5,4);
TASK_PP(16'h11EC6,4);
TASK_PP(16'h11EC7,4);
TASK_PP(16'h11EC8,4);
TASK_PP(16'h11EC9,4);
TASK_PP(16'h11ECA,4);
TASK_PP(16'h11ECB,4);
TASK_PP(16'h11ECC,4);
TASK_PP(16'h11ECD,4);
TASK_PP(16'h11ECE,4);
TASK_PP(16'h11ECF,4);
TASK_PP(16'h11ED0,4);
TASK_PP(16'h11ED1,4);
TASK_PP(16'h11ED2,4);
TASK_PP(16'h11ED3,4);
TASK_PP(16'h11ED4,4);
TASK_PP(16'h11ED5,4);
TASK_PP(16'h11ED6,4);
TASK_PP(16'h11ED7,4);
TASK_PP(16'h11ED8,4);
TASK_PP(16'h11ED9,4);
TASK_PP(16'h11EDA,4);
TASK_PP(16'h11EDB,4);
TASK_PP(16'h11EDC,4);
TASK_PP(16'h11EDD,4);
TASK_PP(16'h11EDE,4);
TASK_PP(16'h11EDF,4);
TASK_PP(16'h11EE0,4);
TASK_PP(16'h11EE1,4);
TASK_PP(16'h11EE2,4);
TASK_PP(16'h11EE3,4);
TASK_PP(16'h11EE4,4);
TASK_PP(16'h11EE5,4);
TASK_PP(16'h11EE6,4);
TASK_PP(16'h11EE7,4);
TASK_PP(16'h11EE8,4);
TASK_PP(16'h11EE9,4);
TASK_PP(16'h11EEA,4);
TASK_PP(16'h11EEB,4);
TASK_PP(16'h11EEC,4);
TASK_PP(16'h11EED,4);
TASK_PP(16'h11EEE,4);
TASK_PP(16'h11EEF,4);
TASK_PP(16'h11EF0,4);
TASK_PP(16'h11EF1,4);
TASK_PP(16'h11EF2,4);
TASK_PP(16'h11EF3,4);
TASK_PP(16'h11EF4,4);
TASK_PP(16'h11EF5,4);
TASK_PP(16'h11EF6,4);
TASK_PP(16'h11EF7,4);
TASK_PP(16'h11EF8,4);
TASK_PP(16'h11EF9,4);
TASK_PP(16'h11EFA,4);
TASK_PP(16'h11EFB,4);
TASK_PP(16'h11EFC,4);
TASK_PP(16'h11EFD,4);
TASK_PP(16'h11EFE,4);
TASK_PP(16'h11EFF,4);
TASK_PP(16'h11F00,4);
TASK_PP(16'h11F01,4);
TASK_PP(16'h11F02,4);
TASK_PP(16'h11F03,4);
TASK_PP(16'h11F04,4);
TASK_PP(16'h11F05,4);
TASK_PP(16'h11F06,4);
TASK_PP(16'h11F07,4);
TASK_PP(16'h11F08,4);
TASK_PP(16'h11F09,4);
TASK_PP(16'h11F0A,4);
TASK_PP(16'h11F0B,4);
TASK_PP(16'h11F0C,4);
TASK_PP(16'h11F0D,4);
TASK_PP(16'h11F0E,4);
TASK_PP(16'h11F0F,4);
TASK_PP(16'h11F10,4);
TASK_PP(16'h11F11,4);
TASK_PP(16'h11F12,4);
TASK_PP(16'h11F13,4);
TASK_PP(16'h11F14,4);
TASK_PP(16'h11F15,4);
TASK_PP(16'h11F16,4);
TASK_PP(16'h11F17,4);
TASK_PP(16'h11F18,4);
TASK_PP(16'h11F19,4);
TASK_PP(16'h11F1A,4);
TASK_PP(16'h11F1B,4);
TASK_PP(16'h11F1C,4);
TASK_PP(16'h11F1D,4);
TASK_PP(16'h11F1E,4);
TASK_PP(16'h11F1F,4);
TASK_PP(16'h11F20,4);
TASK_PP(16'h11F21,4);
TASK_PP(16'h11F22,4);
TASK_PP(16'h11F23,4);
TASK_PP(16'h11F24,4);
TASK_PP(16'h11F25,4);
TASK_PP(16'h11F26,4);
TASK_PP(16'h11F27,4);
TASK_PP(16'h11F28,4);
TASK_PP(16'h11F29,4);
TASK_PP(16'h11F2A,4);
TASK_PP(16'h11F2B,4);
TASK_PP(16'h11F2C,4);
TASK_PP(16'h11F2D,4);
TASK_PP(16'h11F2E,4);
TASK_PP(16'h11F2F,4);
TASK_PP(16'h11F30,4);
TASK_PP(16'h11F31,4);
TASK_PP(16'h11F32,4);
TASK_PP(16'h11F33,4);
TASK_PP(16'h11F34,4);
TASK_PP(16'h11F35,4);
TASK_PP(16'h11F36,4);
TASK_PP(16'h11F37,4);
TASK_PP(16'h11F38,4);
TASK_PP(16'h11F39,4);
TASK_PP(16'h11F3A,4);
TASK_PP(16'h11F3B,4);
TASK_PP(16'h11F3C,4);
TASK_PP(16'h11F3D,4);
TASK_PP(16'h11F3E,4);
TASK_PP(16'h11F3F,4);
TASK_PP(16'h11F40,4);
TASK_PP(16'h11F41,4);
TASK_PP(16'h11F42,4);
TASK_PP(16'h11F43,4);
TASK_PP(16'h11F44,4);
TASK_PP(16'h11F45,4);
TASK_PP(16'h11F46,4);
TASK_PP(16'h11F47,4);
TASK_PP(16'h11F48,4);
TASK_PP(16'h11F49,4);
TASK_PP(16'h11F4A,4);
TASK_PP(16'h11F4B,4);
TASK_PP(16'h11F4C,4);
TASK_PP(16'h11F4D,4);
TASK_PP(16'h11F4E,4);
TASK_PP(16'h11F4F,4);
TASK_PP(16'h11F50,4);
TASK_PP(16'h11F51,4);
TASK_PP(16'h11F52,4);
TASK_PP(16'h11F53,4);
TASK_PP(16'h11F54,4);
TASK_PP(16'h11F55,4);
TASK_PP(16'h11F56,4);
TASK_PP(16'h11F57,4);
TASK_PP(16'h11F58,4);
TASK_PP(16'h11F59,4);
TASK_PP(16'h11F5A,4);
TASK_PP(16'h11F5B,4);
TASK_PP(16'h11F5C,4);
TASK_PP(16'h11F5D,4);
TASK_PP(16'h11F5E,4);
TASK_PP(16'h11F5F,4);
TASK_PP(16'h11F60,4);
TASK_PP(16'h11F61,4);
TASK_PP(16'h11F62,4);
TASK_PP(16'h11F63,4);
TASK_PP(16'h11F64,4);
TASK_PP(16'h11F65,4);
TASK_PP(16'h11F66,4);
TASK_PP(16'h11F67,4);
TASK_PP(16'h11F68,4);
TASK_PP(16'h11F69,4);
TASK_PP(16'h11F6A,4);
TASK_PP(16'h11F6B,4);
TASK_PP(16'h11F6C,4);
TASK_PP(16'h11F6D,4);
TASK_PP(16'h11F6E,4);
TASK_PP(16'h11F6F,4);
TASK_PP(16'h11F70,4);
TASK_PP(16'h11F71,4);
TASK_PP(16'h11F72,4);
TASK_PP(16'h11F73,4);
TASK_PP(16'h11F74,4);
TASK_PP(16'h11F75,4);
TASK_PP(16'h11F76,4);
TASK_PP(16'h11F77,4);
TASK_PP(16'h11F78,4);
TASK_PP(16'h11F79,4);
TASK_PP(16'h11F7A,4);
TASK_PP(16'h11F7B,4);
TASK_PP(16'h11F7C,4);
TASK_PP(16'h11F7D,4);
TASK_PP(16'h11F7E,4);
TASK_PP(16'h11F7F,4);
TASK_PP(16'h11F80,4);
TASK_PP(16'h11F81,4);
TASK_PP(16'h11F82,4);
TASK_PP(16'h11F83,4);
TASK_PP(16'h11F84,4);
TASK_PP(16'h11F85,4);
TASK_PP(16'h11F86,4);
TASK_PP(16'h11F87,4);
TASK_PP(16'h11F88,4);
TASK_PP(16'h11F89,4);
TASK_PP(16'h11F8A,4);
TASK_PP(16'h11F8B,4);
TASK_PP(16'h11F8C,4);
TASK_PP(16'h11F8D,4);
TASK_PP(16'h11F8E,4);
TASK_PP(16'h11F8F,4);
TASK_PP(16'h11F90,4);
TASK_PP(16'h11F91,4);
TASK_PP(16'h11F92,4);
TASK_PP(16'h11F93,4);
TASK_PP(16'h11F94,4);
TASK_PP(16'h11F95,4);
TASK_PP(16'h11F96,4);
TASK_PP(16'h11F97,4);
TASK_PP(16'h11F98,4);
TASK_PP(16'h11F99,4);
TASK_PP(16'h11F9A,4);
TASK_PP(16'h11F9B,4);
TASK_PP(16'h11F9C,4);
TASK_PP(16'h11F9D,4);
TASK_PP(16'h11F9E,4);
TASK_PP(16'h11F9F,4);
TASK_PP(16'h11FA0,4);
TASK_PP(16'h11FA1,4);
TASK_PP(16'h11FA2,4);
TASK_PP(16'h11FA3,4);
TASK_PP(16'h11FA4,4);
TASK_PP(16'h11FA5,4);
TASK_PP(16'h11FA6,4);
TASK_PP(16'h11FA7,4);
TASK_PP(16'h11FA8,4);
TASK_PP(16'h11FA9,4);
TASK_PP(16'h11FAA,4);
TASK_PP(16'h11FAB,4);
TASK_PP(16'h11FAC,4);
TASK_PP(16'h11FAD,4);
TASK_PP(16'h11FAE,4);
TASK_PP(16'h11FAF,4);
TASK_PP(16'h11FB0,4);
TASK_PP(16'h11FB1,4);
TASK_PP(16'h11FB2,4);
TASK_PP(16'h11FB3,4);
TASK_PP(16'h11FB4,4);
TASK_PP(16'h11FB5,4);
TASK_PP(16'h11FB6,4);
TASK_PP(16'h11FB7,4);
TASK_PP(16'h11FB8,4);
TASK_PP(16'h11FB9,4);
TASK_PP(16'h11FBA,4);
TASK_PP(16'h11FBB,4);
TASK_PP(16'h11FBC,4);
TASK_PP(16'h11FBD,4);
TASK_PP(16'h11FBE,4);
TASK_PP(16'h11FBF,4);
TASK_PP(16'h11FC0,4);
TASK_PP(16'h11FC1,4);
TASK_PP(16'h11FC2,4);
TASK_PP(16'h11FC3,4);
TASK_PP(16'h11FC4,4);
TASK_PP(16'h11FC5,4);
TASK_PP(16'h11FC6,4);
TASK_PP(16'h11FC7,4);
TASK_PP(16'h11FC8,4);
TASK_PP(16'h11FC9,4);
TASK_PP(16'h11FCA,4);
TASK_PP(16'h11FCB,4);
TASK_PP(16'h11FCC,4);
TASK_PP(16'h11FCD,4);
TASK_PP(16'h11FCE,4);
TASK_PP(16'h11FCF,4);
TASK_PP(16'h11FD0,4);
TASK_PP(16'h11FD1,4);
TASK_PP(16'h11FD2,4);
TASK_PP(16'h11FD3,4);
TASK_PP(16'h11FD4,4);
TASK_PP(16'h11FD5,4);
TASK_PP(16'h11FD6,4);
TASK_PP(16'h11FD7,4);
TASK_PP(16'h11FD8,4);
TASK_PP(16'h11FD9,4);
TASK_PP(16'h11FDA,4);
TASK_PP(16'h11FDB,4);
TASK_PP(16'h11FDC,4);
TASK_PP(16'h11FDD,4);
TASK_PP(16'h11FDE,4);
TASK_PP(16'h11FDF,4);
TASK_PP(16'h11FE0,4);
TASK_PP(16'h11FE1,4);
TASK_PP(16'h11FE2,4);
TASK_PP(16'h11FE3,4);
TASK_PP(16'h11FE4,4);
TASK_PP(16'h11FE5,4);
TASK_PP(16'h11FE6,4);
TASK_PP(16'h11FE7,4);
TASK_PP(16'h11FE8,4);
TASK_PP(16'h11FE9,4);
TASK_PP(16'h11FEA,4);
TASK_PP(16'h11FEB,4);
TASK_PP(16'h11FEC,4);
TASK_PP(16'h11FED,4);
TASK_PP(16'h11FEE,4);
TASK_PP(16'h11FEF,4);
TASK_PP(16'h11FF0,4);
TASK_PP(16'h11FF1,4);
TASK_PP(16'h11FF2,4);
TASK_PP(16'h11FF3,4);
TASK_PP(16'h11FF4,4);
TASK_PP(16'h11FF5,4);
TASK_PP(16'h11FF6,4);
TASK_PP(16'h11FF7,4);
TASK_PP(16'h11FF8,4);
TASK_PP(16'h11FF9,4);
TASK_PP(16'h11FFA,4);
TASK_PP(16'h11FFB,4);
TASK_PP(16'h11FFC,4);
TASK_PP(16'h11FFD,4);
TASK_PP(16'h11FFE,4);
TASK_PP(16'h11FFF,4);
TASK_PP(16'h12000,4);
TASK_PP(16'h12001,4);
TASK_PP(16'h12002,4);
TASK_PP(16'h12003,4);
TASK_PP(16'h12004,4);
TASK_PP(16'h12005,4);
TASK_PP(16'h12006,4);
TASK_PP(16'h12007,4);
TASK_PP(16'h12008,4);
TASK_PP(16'h12009,4);
TASK_PP(16'h1200A,4);
TASK_PP(16'h1200B,4);
TASK_PP(16'h1200C,4);
TASK_PP(16'h1200D,4);
TASK_PP(16'h1200E,4);
TASK_PP(16'h1200F,4);
TASK_PP(16'h12010,4);
TASK_PP(16'h12011,4);
TASK_PP(16'h12012,4);
TASK_PP(16'h12013,4);
TASK_PP(16'h12014,4);
TASK_PP(16'h12015,4);
TASK_PP(16'h12016,4);
TASK_PP(16'h12017,4);
TASK_PP(16'h12018,4);
TASK_PP(16'h12019,4);
TASK_PP(16'h1201A,4);
TASK_PP(16'h1201B,4);
TASK_PP(16'h1201C,4);
TASK_PP(16'h1201D,4);
TASK_PP(16'h1201E,4);
TASK_PP(16'h1201F,4);
TASK_PP(16'h12020,4);
TASK_PP(16'h12021,4);
TASK_PP(16'h12022,4);
TASK_PP(16'h12023,4);
TASK_PP(16'h12024,4);
TASK_PP(16'h12025,4);
TASK_PP(16'h12026,4);
TASK_PP(16'h12027,4);
TASK_PP(16'h12028,4);
TASK_PP(16'h12029,4);
TASK_PP(16'h1202A,4);
TASK_PP(16'h1202B,4);
TASK_PP(16'h1202C,4);
TASK_PP(16'h1202D,4);
TASK_PP(16'h1202E,4);
TASK_PP(16'h1202F,4);
TASK_PP(16'h12030,4);
TASK_PP(16'h12031,4);
TASK_PP(16'h12032,4);
TASK_PP(16'h12033,4);
TASK_PP(16'h12034,4);
TASK_PP(16'h12035,4);
TASK_PP(16'h12036,4);
TASK_PP(16'h12037,4);
TASK_PP(16'h12038,4);
TASK_PP(16'h12039,4);
TASK_PP(16'h1203A,4);
TASK_PP(16'h1203B,4);
TASK_PP(16'h1203C,4);
TASK_PP(16'h1203D,4);
TASK_PP(16'h1203E,4);
TASK_PP(16'h1203F,4);
TASK_PP(16'h12040,4);
TASK_PP(16'h12041,4);
TASK_PP(16'h12042,4);
TASK_PP(16'h12043,4);
TASK_PP(16'h12044,4);
TASK_PP(16'h12045,4);
TASK_PP(16'h12046,4);
TASK_PP(16'h12047,4);
TASK_PP(16'h12048,4);
TASK_PP(16'h12049,4);
TASK_PP(16'h1204A,4);
TASK_PP(16'h1204B,4);
TASK_PP(16'h1204C,4);
TASK_PP(16'h1204D,4);
TASK_PP(16'h1204E,4);
TASK_PP(16'h1204F,4);
TASK_PP(16'h12050,4);
TASK_PP(16'h12051,4);
TASK_PP(16'h12052,4);
TASK_PP(16'h12053,4);
TASK_PP(16'h12054,4);
TASK_PP(16'h12055,4);
TASK_PP(16'h12056,4);
TASK_PP(16'h12057,4);
TASK_PP(16'h12058,4);
TASK_PP(16'h12059,4);
TASK_PP(16'h1205A,4);
TASK_PP(16'h1205B,4);
TASK_PP(16'h1205C,4);
TASK_PP(16'h1205D,4);
TASK_PP(16'h1205E,4);
TASK_PP(16'h1205F,4);
TASK_PP(16'h12060,4);
TASK_PP(16'h12061,4);
TASK_PP(16'h12062,4);
TASK_PP(16'h12063,4);
TASK_PP(16'h12064,4);
TASK_PP(16'h12065,4);
TASK_PP(16'h12066,4);
TASK_PP(16'h12067,4);
TASK_PP(16'h12068,4);
TASK_PP(16'h12069,4);
TASK_PP(16'h1206A,4);
TASK_PP(16'h1206B,4);
TASK_PP(16'h1206C,4);
TASK_PP(16'h1206D,4);
TASK_PP(16'h1206E,4);
TASK_PP(16'h1206F,4);
TASK_PP(16'h12070,4);
TASK_PP(16'h12071,4);
TASK_PP(16'h12072,4);
TASK_PP(16'h12073,4);
TASK_PP(16'h12074,4);
TASK_PP(16'h12075,4);
TASK_PP(16'h12076,4);
TASK_PP(16'h12077,4);
TASK_PP(16'h12078,4);
TASK_PP(16'h12079,4);
TASK_PP(16'h1207A,4);
TASK_PP(16'h1207B,4);
TASK_PP(16'h1207C,4);
TASK_PP(16'h1207D,4);
TASK_PP(16'h1207E,4);
TASK_PP(16'h1207F,4);
TASK_PP(16'h12080,4);
TASK_PP(16'h12081,4);
TASK_PP(16'h12082,4);
TASK_PP(16'h12083,4);
TASK_PP(16'h12084,4);
TASK_PP(16'h12085,4);
TASK_PP(16'h12086,4);
TASK_PP(16'h12087,4);
TASK_PP(16'h12088,4);
TASK_PP(16'h12089,4);
TASK_PP(16'h1208A,4);
TASK_PP(16'h1208B,4);
TASK_PP(16'h1208C,4);
TASK_PP(16'h1208D,4);
TASK_PP(16'h1208E,4);
TASK_PP(16'h1208F,4);
TASK_PP(16'h12090,4);
TASK_PP(16'h12091,4);
TASK_PP(16'h12092,4);
TASK_PP(16'h12093,4);
TASK_PP(16'h12094,4);
TASK_PP(16'h12095,4);
TASK_PP(16'h12096,4);
TASK_PP(16'h12097,4);
TASK_PP(16'h12098,4);
TASK_PP(16'h12099,4);
TASK_PP(16'h1209A,4);
TASK_PP(16'h1209B,4);
TASK_PP(16'h1209C,4);
TASK_PP(16'h1209D,4);
TASK_PP(16'h1209E,4);
TASK_PP(16'h1209F,4);
TASK_PP(16'h120A0,4);
TASK_PP(16'h120A1,4);
TASK_PP(16'h120A2,4);
TASK_PP(16'h120A3,4);
TASK_PP(16'h120A4,4);
TASK_PP(16'h120A5,4);
TASK_PP(16'h120A6,4);
TASK_PP(16'h120A7,4);
TASK_PP(16'h120A8,4);
TASK_PP(16'h120A9,4);
TASK_PP(16'h120AA,4);
TASK_PP(16'h120AB,4);
TASK_PP(16'h120AC,4);
TASK_PP(16'h120AD,4);
TASK_PP(16'h120AE,4);
TASK_PP(16'h120AF,4);
TASK_PP(16'h120B0,4);
TASK_PP(16'h120B1,4);
TASK_PP(16'h120B2,4);
TASK_PP(16'h120B3,4);
TASK_PP(16'h120B4,4);
TASK_PP(16'h120B5,4);
TASK_PP(16'h120B6,4);
TASK_PP(16'h120B7,4);
TASK_PP(16'h120B8,4);
TASK_PP(16'h120B9,4);
TASK_PP(16'h120BA,4);
TASK_PP(16'h120BB,4);
TASK_PP(16'h120BC,4);
TASK_PP(16'h120BD,4);
TASK_PP(16'h120BE,4);
TASK_PP(16'h120BF,4);
TASK_PP(16'h120C0,4);
TASK_PP(16'h120C1,4);
TASK_PP(16'h120C2,4);
TASK_PP(16'h120C3,4);
TASK_PP(16'h120C4,4);
TASK_PP(16'h120C5,4);
TASK_PP(16'h120C6,4);
TASK_PP(16'h120C7,4);
TASK_PP(16'h120C8,4);
TASK_PP(16'h120C9,4);
TASK_PP(16'h120CA,4);
TASK_PP(16'h120CB,4);
TASK_PP(16'h120CC,4);
TASK_PP(16'h120CD,4);
TASK_PP(16'h120CE,4);
TASK_PP(16'h120CF,4);
TASK_PP(16'h120D0,4);
TASK_PP(16'h120D1,4);
TASK_PP(16'h120D2,4);
TASK_PP(16'h120D3,4);
TASK_PP(16'h120D4,4);
TASK_PP(16'h120D5,4);
TASK_PP(16'h120D6,4);
TASK_PP(16'h120D7,4);
TASK_PP(16'h120D8,4);
TASK_PP(16'h120D9,4);
TASK_PP(16'h120DA,4);
TASK_PP(16'h120DB,4);
TASK_PP(16'h120DC,4);
TASK_PP(16'h120DD,4);
TASK_PP(16'h120DE,4);
TASK_PP(16'h120DF,4);
TASK_PP(16'h120E0,4);
TASK_PP(16'h120E1,4);
TASK_PP(16'h120E2,4);
TASK_PP(16'h120E3,4);
TASK_PP(16'h120E4,4);
TASK_PP(16'h120E5,4);
TASK_PP(16'h120E6,4);
TASK_PP(16'h120E7,4);
TASK_PP(16'h120E8,4);
TASK_PP(16'h120E9,4);
TASK_PP(16'h120EA,4);
TASK_PP(16'h120EB,4);
TASK_PP(16'h120EC,4);
TASK_PP(16'h120ED,4);
TASK_PP(16'h120EE,4);
TASK_PP(16'h120EF,4);
TASK_PP(16'h120F0,4);
TASK_PP(16'h120F1,4);
TASK_PP(16'h120F2,4);
TASK_PP(16'h120F3,4);
TASK_PP(16'h120F4,4);
TASK_PP(16'h120F5,4);
TASK_PP(16'h120F6,4);
TASK_PP(16'h120F7,4);
TASK_PP(16'h120F8,4);
TASK_PP(16'h120F9,4);
TASK_PP(16'h120FA,4);
TASK_PP(16'h120FB,4);
TASK_PP(16'h120FC,4);
TASK_PP(16'h120FD,4);
TASK_PP(16'h120FE,4);
TASK_PP(16'h120FF,4);
TASK_PP(16'h12100,4);
TASK_PP(16'h12101,4);
TASK_PP(16'h12102,4);
TASK_PP(16'h12103,4);
TASK_PP(16'h12104,4);
TASK_PP(16'h12105,4);
TASK_PP(16'h12106,4);
TASK_PP(16'h12107,4);
TASK_PP(16'h12108,4);
TASK_PP(16'h12109,4);
TASK_PP(16'h1210A,4);
TASK_PP(16'h1210B,4);
TASK_PP(16'h1210C,4);
TASK_PP(16'h1210D,4);
TASK_PP(16'h1210E,4);
TASK_PP(16'h1210F,4);
TASK_PP(16'h12110,4);
TASK_PP(16'h12111,4);
TASK_PP(16'h12112,4);
TASK_PP(16'h12113,4);
TASK_PP(16'h12114,4);
TASK_PP(16'h12115,4);
TASK_PP(16'h12116,4);
TASK_PP(16'h12117,4);
TASK_PP(16'h12118,4);
TASK_PP(16'h12119,4);
TASK_PP(16'h1211A,4);
TASK_PP(16'h1211B,4);
TASK_PP(16'h1211C,4);
TASK_PP(16'h1211D,4);
TASK_PP(16'h1211E,4);
TASK_PP(16'h1211F,4);
TASK_PP(16'h12120,4);
TASK_PP(16'h12121,4);
TASK_PP(16'h12122,4);
TASK_PP(16'h12123,4);
TASK_PP(16'h12124,4);
TASK_PP(16'h12125,4);
TASK_PP(16'h12126,4);
TASK_PP(16'h12127,4);
TASK_PP(16'h12128,4);
TASK_PP(16'h12129,4);
TASK_PP(16'h1212A,4);
TASK_PP(16'h1212B,4);
TASK_PP(16'h1212C,4);
TASK_PP(16'h1212D,4);
TASK_PP(16'h1212E,4);
TASK_PP(16'h1212F,4);
TASK_PP(16'h12130,4);
TASK_PP(16'h12131,4);
TASK_PP(16'h12132,4);
TASK_PP(16'h12133,4);
TASK_PP(16'h12134,4);
TASK_PP(16'h12135,4);
TASK_PP(16'h12136,4);
TASK_PP(16'h12137,4);
TASK_PP(16'h12138,4);
TASK_PP(16'h12139,4);
TASK_PP(16'h1213A,4);
TASK_PP(16'h1213B,4);
TASK_PP(16'h1213C,4);
TASK_PP(16'h1213D,4);
TASK_PP(16'h1213E,4);
TASK_PP(16'h1213F,4);
TASK_PP(16'h12140,4);
TASK_PP(16'h12141,4);
TASK_PP(16'h12142,4);
TASK_PP(16'h12143,4);
TASK_PP(16'h12144,4);
TASK_PP(16'h12145,4);
TASK_PP(16'h12146,4);
TASK_PP(16'h12147,4);
TASK_PP(16'h12148,4);
TASK_PP(16'h12149,4);
TASK_PP(16'h1214A,4);
TASK_PP(16'h1214B,4);
TASK_PP(16'h1214C,4);
TASK_PP(16'h1214D,4);
TASK_PP(16'h1214E,4);
TASK_PP(16'h1214F,4);
TASK_PP(16'h12150,4);
TASK_PP(16'h12151,4);
TASK_PP(16'h12152,4);
TASK_PP(16'h12153,4);
TASK_PP(16'h12154,4);
TASK_PP(16'h12155,4);
TASK_PP(16'h12156,4);
TASK_PP(16'h12157,4);
TASK_PP(16'h12158,4);
TASK_PP(16'h12159,4);
TASK_PP(16'h1215A,4);
TASK_PP(16'h1215B,4);
TASK_PP(16'h1215C,4);
TASK_PP(16'h1215D,4);
TASK_PP(16'h1215E,4);
TASK_PP(16'h1215F,4);
TASK_PP(16'h12160,4);
TASK_PP(16'h12161,4);
TASK_PP(16'h12162,4);
TASK_PP(16'h12163,4);
TASK_PP(16'h12164,4);
TASK_PP(16'h12165,4);
TASK_PP(16'h12166,4);
TASK_PP(16'h12167,4);
TASK_PP(16'h12168,4);
TASK_PP(16'h12169,4);
TASK_PP(16'h1216A,4);
TASK_PP(16'h1216B,4);
TASK_PP(16'h1216C,4);
TASK_PP(16'h1216D,4);
TASK_PP(16'h1216E,4);
TASK_PP(16'h1216F,4);
TASK_PP(16'h12170,4);
TASK_PP(16'h12171,4);
TASK_PP(16'h12172,4);
TASK_PP(16'h12173,4);
TASK_PP(16'h12174,4);
TASK_PP(16'h12175,4);
TASK_PP(16'h12176,4);
TASK_PP(16'h12177,4);
TASK_PP(16'h12178,4);
TASK_PP(16'h12179,4);
TASK_PP(16'h1217A,4);
TASK_PP(16'h1217B,4);
TASK_PP(16'h1217C,4);
TASK_PP(16'h1217D,4);
TASK_PP(16'h1217E,4);
TASK_PP(16'h1217F,4);
TASK_PP(16'h12180,4);
TASK_PP(16'h12181,4);
TASK_PP(16'h12182,4);
TASK_PP(16'h12183,4);
TASK_PP(16'h12184,4);
TASK_PP(16'h12185,4);
TASK_PP(16'h12186,4);
TASK_PP(16'h12187,4);
TASK_PP(16'h12188,4);
TASK_PP(16'h12189,4);
TASK_PP(16'h1218A,4);
TASK_PP(16'h1218B,4);
TASK_PP(16'h1218C,4);
TASK_PP(16'h1218D,4);
TASK_PP(16'h1218E,4);
TASK_PP(16'h1218F,4);
TASK_PP(16'h12190,4);
TASK_PP(16'h12191,4);
TASK_PP(16'h12192,4);
TASK_PP(16'h12193,4);
TASK_PP(16'h12194,4);
TASK_PP(16'h12195,4);
TASK_PP(16'h12196,4);
TASK_PP(16'h12197,4);
TASK_PP(16'h12198,4);
TASK_PP(16'h12199,4);
TASK_PP(16'h1219A,4);
TASK_PP(16'h1219B,4);
TASK_PP(16'h1219C,4);
TASK_PP(16'h1219D,4);
TASK_PP(16'h1219E,4);
TASK_PP(16'h1219F,4);
TASK_PP(16'h121A0,4);
TASK_PP(16'h121A1,4);
TASK_PP(16'h121A2,4);
TASK_PP(16'h121A3,4);
TASK_PP(16'h121A4,4);
TASK_PP(16'h121A5,4);
TASK_PP(16'h121A6,4);
TASK_PP(16'h121A7,4);
TASK_PP(16'h121A8,4);
TASK_PP(16'h121A9,4);
TASK_PP(16'h121AA,4);
TASK_PP(16'h121AB,4);
TASK_PP(16'h121AC,4);
TASK_PP(16'h121AD,4);
TASK_PP(16'h121AE,4);
TASK_PP(16'h121AF,4);
TASK_PP(16'h121B0,4);
TASK_PP(16'h121B1,4);
TASK_PP(16'h121B2,4);
TASK_PP(16'h121B3,4);
TASK_PP(16'h121B4,4);
TASK_PP(16'h121B5,4);
TASK_PP(16'h121B6,4);
TASK_PP(16'h121B7,4);
TASK_PP(16'h121B8,4);
TASK_PP(16'h121B9,4);
TASK_PP(16'h121BA,4);
TASK_PP(16'h121BB,4);
TASK_PP(16'h121BC,4);
TASK_PP(16'h121BD,4);
TASK_PP(16'h121BE,4);
TASK_PP(16'h121BF,4);
TASK_PP(16'h121C0,4);
TASK_PP(16'h121C1,4);
TASK_PP(16'h121C2,4);
TASK_PP(16'h121C3,4);
TASK_PP(16'h121C4,4);
TASK_PP(16'h121C5,4);
TASK_PP(16'h121C6,4);
TASK_PP(16'h121C7,4);
TASK_PP(16'h121C8,4);
TASK_PP(16'h121C9,4);
TASK_PP(16'h121CA,4);
TASK_PP(16'h121CB,4);
TASK_PP(16'h121CC,4);
TASK_PP(16'h121CD,4);
TASK_PP(16'h121CE,4);
TASK_PP(16'h121CF,4);
TASK_PP(16'h121D0,4);
TASK_PP(16'h121D1,4);
TASK_PP(16'h121D2,4);
TASK_PP(16'h121D3,4);
TASK_PP(16'h121D4,4);
TASK_PP(16'h121D5,4);
TASK_PP(16'h121D6,4);
TASK_PP(16'h121D7,4);
TASK_PP(16'h121D8,4);
TASK_PP(16'h121D9,4);
TASK_PP(16'h121DA,4);
TASK_PP(16'h121DB,4);
TASK_PP(16'h121DC,4);
TASK_PP(16'h121DD,4);
TASK_PP(16'h121DE,4);
TASK_PP(16'h121DF,4);
TASK_PP(16'h121E0,4);
TASK_PP(16'h121E1,4);
TASK_PP(16'h121E2,4);
TASK_PP(16'h121E3,4);
TASK_PP(16'h121E4,4);
TASK_PP(16'h121E5,4);
TASK_PP(16'h121E6,4);
TASK_PP(16'h121E7,4);
TASK_PP(16'h121E8,4);
TASK_PP(16'h121E9,4);
TASK_PP(16'h121EA,4);
TASK_PP(16'h121EB,4);
TASK_PP(16'h121EC,4);
TASK_PP(16'h121ED,4);
TASK_PP(16'h121EE,4);
TASK_PP(16'h121EF,4);
TASK_PP(16'h121F0,4);
TASK_PP(16'h121F1,4);
TASK_PP(16'h121F2,4);
TASK_PP(16'h121F3,4);
TASK_PP(16'h121F4,4);
TASK_PP(16'h121F5,4);
TASK_PP(16'h121F6,4);
TASK_PP(16'h121F7,4);
TASK_PP(16'h121F8,4);
TASK_PP(16'h121F9,4);
TASK_PP(16'h121FA,4);
TASK_PP(16'h121FB,4);
TASK_PP(16'h121FC,4);
TASK_PP(16'h121FD,4);
TASK_PP(16'h121FE,4);
TASK_PP(16'h121FF,4);
TASK_PP(16'h12200,4);
TASK_PP(16'h12201,4);
TASK_PP(16'h12202,4);
TASK_PP(16'h12203,4);
TASK_PP(16'h12204,4);
TASK_PP(16'h12205,4);
TASK_PP(16'h12206,4);
TASK_PP(16'h12207,4);
TASK_PP(16'h12208,4);
TASK_PP(16'h12209,4);
TASK_PP(16'h1220A,4);
TASK_PP(16'h1220B,4);
TASK_PP(16'h1220C,4);
TASK_PP(16'h1220D,4);
TASK_PP(16'h1220E,4);
TASK_PP(16'h1220F,4);
TASK_PP(16'h12210,4);
TASK_PP(16'h12211,4);
TASK_PP(16'h12212,4);
TASK_PP(16'h12213,4);
TASK_PP(16'h12214,4);
TASK_PP(16'h12215,4);
TASK_PP(16'h12216,4);
TASK_PP(16'h12217,4);
TASK_PP(16'h12218,4);
TASK_PP(16'h12219,4);
TASK_PP(16'h1221A,4);
TASK_PP(16'h1221B,4);
TASK_PP(16'h1221C,4);
TASK_PP(16'h1221D,4);
TASK_PP(16'h1221E,4);
TASK_PP(16'h1221F,4);
TASK_PP(16'h12220,4);
TASK_PP(16'h12221,4);
TASK_PP(16'h12222,4);
TASK_PP(16'h12223,4);
TASK_PP(16'h12224,4);
TASK_PP(16'h12225,4);
TASK_PP(16'h12226,4);
TASK_PP(16'h12227,4);
TASK_PP(16'h12228,4);
TASK_PP(16'h12229,4);
TASK_PP(16'h1222A,4);
TASK_PP(16'h1222B,4);
TASK_PP(16'h1222C,4);
TASK_PP(16'h1222D,4);
TASK_PP(16'h1222E,4);
TASK_PP(16'h1222F,4);
TASK_PP(16'h12230,4);
TASK_PP(16'h12231,4);
TASK_PP(16'h12232,4);
TASK_PP(16'h12233,4);
TASK_PP(16'h12234,4);
TASK_PP(16'h12235,4);
TASK_PP(16'h12236,4);
TASK_PP(16'h12237,4);
TASK_PP(16'h12238,4);
TASK_PP(16'h12239,4);
TASK_PP(16'h1223A,4);
TASK_PP(16'h1223B,4);
TASK_PP(16'h1223C,4);
TASK_PP(16'h1223D,4);
TASK_PP(16'h1223E,4);
TASK_PP(16'h1223F,4);
TASK_PP(16'h12240,4);
TASK_PP(16'h12241,4);
TASK_PP(16'h12242,4);
TASK_PP(16'h12243,4);
TASK_PP(16'h12244,4);
TASK_PP(16'h12245,4);
TASK_PP(16'h12246,4);
TASK_PP(16'h12247,4);
TASK_PP(16'h12248,4);
TASK_PP(16'h12249,4);
TASK_PP(16'h1224A,4);
TASK_PP(16'h1224B,4);
TASK_PP(16'h1224C,4);
TASK_PP(16'h1224D,4);
TASK_PP(16'h1224E,4);
TASK_PP(16'h1224F,4);
TASK_PP(16'h12250,4);
TASK_PP(16'h12251,4);
TASK_PP(16'h12252,4);
TASK_PP(16'h12253,4);
TASK_PP(16'h12254,4);
TASK_PP(16'h12255,4);
TASK_PP(16'h12256,4);
TASK_PP(16'h12257,4);
TASK_PP(16'h12258,4);
TASK_PP(16'h12259,4);
TASK_PP(16'h1225A,4);
TASK_PP(16'h1225B,4);
TASK_PP(16'h1225C,4);
TASK_PP(16'h1225D,4);
TASK_PP(16'h1225E,4);
TASK_PP(16'h1225F,4);
TASK_PP(16'h12260,4);
TASK_PP(16'h12261,4);
TASK_PP(16'h12262,4);
TASK_PP(16'h12263,4);
TASK_PP(16'h12264,4);
TASK_PP(16'h12265,4);
TASK_PP(16'h12266,4);
TASK_PP(16'h12267,4);
TASK_PP(16'h12268,4);
TASK_PP(16'h12269,4);
TASK_PP(16'h1226A,4);
TASK_PP(16'h1226B,4);
TASK_PP(16'h1226C,4);
TASK_PP(16'h1226D,4);
TASK_PP(16'h1226E,4);
TASK_PP(16'h1226F,4);
TASK_PP(16'h12270,4);
TASK_PP(16'h12271,4);
TASK_PP(16'h12272,4);
TASK_PP(16'h12273,4);
TASK_PP(16'h12274,4);
TASK_PP(16'h12275,4);
TASK_PP(16'h12276,4);
TASK_PP(16'h12277,4);
TASK_PP(16'h12278,4);
TASK_PP(16'h12279,4);
TASK_PP(16'h1227A,4);
TASK_PP(16'h1227B,4);
TASK_PP(16'h1227C,4);
TASK_PP(16'h1227D,4);
TASK_PP(16'h1227E,4);
TASK_PP(16'h1227F,4);
TASK_PP(16'h12280,4);
TASK_PP(16'h12281,4);
TASK_PP(16'h12282,4);
TASK_PP(16'h12283,4);
TASK_PP(16'h12284,4);
TASK_PP(16'h12285,4);
TASK_PP(16'h12286,4);
TASK_PP(16'h12287,4);
TASK_PP(16'h12288,4);
TASK_PP(16'h12289,4);
TASK_PP(16'h1228A,4);
TASK_PP(16'h1228B,4);
TASK_PP(16'h1228C,4);
TASK_PP(16'h1228D,4);
TASK_PP(16'h1228E,4);
TASK_PP(16'h1228F,4);
TASK_PP(16'h12290,4);
TASK_PP(16'h12291,4);
TASK_PP(16'h12292,4);
TASK_PP(16'h12293,4);
TASK_PP(16'h12294,4);
TASK_PP(16'h12295,4);
TASK_PP(16'h12296,4);
TASK_PP(16'h12297,4);
TASK_PP(16'h12298,4);
TASK_PP(16'h12299,4);
TASK_PP(16'h1229A,4);
TASK_PP(16'h1229B,4);
TASK_PP(16'h1229C,4);
TASK_PP(16'h1229D,4);
TASK_PP(16'h1229E,4);
TASK_PP(16'h1229F,4);
TASK_PP(16'h122A0,4);
TASK_PP(16'h122A1,4);
TASK_PP(16'h122A2,4);
TASK_PP(16'h122A3,4);
TASK_PP(16'h122A4,4);
TASK_PP(16'h122A5,4);
TASK_PP(16'h122A6,4);
TASK_PP(16'h122A7,4);
TASK_PP(16'h122A8,4);
TASK_PP(16'h122A9,4);
TASK_PP(16'h122AA,4);
TASK_PP(16'h122AB,4);
TASK_PP(16'h122AC,4);
TASK_PP(16'h122AD,4);
TASK_PP(16'h122AE,4);
TASK_PP(16'h122AF,4);
TASK_PP(16'h122B0,4);
TASK_PP(16'h122B1,4);
TASK_PP(16'h122B2,4);
TASK_PP(16'h122B3,4);
TASK_PP(16'h122B4,4);
TASK_PP(16'h122B5,4);
TASK_PP(16'h122B6,4);
TASK_PP(16'h122B7,4);
TASK_PP(16'h122B8,4);
TASK_PP(16'h122B9,4);
TASK_PP(16'h122BA,4);
TASK_PP(16'h122BB,4);
TASK_PP(16'h122BC,4);
TASK_PP(16'h122BD,4);
TASK_PP(16'h122BE,4);
TASK_PP(16'h122BF,4);
TASK_PP(16'h122C0,4);
TASK_PP(16'h122C1,4);
TASK_PP(16'h122C2,4);
TASK_PP(16'h122C3,4);
TASK_PP(16'h122C4,4);
TASK_PP(16'h122C5,4);
TASK_PP(16'h122C6,4);
TASK_PP(16'h122C7,4);
TASK_PP(16'h122C8,4);
TASK_PP(16'h122C9,4);
TASK_PP(16'h122CA,4);
TASK_PP(16'h122CB,4);
TASK_PP(16'h122CC,4);
TASK_PP(16'h122CD,4);
TASK_PP(16'h122CE,4);
TASK_PP(16'h122CF,4);
TASK_PP(16'h122D0,4);
TASK_PP(16'h122D1,4);
TASK_PP(16'h122D2,4);
TASK_PP(16'h122D3,4);
TASK_PP(16'h122D4,4);
TASK_PP(16'h122D5,4);
TASK_PP(16'h122D6,4);
TASK_PP(16'h122D7,4);
TASK_PP(16'h122D8,4);
TASK_PP(16'h122D9,4);
TASK_PP(16'h122DA,4);
TASK_PP(16'h122DB,4);
TASK_PP(16'h122DC,4);
TASK_PP(16'h122DD,4);
TASK_PP(16'h122DE,4);
TASK_PP(16'h122DF,4);
TASK_PP(16'h122E0,4);
TASK_PP(16'h122E1,4);
TASK_PP(16'h122E2,4);
TASK_PP(16'h122E3,4);
TASK_PP(16'h122E4,4);
TASK_PP(16'h122E5,4);
TASK_PP(16'h122E6,4);
TASK_PP(16'h122E7,4);
TASK_PP(16'h122E8,4);
TASK_PP(16'h122E9,4);
TASK_PP(16'h122EA,4);
TASK_PP(16'h122EB,4);
TASK_PP(16'h122EC,4);
TASK_PP(16'h122ED,4);
TASK_PP(16'h122EE,4);
TASK_PP(16'h122EF,4);
TASK_PP(16'h122F0,4);
TASK_PP(16'h122F1,4);
TASK_PP(16'h122F2,4);
TASK_PP(16'h122F3,4);
TASK_PP(16'h122F4,4);
TASK_PP(16'h122F5,4);
TASK_PP(16'h122F6,4);
TASK_PP(16'h122F7,4);
TASK_PP(16'h122F8,4);
TASK_PP(16'h122F9,4);
TASK_PP(16'h122FA,4);
TASK_PP(16'h122FB,4);
TASK_PP(16'h122FC,4);
TASK_PP(16'h122FD,4);
TASK_PP(16'h122FE,4);
TASK_PP(16'h122FF,4);
TASK_PP(16'h12300,4);
TASK_PP(16'h12301,4);
TASK_PP(16'h12302,4);
TASK_PP(16'h12303,4);
TASK_PP(16'h12304,4);
TASK_PP(16'h12305,4);
TASK_PP(16'h12306,4);
TASK_PP(16'h12307,4);
TASK_PP(16'h12308,4);
TASK_PP(16'h12309,4);
TASK_PP(16'h1230A,4);
TASK_PP(16'h1230B,4);
TASK_PP(16'h1230C,4);
TASK_PP(16'h1230D,4);
TASK_PP(16'h1230E,4);
TASK_PP(16'h1230F,4);
TASK_PP(16'h12310,4);
TASK_PP(16'h12311,4);
TASK_PP(16'h12312,4);
TASK_PP(16'h12313,4);
TASK_PP(16'h12314,4);
TASK_PP(16'h12315,4);
TASK_PP(16'h12316,4);
TASK_PP(16'h12317,4);
TASK_PP(16'h12318,4);
TASK_PP(16'h12319,4);
TASK_PP(16'h1231A,4);
TASK_PP(16'h1231B,4);
TASK_PP(16'h1231C,4);
TASK_PP(16'h1231D,4);
TASK_PP(16'h1231E,4);
TASK_PP(16'h1231F,4);
TASK_PP(16'h12320,4);
TASK_PP(16'h12321,4);
TASK_PP(16'h12322,4);
TASK_PP(16'h12323,4);
TASK_PP(16'h12324,4);
TASK_PP(16'h12325,4);
TASK_PP(16'h12326,4);
TASK_PP(16'h12327,4);
TASK_PP(16'h12328,4);
TASK_PP(16'h12329,4);
TASK_PP(16'h1232A,4);
TASK_PP(16'h1232B,4);
TASK_PP(16'h1232C,4);
TASK_PP(16'h1232D,4);
TASK_PP(16'h1232E,4);
TASK_PP(16'h1232F,4);
TASK_PP(16'h12330,4);
TASK_PP(16'h12331,4);
TASK_PP(16'h12332,4);
TASK_PP(16'h12333,4);
TASK_PP(16'h12334,4);
TASK_PP(16'h12335,4);
TASK_PP(16'h12336,4);
TASK_PP(16'h12337,4);
TASK_PP(16'h12338,4);
TASK_PP(16'h12339,4);
TASK_PP(16'h1233A,4);
TASK_PP(16'h1233B,4);
TASK_PP(16'h1233C,4);
TASK_PP(16'h1233D,4);
TASK_PP(16'h1233E,4);
TASK_PP(16'h1233F,4);
TASK_PP(16'h12340,4);
TASK_PP(16'h12341,4);
TASK_PP(16'h12342,4);
TASK_PP(16'h12343,4);
TASK_PP(16'h12344,4);
TASK_PP(16'h12345,4);
TASK_PP(16'h12346,4);
TASK_PP(16'h12347,4);
TASK_PP(16'h12348,4);
TASK_PP(16'h12349,4);
TASK_PP(16'h1234A,4);
TASK_PP(16'h1234B,4);
TASK_PP(16'h1234C,4);
TASK_PP(16'h1234D,4);
TASK_PP(16'h1234E,4);
TASK_PP(16'h1234F,4);
TASK_PP(16'h12350,4);
TASK_PP(16'h12351,4);
TASK_PP(16'h12352,4);
TASK_PP(16'h12353,4);
TASK_PP(16'h12354,4);
TASK_PP(16'h12355,4);
TASK_PP(16'h12356,4);
TASK_PP(16'h12357,4);
TASK_PP(16'h12358,4);
TASK_PP(16'h12359,4);
TASK_PP(16'h1235A,4);
TASK_PP(16'h1235B,4);
TASK_PP(16'h1235C,4);
TASK_PP(16'h1235D,4);
TASK_PP(16'h1235E,4);
TASK_PP(16'h1235F,4);
TASK_PP(16'h12360,4);
TASK_PP(16'h12361,4);
TASK_PP(16'h12362,4);
TASK_PP(16'h12363,4);
TASK_PP(16'h12364,4);
TASK_PP(16'h12365,4);
TASK_PP(16'h12366,4);
TASK_PP(16'h12367,4);
TASK_PP(16'h12368,4);
TASK_PP(16'h12369,4);
TASK_PP(16'h1236A,4);
TASK_PP(16'h1236B,4);
TASK_PP(16'h1236C,4);
TASK_PP(16'h1236D,4);
TASK_PP(16'h1236E,4);
TASK_PP(16'h1236F,4);
TASK_PP(16'h12370,4);
TASK_PP(16'h12371,4);
TASK_PP(16'h12372,4);
TASK_PP(16'h12373,4);
TASK_PP(16'h12374,4);
TASK_PP(16'h12375,4);
TASK_PP(16'h12376,4);
TASK_PP(16'h12377,4);
TASK_PP(16'h12378,4);
TASK_PP(16'h12379,4);
TASK_PP(16'h1237A,4);
TASK_PP(16'h1237B,4);
TASK_PP(16'h1237C,4);
TASK_PP(16'h1237D,4);
TASK_PP(16'h1237E,4);
TASK_PP(16'h1237F,4);
TASK_PP(16'h12380,4);
TASK_PP(16'h12381,4);
TASK_PP(16'h12382,4);
TASK_PP(16'h12383,4);
TASK_PP(16'h12384,4);
TASK_PP(16'h12385,4);
TASK_PP(16'h12386,4);
TASK_PP(16'h12387,4);
TASK_PP(16'h12388,4);
TASK_PP(16'h12389,4);
TASK_PP(16'h1238A,4);
TASK_PP(16'h1238B,4);
TASK_PP(16'h1238C,4);
TASK_PP(16'h1238D,4);
TASK_PP(16'h1238E,4);
TASK_PP(16'h1238F,4);
TASK_PP(16'h12390,4);
TASK_PP(16'h12391,4);
TASK_PP(16'h12392,4);
TASK_PP(16'h12393,4);
TASK_PP(16'h12394,4);
TASK_PP(16'h12395,4);
TASK_PP(16'h12396,4);
TASK_PP(16'h12397,4);
TASK_PP(16'h12398,4);
TASK_PP(16'h12399,4);
TASK_PP(16'h1239A,4);
TASK_PP(16'h1239B,4);
TASK_PP(16'h1239C,4);
TASK_PP(16'h1239D,4);
TASK_PP(16'h1239E,4);
TASK_PP(16'h1239F,4);
TASK_PP(16'h123A0,4);
TASK_PP(16'h123A1,4);
TASK_PP(16'h123A2,4);
TASK_PP(16'h123A3,4);
TASK_PP(16'h123A4,4);
TASK_PP(16'h123A5,4);
TASK_PP(16'h123A6,4);
TASK_PP(16'h123A7,4);
TASK_PP(16'h123A8,4);
TASK_PP(16'h123A9,4);
TASK_PP(16'h123AA,4);
TASK_PP(16'h123AB,4);
TASK_PP(16'h123AC,4);
TASK_PP(16'h123AD,4);
TASK_PP(16'h123AE,4);
TASK_PP(16'h123AF,4);
TASK_PP(16'h123B0,4);
TASK_PP(16'h123B1,4);
TASK_PP(16'h123B2,4);
TASK_PP(16'h123B3,4);
TASK_PP(16'h123B4,4);
TASK_PP(16'h123B5,4);
TASK_PP(16'h123B6,4);
TASK_PP(16'h123B7,4);
TASK_PP(16'h123B8,4);
TASK_PP(16'h123B9,4);
TASK_PP(16'h123BA,4);
TASK_PP(16'h123BB,4);
TASK_PP(16'h123BC,4);
TASK_PP(16'h123BD,4);
TASK_PP(16'h123BE,4);
TASK_PP(16'h123BF,4);
TASK_PP(16'h123C0,4);
TASK_PP(16'h123C1,4);
TASK_PP(16'h123C2,4);
TASK_PP(16'h123C3,4);
TASK_PP(16'h123C4,4);
TASK_PP(16'h123C5,4);
TASK_PP(16'h123C6,4);
TASK_PP(16'h123C7,4);
TASK_PP(16'h123C8,4);
TASK_PP(16'h123C9,4);
TASK_PP(16'h123CA,4);
TASK_PP(16'h123CB,4);
TASK_PP(16'h123CC,4);
TASK_PP(16'h123CD,4);
TASK_PP(16'h123CE,4);
TASK_PP(16'h123CF,4);
TASK_PP(16'h123D0,4);
TASK_PP(16'h123D1,4);
TASK_PP(16'h123D2,4);
TASK_PP(16'h123D3,4);
TASK_PP(16'h123D4,4);
TASK_PP(16'h123D5,4);
TASK_PP(16'h123D6,4);
TASK_PP(16'h123D7,4);
TASK_PP(16'h123D8,4);
TASK_PP(16'h123D9,4);
TASK_PP(16'h123DA,4);
TASK_PP(16'h123DB,4);
TASK_PP(16'h123DC,4);
TASK_PP(16'h123DD,4);
TASK_PP(16'h123DE,4);
TASK_PP(16'h123DF,4);
TASK_PP(16'h123E0,4);
TASK_PP(16'h123E1,4);
TASK_PP(16'h123E2,4);
TASK_PP(16'h123E3,4);
TASK_PP(16'h123E4,4);
TASK_PP(16'h123E5,4);
TASK_PP(16'h123E6,4);
TASK_PP(16'h123E7,4);
TASK_PP(16'h123E8,4);
TASK_PP(16'h123E9,4);
TASK_PP(16'h123EA,4);
TASK_PP(16'h123EB,4);
TASK_PP(16'h123EC,4);
TASK_PP(16'h123ED,4);
TASK_PP(16'h123EE,4);
TASK_PP(16'h123EF,4);
TASK_PP(16'h123F0,4);
TASK_PP(16'h123F1,4);
TASK_PP(16'h123F2,4);
TASK_PP(16'h123F3,4);
TASK_PP(16'h123F4,4);
TASK_PP(16'h123F5,4);
TASK_PP(16'h123F6,4);
TASK_PP(16'h123F7,4);
TASK_PP(16'h123F8,4);
TASK_PP(16'h123F9,4);
TASK_PP(16'h123FA,4);
TASK_PP(16'h123FB,4);
TASK_PP(16'h123FC,4);
TASK_PP(16'h123FD,4);
TASK_PP(16'h123FE,4);
TASK_PP(16'h123FF,4);
TASK_PP(16'h12400,4);
TASK_PP(16'h12401,4);
TASK_PP(16'h12402,4);
TASK_PP(16'h12403,4);
TASK_PP(16'h12404,4);
TASK_PP(16'h12405,4);
TASK_PP(16'h12406,4);
TASK_PP(16'h12407,4);
TASK_PP(16'h12408,4);
TASK_PP(16'h12409,4);
TASK_PP(16'h1240A,4);
TASK_PP(16'h1240B,4);
TASK_PP(16'h1240C,4);
TASK_PP(16'h1240D,4);
TASK_PP(16'h1240E,4);
TASK_PP(16'h1240F,4);
TASK_PP(16'h12410,4);
TASK_PP(16'h12411,4);
TASK_PP(16'h12412,4);
TASK_PP(16'h12413,4);
TASK_PP(16'h12414,4);
TASK_PP(16'h12415,4);
TASK_PP(16'h12416,4);
TASK_PP(16'h12417,4);
TASK_PP(16'h12418,4);
TASK_PP(16'h12419,4);
TASK_PP(16'h1241A,4);
TASK_PP(16'h1241B,4);
TASK_PP(16'h1241C,4);
TASK_PP(16'h1241D,4);
TASK_PP(16'h1241E,4);
TASK_PP(16'h1241F,4);
TASK_PP(16'h12420,4);
TASK_PP(16'h12421,4);
TASK_PP(16'h12422,4);
TASK_PP(16'h12423,4);
TASK_PP(16'h12424,4);
TASK_PP(16'h12425,4);
TASK_PP(16'h12426,4);
TASK_PP(16'h12427,4);
TASK_PP(16'h12428,4);
TASK_PP(16'h12429,4);
TASK_PP(16'h1242A,4);
TASK_PP(16'h1242B,4);
TASK_PP(16'h1242C,4);
TASK_PP(16'h1242D,4);
TASK_PP(16'h1242E,4);
TASK_PP(16'h1242F,4);
TASK_PP(16'h12430,4);
TASK_PP(16'h12431,4);
TASK_PP(16'h12432,4);
TASK_PP(16'h12433,4);
TASK_PP(16'h12434,4);
TASK_PP(16'h12435,4);
TASK_PP(16'h12436,4);
TASK_PP(16'h12437,4);
TASK_PP(16'h12438,4);
TASK_PP(16'h12439,4);
TASK_PP(16'h1243A,4);
TASK_PP(16'h1243B,4);
TASK_PP(16'h1243C,4);
TASK_PP(16'h1243D,4);
TASK_PP(16'h1243E,4);
TASK_PP(16'h1243F,4);
TASK_PP(16'h12440,4);
TASK_PP(16'h12441,4);
TASK_PP(16'h12442,4);
TASK_PP(16'h12443,4);
TASK_PP(16'h12444,4);
TASK_PP(16'h12445,4);
TASK_PP(16'h12446,4);
TASK_PP(16'h12447,4);
TASK_PP(16'h12448,4);
TASK_PP(16'h12449,4);
TASK_PP(16'h1244A,4);
TASK_PP(16'h1244B,4);
TASK_PP(16'h1244C,4);
TASK_PP(16'h1244D,4);
TASK_PP(16'h1244E,4);
TASK_PP(16'h1244F,4);
TASK_PP(16'h12450,4);
TASK_PP(16'h12451,4);
TASK_PP(16'h12452,4);
TASK_PP(16'h12453,4);
TASK_PP(16'h12454,4);
TASK_PP(16'h12455,4);
TASK_PP(16'h12456,4);
TASK_PP(16'h12457,4);
TASK_PP(16'h12458,4);
TASK_PP(16'h12459,4);
TASK_PP(16'h1245A,4);
TASK_PP(16'h1245B,4);
TASK_PP(16'h1245C,4);
TASK_PP(16'h1245D,4);
TASK_PP(16'h1245E,4);
TASK_PP(16'h1245F,4);
TASK_PP(16'h12460,4);
TASK_PP(16'h12461,4);
TASK_PP(16'h12462,4);
TASK_PP(16'h12463,4);
TASK_PP(16'h12464,4);
TASK_PP(16'h12465,4);
TASK_PP(16'h12466,4);
TASK_PP(16'h12467,4);
TASK_PP(16'h12468,4);
TASK_PP(16'h12469,4);
TASK_PP(16'h1246A,4);
TASK_PP(16'h1246B,4);
TASK_PP(16'h1246C,4);
TASK_PP(16'h1246D,4);
TASK_PP(16'h1246E,4);
TASK_PP(16'h1246F,4);
TASK_PP(16'h12470,4);
TASK_PP(16'h12471,4);
TASK_PP(16'h12472,4);
TASK_PP(16'h12473,4);
TASK_PP(16'h12474,4);
TASK_PP(16'h12475,4);
TASK_PP(16'h12476,4);
TASK_PP(16'h12477,4);
TASK_PP(16'h12478,4);
TASK_PP(16'h12479,4);
TASK_PP(16'h1247A,4);
TASK_PP(16'h1247B,4);
TASK_PP(16'h1247C,4);
TASK_PP(16'h1247D,4);
TASK_PP(16'h1247E,4);
TASK_PP(16'h1247F,4);
TASK_PP(16'h12480,4);
TASK_PP(16'h12481,4);
TASK_PP(16'h12482,4);
TASK_PP(16'h12483,4);
TASK_PP(16'h12484,4);
TASK_PP(16'h12485,4);
TASK_PP(16'h12486,4);
TASK_PP(16'h12487,4);
TASK_PP(16'h12488,4);
TASK_PP(16'h12489,4);
TASK_PP(16'h1248A,4);
TASK_PP(16'h1248B,4);
TASK_PP(16'h1248C,4);
TASK_PP(16'h1248D,4);
TASK_PP(16'h1248E,4);
TASK_PP(16'h1248F,4);
TASK_PP(16'h12490,4);
TASK_PP(16'h12491,4);
TASK_PP(16'h12492,4);
TASK_PP(16'h12493,4);
TASK_PP(16'h12494,4);
TASK_PP(16'h12495,4);
TASK_PP(16'h12496,4);
TASK_PP(16'h12497,4);
TASK_PP(16'h12498,4);
TASK_PP(16'h12499,4);
TASK_PP(16'h1249A,4);
TASK_PP(16'h1249B,4);
TASK_PP(16'h1249C,4);
TASK_PP(16'h1249D,4);
TASK_PP(16'h1249E,4);
TASK_PP(16'h1249F,4);
TASK_PP(16'h124A0,4);
TASK_PP(16'h124A1,4);
TASK_PP(16'h124A2,4);
TASK_PP(16'h124A3,4);
TASK_PP(16'h124A4,4);
TASK_PP(16'h124A5,4);
TASK_PP(16'h124A6,4);
TASK_PP(16'h124A7,4);
TASK_PP(16'h124A8,4);
TASK_PP(16'h124A9,4);
TASK_PP(16'h124AA,4);
TASK_PP(16'h124AB,4);
TASK_PP(16'h124AC,4);
TASK_PP(16'h124AD,4);
TASK_PP(16'h124AE,4);
TASK_PP(16'h124AF,4);
TASK_PP(16'h124B0,4);
TASK_PP(16'h124B1,4);
TASK_PP(16'h124B2,4);
TASK_PP(16'h124B3,4);
TASK_PP(16'h124B4,4);
TASK_PP(16'h124B5,4);
TASK_PP(16'h124B6,4);
TASK_PP(16'h124B7,4);
TASK_PP(16'h124B8,4);
TASK_PP(16'h124B9,4);
TASK_PP(16'h124BA,4);
TASK_PP(16'h124BB,4);
TASK_PP(16'h124BC,4);
TASK_PP(16'h124BD,4);
TASK_PP(16'h124BE,4);
TASK_PP(16'h124BF,4);
TASK_PP(16'h124C0,4);
TASK_PP(16'h124C1,4);
TASK_PP(16'h124C2,4);
TASK_PP(16'h124C3,4);
TASK_PP(16'h124C4,4);
TASK_PP(16'h124C5,4);
TASK_PP(16'h124C6,4);
TASK_PP(16'h124C7,4);
TASK_PP(16'h124C8,4);
TASK_PP(16'h124C9,4);
TASK_PP(16'h124CA,4);
TASK_PP(16'h124CB,4);
TASK_PP(16'h124CC,4);
TASK_PP(16'h124CD,4);
TASK_PP(16'h124CE,4);
TASK_PP(16'h124CF,4);
TASK_PP(16'h124D0,4);
TASK_PP(16'h124D1,4);
TASK_PP(16'h124D2,4);
TASK_PP(16'h124D3,4);
TASK_PP(16'h124D4,4);
TASK_PP(16'h124D5,4);
TASK_PP(16'h124D6,4);
TASK_PP(16'h124D7,4);
TASK_PP(16'h124D8,4);
TASK_PP(16'h124D9,4);
TASK_PP(16'h124DA,4);
TASK_PP(16'h124DB,4);
TASK_PP(16'h124DC,4);
TASK_PP(16'h124DD,4);
TASK_PP(16'h124DE,4);
TASK_PP(16'h124DF,4);
TASK_PP(16'h124E0,4);
TASK_PP(16'h124E1,4);
TASK_PP(16'h124E2,4);
TASK_PP(16'h124E3,4);
TASK_PP(16'h124E4,4);
TASK_PP(16'h124E5,4);
TASK_PP(16'h124E6,4);
TASK_PP(16'h124E7,4);
TASK_PP(16'h124E8,4);
TASK_PP(16'h124E9,4);
TASK_PP(16'h124EA,4);
TASK_PP(16'h124EB,4);
TASK_PP(16'h124EC,4);
TASK_PP(16'h124ED,4);
TASK_PP(16'h124EE,4);
TASK_PP(16'h124EF,4);
TASK_PP(16'h124F0,4);
TASK_PP(16'h124F1,4);
TASK_PP(16'h124F2,4);
TASK_PP(16'h124F3,4);
TASK_PP(16'h124F4,4);
TASK_PP(16'h124F5,4);
TASK_PP(16'h124F6,4);
TASK_PP(16'h124F7,4);
TASK_PP(16'h124F8,4);
TASK_PP(16'h124F9,4);
TASK_PP(16'h124FA,4);
TASK_PP(16'h124FB,4);
TASK_PP(16'h124FC,4);
TASK_PP(16'h124FD,4);
TASK_PP(16'h124FE,4);
TASK_PP(16'h124FF,4);
TASK_PP(16'h12500,4);
TASK_PP(16'h12501,4);
TASK_PP(16'h12502,4);
TASK_PP(16'h12503,4);
TASK_PP(16'h12504,4);
TASK_PP(16'h12505,4);
TASK_PP(16'h12506,4);
TASK_PP(16'h12507,4);
TASK_PP(16'h12508,4);
TASK_PP(16'h12509,4);
TASK_PP(16'h1250A,4);
TASK_PP(16'h1250B,4);
TASK_PP(16'h1250C,4);
TASK_PP(16'h1250D,4);
TASK_PP(16'h1250E,4);
TASK_PP(16'h1250F,4);
TASK_PP(16'h12510,4);
TASK_PP(16'h12511,4);
TASK_PP(16'h12512,4);
TASK_PP(16'h12513,4);
TASK_PP(16'h12514,4);
TASK_PP(16'h12515,4);
TASK_PP(16'h12516,4);
TASK_PP(16'h12517,4);
TASK_PP(16'h12518,4);
TASK_PP(16'h12519,4);
TASK_PP(16'h1251A,4);
TASK_PP(16'h1251B,4);
TASK_PP(16'h1251C,4);
TASK_PP(16'h1251D,4);
TASK_PP(16'h1251E,4);
TASK_PP(16'h1251F,4);
TASK_PP(16'h12520,4);
TASK_PP(16'h12521,4);
TASK_PP(16'h12522,4);
TASK_PP(16'h12523,4);
TASK_PP(16'h12524,4);
TASK_PP(16'h12525,4);
TASK_PP(16'h12526,4);
TASK_PP(16'h12527,4);
TASK_PP(16'h12528,4);
TASK_PP(16'h12529,4);
TASK_PP(16'h1252A,4);
TASK_PP(16'h1252B,4);
TASK_PP(16'h1252C,4);
TASK_PP(16'h1252D,4);
TASK_PP(16'h1252E,4);
TASK_PP(16'h1252F,4);
TASK_PP(16'h12530,4);
TASK_PP(16'h12531,4);
TASK_PP(16'h12532,4);
TASK_PP(16'h12533,4);
TASK_PP(16'h12534,4);
TASK_PP(16'h12535,4);
TASK_PP(16'h12536,4);
TASK_PP(16'h12537,4);
TASK_PP(16'h12538,4);
TASK_PP(16'h12539,4);
TASK_PP(16'h1253A,4);
TASK_PP(16'h1253B,4);
TASK_PP(16'h1253C,4);
TASK_PP(16'h1253D,4);
TASK_PP(16'h1253E,4);
TASK_PP(16'h1253F,4);
TASK_PP(16'h12540,4);
TASK_PP(16'h12541,4);
TASK_PP(16'h12542,4);
TASK_PP(16'h12543,4);
TASK_PP(16'h12544,4);
TASK_PP(16'h12545,4);
TASK_PP(16'h12546,4);
TASK_PP(16'h12547,4);
TASK_PP(16'h12548,4);
TASK_PP(16'h12549,4);
TASK_PP(16'h1254A,4);
TASK_PP(16'h1254B,4);
TASK_PP(16'h1254C,4);
TASK_PP(16'h1254D,4);
TASK_PP(16'h1254E,4);
TASK_PP(16'h1254F,4);
TASK_PP(16'h12550,4);
TASK_PP(16'h12551,4);
TASK_PP(16'h12552,4);
TASK_PP(16'h12553,4);
TASK_PP(16'h12554,4);
TASK_PP(16'h12555,4);
TASK_PP(16'h12556,4);
TASK_PP(16'h12557,4);
TASK_PP(16'h12558,4);
TASK_PP(16'h12559,4);
TASK_PP(16'h1255A,4);
TASK_PP(16'h1255B,4);
TASK_PP(16'h1255C,4);
TASK_PP(16'h1255D,4);
TASK_PP(16'h1255E,4);
TASK_PP(16'h1255F,4);
TASK_PP(16'h12560,4);
TASK_PP(16'h12561,4);
TASK_PP(16'h12562,4);
TASK_PP(16'h12563,4);
TASK_PP(16'h12564,4);
TASK_PP(16'h12565,4);
TASK_PP(16'h12566,4);
TASK_PP(16'h12567,4);
TASK_PP(16'h12568,4);
TASK_PP(16'h12569,4);
TASK_PP(16'h1256A,4);
TASK_PP(16'h1256B,4);
TASK_PP(16'h1256C,4);
TASK_PP(16'h1256D,4);
TASK_PP(16'h1256E,4);
TASK_PP(16'h1256F,4);
TASK_PP(16'h12570,4);
TASK_PP(16'h12571,4);
TASK_PP(16'h12572,4);
TASK_PP(16'h12573,4);
TASK_PP(16'h12574,4);
TASK_PP(16'h12575,4);
TASK_PP(16'h12576,4);
TASK_PP(16'h12577,4);
TASK_PP(16'h12578,4);
TASK_PP(16'h12579,4);
TASK_PP(16'h1257A,4);
TASK_PP(16'h1257B,4);
TASK_PP(16'h1257C,4);
TASK_PP(16'h1257D,4);
TASK_PP(16'h1257E,4);
TASK_PP(16'h1257F,4);
TASK_PP(16'h12580,4);
TASK_PP(16'h12581,4);
TASK_PP(16'h12582,4);
TASK_PP(16'h12583,4);
TASK_PP(16'h12584,4);
TASK_PP(16'h12585,4);
TASK_PP(16'h12586,4);
TASK_PP(16'h12587,4);
TASK_PP(16'h12588,4);
TASK_PP(16'h12589,4);
TASK_PP(16'h1258A,4);
TASK_PP(16'h1258B,4);
TASK_PP(16'h1258C,4);
TASK_PP(16'h1258D,4);
TASK_PP(16'h1258E,4);
TASK_PP(16'h1258F,4);
TASK_PP(16'h12590,4);
TASK_PP(16'h12591,4);
TASK_PP(16'h12592,4);
TASK_PP(16'h12593,4);
TASK_PP(16'h12594,4);
TASK_PP(16'h12595,4);
TASK_PP(16'h12596,4);
TASK_PP(16'h12597,4);
TASK_PP(16'h12598,4);
TASK_PP(16'h12599,4);
TASK_PP(16'h1259A,4);
TASK_PP(16'h1259B,4);
TASK_PP(16'h1259C,4);
TASK_PP(16'h1259D,4);
TASK_PP(16'h1259E,4);
TASK_PP(16'h1259F,4);
TASK_PP(16'h125A0,4);
TASK_PP(16'h125A1,4);
TASK_PP(16'h125A2,4);
TASK_PP(16'h125A3,4);
TASK_PP(16'h125A4,4);
TASK_PP(16'h125A5,4);
TASK_PP(16'h125A6,4);
TASK_PP(16'h125A7,4);
TASK_PP(16'h125A8,4);
TASK_PP(16'h125A9,4);
TASK_PP(16'h125AA,4);
TASK_PP(16'h125AB,4);
TASK_PP(16'h125AC,4);
TASK_PP(16'h125AD,4);
TASK_PP(16'h125AE,4);
TASK_PP(16'h125AF,4);
TASK_PP(16'h125B0,4);
TASK_PP(16'h125B1,4);
TASK_PP(16'h125B2,4);
TASK_PP(16'h125B3,4);
TASK_PP(16'h125B4,4);
TASK_PP(16'h125B5,4);
TASK_PP(16'h125B6,4);
TASK_PP(16'h125B7,4);
TASK_PP(16'h125B8,4);
TASK_PP(16'h125B9,4);
TASK_PP(16'h125BA,4);
TASK_PP(16'h125BB,4);
TASK_PP(16'h125BC,4);
TASK_PP(16'h125BD,4);
TASK_PP(16'h125BE,4);
TASK_PP(16'h125BF,4);
TASK_PP(16'h125C0,4);
TASK_PP(16'h125C1,4);
TASK_PP(16'h125C2,4);
TASK_PP(16'h125C3,4);
TASK_PP(16'h125C4,4);
TASK_PP(16'h125C5,4);
TASK_PP(16'h125C6,4);
TASK_PP(16'h125C7,4);
TASK_PP(16'h125C8,4);
TASK_PP(16'h125C9,4);
TASK_PP(16'h125CA,4);
TASK_PP(16'h125CB,4);
TASK_PP(16'h125CC,4);
TASK_PP(16'h125CD,4);
TASK_PP(16'h125CE,4);
TASK_PP(16'h125CF,4);
TASK_PP(16'h125D0,4);
TASK_PP(16'h125D1,4);
TASK_PP(16'h125D2,4);
TASK_PP(16'h125D3,4);
TASK_PP(16'h125D4,4);
TASK_PP(16'h125D5,4);
TASK_PP(16'h125D6,4);
TASK_PP(16'h125D7,4);
TASK_PP(16'h125D8,4);
TASK_PP(16'h125D9,4);
TASK_PP(16'h125DA,4);
TASK_PP(16'h125DB,4);
TASK_PP(16'h125DC,4);
TASK_PP(16'h125DD,4);
TASK_PP(16'h125DE,4);
TASK_PP(16'h125DF,4);
TASK_PP(16'h125E0,4);
TASK_PP(16'h125E1,4);
TASK_PP(16'h125E2,4);
TASK_PP(16'h125E3,4);
TASK_PP(16'h125E4,4);
TASK_PP(16'h125E5,4);
TASK_PP(16'h125E6,4);
TASK_PP(16'h125E7,4);
TASK_PP(16'h125E8,4);
TASK_PP(16'h125E9,4);
TASK_PP(16'h125EA,4);
TASK_PP(16'h125EB,4);
TASK_PP(16'h125EC,4);
TASK_PP(16'h125ED,4);
TASK_PP(16'h125EE,4);
TASK_PP(16'h125EF,4);
TASK_PP(16'h125F0,4);
TASK_PP(16'h125F1,4);
TASK_PP(16'h125F2,4);
TASK_PP(16'h125F3,4);
TASK_PP(16'h125F4,4);
TASK_PP(16'h125F5,4);
TASK_PP(16'h125F6,4);
TASK_PP(16'h125F7,4);
TASK_PP(16'h125F8,4);
TASK_PP(16'h125F9,4);
TASK_PP(16'h125FA,4);
TASK_PP(16'h125FB,4);
TASK_PP(16'h125FC,4);
TASK_PP(16'h125FD,4);
TASK_PP(16'h125FE,4);
TASK_PP(16'h125FF,4);
TASK_PP(16'h12600,4);
TASK_PP(16'h12601,4);
TASK_PP(16'h12602,4);
TASK_PP(16'h12603,4);
TASK_PP(16'h12604,4);
TASK_PP(16'h12605,4);
TASK_PP(16'h12606,4);
TASK_PP(16'h12607,4);
TASK_PP(16'h12608,4);
TASK_PP(16'h12609,4);
TASK_PP(16'h1260A,4);
TASK_PP(16'h1260B,4);
TASK_PP(16'h1260C,4);
TASK_PP(16'h1260D,4);
TASK_PP(16'h1260E,4);
TASK_PP(16'h1260F,4);
TASK_PP(16'h12610,4);
TASK_PP(16'h12611,4);
TASK_PP(16'h12612,4);
TASK_PP(16'h12613,4);
TASK_PP(16'h12614,4);
TASK_PP(16'h12615,4);
TASK_PP(16'h12616,4);
TASK_PP(16'h12617,4);
TASK_PP(16'h12618,4);
TASK_PP(16'h12619,4);
TASK_PP(16'h1261A,4);
TASK_PP(16'h1261B,4);
TASK_PP(16'h1261C,4);
TASK_PP(16'h1261D,4);
TASK_PP(16'h1261E,4);
TASK_PP(16'h1261F,4);
TASK_PP(16'h12620,4);
TASK_PP(16'h12621,4);
TASK_PP(16'h12622,4);
TASK_PP(16'h12623,4);
TASK_PP(16'h12624,4);
TASK_PP(16'h12625,4);
TASK_PP(16'h12626,4);
TASK_PP(16'h12627,4);
TASK_PP(16'h12628,4);
TASK_PP(16'h12629,4);
TASK_PP(16'h1262A,4);
TASK_PP(16'h1262B,4);
TASK_PP(16'h1262C,4);
TASK_PP(16'h1262D,4);
TASK_PP(16'h1262E,4);
TASK_PP(16'h1262F,4);
TASK_PP(16'h12630,4);
TASK_PP(16'h12631,4);
TASK_PP(16'h12632,4);
TASK_PP(16'h12633,4);
TASK_PP(16'h12634,4);
TASK_PP(16'h12635,4);
TASK_PP(16'h12636,4);
TASK_PP(16'h12637,4);
TASK_PP(16'h12638,4);
TASK_PP(16'h12639,4);
TASK_PP(16'h1263A,4);
TASK_PP(16'h1263B,4);
TASK_PP(16'h1263C,4);
TASK_PP(16'h1263D,4);
TASK_PP(16'h1263E,4);
TASK_PP(16'h1263F,4);
TASK_PP(16'h12640,4);
TASK_PP(16'h12641,4);
TASK_PP(16'h12642,4);
TASK_PP(16'h12643,4);
TASK_PP(16'h12644,4);
TASK_PP(16'h12645,4);
TASK_PP(16'h12646,4);
TASK_PP(16'h12647,4);
TASK_PP(16'h12648,4);
TASK_PP(16'h12649,4);
TASK_PP(16'h1264A,4);
TASK_PP(16'h1264B,4);
TASK_PP(16'h1264C,4);
TASK_PP(16'h1264D,4);
TASK_PP(16'h1264E,4);
TASK_PP(16'h1264F,4);
TASK_PP(16'h12650,4);
TASK_PP(16'h12651,4);
TASK_PP(16'h12652,4);
TASK_PP(16'h12653,4);
TASK_PP(16'h12654,4);
TASK_PP(16'h12655,4);
TASK_PP(16'h12656,4);
TASK_PP(16'h12657,4);
TASK_PP(16'h12658,4);
TASK_PP(16'h12659,4);
TASK_PP(16'h1265A,4);
TASK_PP(16'h1265B,4);
TASK_PP(16'h1265C,4);
TASK_PP(16'h1265D,4);
TASK_PP(16'h1265E,4);
TASK_PP(16'h1265F,4);
TASK_PP(16'h12660,4);
TASK_PP(16'h12661,4);
TASK_PP(16'h12662,4);
TASK_PP(16'h12663,4);
TASK_PP(16'h12664,4);
TASK_PP(16'h12665,4);
TASK_PP(16'h12666,4);
TASK_PP(16'h12667,4);
TASK_PP(16'h12668,4);
TASK_PP(16'h12669,4);
TASK_PP(16'h1266A,4);
TASK_PP(16'h1266B,4);
TASK_PP(16'h1266C,4);
TASK_PP(16'h1266D,4);
TASK_PP(16'h1266E,4);
TASK_PP(16'h1266F,4);
TASK_PP(16'h12670,4);
TASK_PP(16'h12671,4);
TASK_PP(16'h12672,4);
TASK_PP(16'h12673,4);
TASK_PP(16'h12674,4);
TASK_PP(16'h12675,4);
TASK_PP(16'h12676,4);
TASK_PP(16'h12677,4);
TASK_PP(16'h12678,4);
TASK_PP(16'h12679,4);
TASK_PP(16'h1267A,4);
TASK_PP(16'h1267B,4);
TASK_PP(16'h1267C,4);
TASK_PP(16'h1267D,4);
TASK_PP(16'h1267E,4);
TASK_PP(16'h1267F,4);
TASK_PP(16'h12680,4);
TASK_PP(16'h12681,4);
TASK_PP(16'h12682,4);
TASK_PP(16'h12683,4);
TASK_PP(16'h12684,4);
TASK_PP(16'h12685,4);
TASK_PP(16'h12686,4);
TASK_PP(16'h12687,4);
TASK_PP(16'h12688,4);
TASK_PP(16'h12689,4);
TASK_PP(16'h1268A,4);
TASK_PP(16'h1268B,4);
TASK_PP(16'h1268C,4);
TASK_PP(16'h1268D,4);
TASK_PP(16'h1268E,4);
TASK_PP(16'h1268F,4);
TASK_PP(16'h12690,4);
TASK_PP(16'h12691,4);
TASK_PP(16'h12692,4);
TASK_PP(16'h12693,4);
TASK_PP(16'h12694,4);
TASK_PP(16'h12695,4);
TASK_PP(16'h12696,4);
TASK_PP(16'h12697,4);
TASK_PP(16'h12698,4);
TASK_PP(16'h12699,4);
TASK_PP(16'h1269A,4);
TASK_PP(16'h1269B,4);
TASK_PP(16'h1269C,4);
TASK_PP(16'h1269D,4);
TASK_PP(16'h1269E,4);
TASK_PP(16'h1269F,4);
TASK_PP(16'h126A0,4);
TASK_PP(16'h126A1,4);
TASK_PP(16'h126A2,4);
TASK_PP(16'h126A3,4);
TASK_PP(16'h126A4,4);
TASK_PP(16'h126A5,4);
TASK_PP(16'h126A6,4);
TASK_PP(16'h126A7,4);
TASK_PP(16'h126A8,4);
TASK_PP(16'h126A9,4);
TASK_PP(16'h126AA,4);
TASK_PP(16'h126AB,4);
TASK_PP(16'h126AC,4);
TASK_PP(16'h126AD,4);
TASK_PP(16'h126AE,4);
TASK_PP(16'h126AF,4);
TASK_PP(16'h126B0,4);
TASK_PP(16'h126B1,4);
TASK_PP(16'h126B2,4);
TASK_PP(16'h126B3,4);
TASK_PP(16'h126B4,4);
TASK_PP(16'h126B5,4);
TASK_PP(16'h126B6,4);
TASK_PP(16'h126B7,4);
TASK_PP(16'h126B8,4);
TASK_PP(16'h126B9,4);
TASK_PP(16'h126BA,4);
TASK_PP(16'h126BB,4);
TASK_PP(16'h126BC,4);
TASK_PP(16'h126BD,4);
TASK_PP(16'h126BE,4);
TASK_PP(16'h126BF,4);
TASK_PP(16'h126C0,4);
TASK_PP(16'h126C1,4);
TASK_PP(16'h126C2,4);
TASK_PP(16'h126C3,4);
TASK_PP(16'h126C4,4);
TASK_PP(16'h126C5,4);
TASK_PP(16'h126C6,4);
TASK_PP(16'h126C7,4);
TASK_PP(16'h126C8,4);
TASK_PP(16'h126C9,4);
TASK_PP(16'h126CA,4);
TASK_PP(16'h126CB,4);
TASK_PP(16'h126CC,4);
TASK_PP(16'h126CD,4);
TASK_PP(16'h126CE,4);
TASK_PP(16'h126CF,4);
TASK_PP(16'h126D0,4);
TASK_PP(16'h126D1,4);
TASK_PP(16'h126D2,4);
TASK_PP(16'h126D3,4);
TASK_PP(16'h126D4,4);
TASK_PP(16'h126D5,4);
TASK_PP(16'h126D6,4);
TASK_PP(16'h126D7,4);
TASK_PP(16'h126D8,4);
TASK_PP(16'h126D9,4);
TASK_PP(16'h126DA,4);
TASK_PP(16'h126DB,4);
TASK_PP(16'h126DC,4);
TASK_PP(16'h126DD,4);
TASK_PP(16'h126DE,4);
TASK_PP(16'h126DF,4);
TASK_PP(16'h126E0,4);
TASK_PP(16'h126E1,4);
TASK_PP(16'h126E2,4);
TASK_PP(16'h126E3,4);
TASK_PP(16'h126E4,4);
TASK_PP(16'h126E5,4);
TASK_PP(16'h126E6,4);
TASK_PP(16'h126E7,4);
TASK_PP(16'h126E8,4);
TASK_PP(16'h126E9,4);
TASK_PP(16'h126EA,4);
TASK_PP(16'h126EB,4);
TASK_PP(16'h126EC,4);
TASK_PP(16'h126ED,4);
TASK_PP(16'h126EE,4);
TASK_PP(16'h126EF,4);
TASK_PP(16'h126F0,4);
TASK_PP(16'h126F1,4);
TASK_PP(16'h126F2,4);
TASK_PP(16'h126F3,4);
TASK_PP(16'h126F4,4);
TASK_PP(16'h126F5,4);
TASK_PP(16'h126F6,4);
TASK_PP(16'h126F7,4);
TASK_PP(16'h126F8,4);
TASK_PP(16'h126F9,4);
TASK_PP(16'h126FA,4);
TASK_PP(16'h126FB,4);
TASK_PP(16'h126FC,4);
TASK_PP(16'h126FD,4);
TASK_PP(16'h126FE,4);
TASK_PP(16'h126FF,4);
TASK_PP(16'h12700,4);
TASK_PP(16'h12701,4);
TASK_PP(16'h12702,4);
TASK_PP(16'h12703,4);
TASK_PP(16'h12704,4);
TASK_PP(16'h12705,4);
TASK_PP(16'h12706,4);
TASK_PP(16'h12707,4);
TASK_PP(16'h12708,4);
TASK_PP(16'h12709,4);
TASK_PP(16'h1270A,4);
TASK_PP(16'h1270B,4);
TASK_PP(16'h1270C,4);
TASK_PP(16'h1270D,4);
TASK_PP(16'h1270E,4);
TASK_PP(16'h1270F,4);
TASK_PP(16'h12710,4);
TASK_PP(16'h12711,4);
TASK_PP(16'h12712,4);
TASK_PP(16'h12713,4);
TASK_PP(16'h12714,4);
TASK_PP(16'h12715,4);
TASK_PP(16'h12716,4);
TASK_PP(16'h12717,4);
TASK_PP(16'h12718,4);
TASK_PP(16'h12719,4);
TASK_PP(16'h1271A,4);
TASK_PP(16'h1271B,4);
TASK_PP(16'h1271C,4);
TASK_PP(16'h1271D,4);
TASK_PP(16'h1271E,4);
TASK_PP(16'h1271F,4);
TASK_PP(16'h12720,4);
TASK_PP(16'h12721,4);
TASK_PP(16'h12722,4);
TASK_PP(16'h12723,4);
TASK_PP(16'h12724,4);
TASK_PP(16'h12725,4);
TASK_PP(16'h12726,4);
TASK_PP(16'h12727,4);
TASK_PP(16'h12728,4);
TASK_PP(16'h12729,4);
TASK_PP(16'h1272A,4);
TASK_PP(16'h1272B,4);
TASK_PP(16'h1272C,4);
TASK_PP(16'h1272D,4);
TASK_PP(16'h1272E,4);
TASK_PP(16'h1272F,4);
TASK_PP(16'h12730,4);
TASK_PP(16'h12731,4);
TASK_PP(16'h12732,4);
TASK_PP(16'h12733,4);
TASK_PP(16'h12734,4);
TASK_PP(16'h12735,4);
TASK_PP(16'h12736,4);
TASK_PP(16'h12737,4);
TASK_PP(16'h12738,4);
TASK_PP(16'h12739,4);
TASK_PP(16'h1273A,4);
TASK_PP(16'h1273B,4);
TASK_PP(16'h1273C,4);
TASK_PP(16'h1273D,4);
TASK_PP(16'h1273E,4);
TASK_PP(16'h1273F,4);
TASK_PP(16'h12740,4);
TASK_PP(16'h12741,4);
TASK_PP(16'h12742,4);
TASK_PP(16'h12743,4);
TASK_PP(16'h12744,4);
TASK_PP(16'h12745,4);
TASK_PP(16'h12746,4);
TASK_PP(16'h12747,4);
TASK_PP(16'h12748,4);
TASK_PP(16'h12749,4);
TASK_PP(16'h1274A,4);
TASK_PP(16'h1274B,4);
TASK_PP(16'h1274C,4);
TASK_PP(16'h1274D,4);
TASK_PP(16'h1274E,4);
TASK_PP(16'h1274F,4);
TASK_PP(16'h12750,4);
TASK_PP(16'h12751,4);
TASK_PP(16'h12752,4);
TASK_PP(16'h12753,4);
TASK_PP(16'h12754,4);
TASK_PP(16'h12755,4);
TASK_PP(16'h12756,4);
TASK_PP(16'h12757,4);
TASK_PP(16'h12758,4);
TASK_PP(16'h12759,4);
TASK_PP(16'h1275A,4);
TASK_PP(16'h1275B,4);
TASK_PP(16'h1275C,4);
TASK_PP(16'h1275D,4);
TASK_PP(16'h1275E,4);
TASK_PP(16'h1275F,4);
TASK_PP(16'h12760,4);
TASK_PP(16'h12761,4);
TASK_PP(16'h12762,4);
TASK_PP(16'h12763,4);
TASK_PP(16'h12764,4);
TASK_PP(16'h12765,4);
TASK_PP(16'h12766,4);
TASK_PP(16'h12767,4);
TASK_PP(16'h12768,4);
TASK_PP(16'h12769,4);
TASK_PP(16'h1276A,4);
TASK_PP(16'h1276B,4);
TASK_PP(16'h1276C,4);
TASK_PP(16'h1276D,4);
TASK_PP(16'h1276E,4);
TASK_PP(16'h1276F,4);
TASK_PP(16'h12770,4);
TASK_PP(16'h12771,4);
TASK_PP(16'h12772,4);
TASK_PP(16'h12773,4);
TASK_PP(16'h12774,4);
TASK_PP(16'h12775,4);
TASK_PP(16'h12776,4);
TASK_PP(16'h12777,4);
TASK_PP(16'h12778,4);
TASK_PP(16'h12779,4);
TASK_PP(16'h1277A,4);
TASK_PP(16'h1277B,4);
TASK_PP(16'h1277C,4);
TASK_PP(16'h1277D,4);
TASK_PP(16'h1277E,4);
TASK_PP(16'h1277F,4);
TASK_PP(16'h12780,4);
TASK_PP(16'h12781,4);
TASK_PP(16'h12782,4);
TASK_PP(16'h12783,4);
TASK_PP(16'h12784,4);
TASK_PP(16'h12785,4);
TASK_PP(16'h12786,4);
TASK_PP(16'h12787,4);
TASK_PP(16'h12788,4);
TASK_PP(16'h12789,4);
TASK_PP(16'h1278A,4);
TASK_PP(16'h1278B,4);
TASK_PP(16'h1278C,4);
TASK_PP(16'h1278D,4);
TASK_PP(16'h1278E,4);
TASK_PP(16'h1278F,4);
TASK_PP(16'h12790,4);
TASK_PP(16'h12791,4);
TASK_PP(16'h12792,4);
TASK_PP(16'h12793,4);
TASK_PP(16'h12794,4);
TASK_PP(16'h12795,4);
TASK_PP(16'h12796,4);
TASK_PP(16'h12797,4);
TASK_PP(16'h12798,4);
TASK_PP(16'h12799,4);
TASK_PP(16'h1279A,4);
TASK_PP(16'h1279B,4);
TASK_PP(16'h1279C,4);
TASK_PP(16'h1279D,4);
TASK_PP(16'h1279E,4);
TASK_PP(16'h1279F,4);
TASK_PP(16'h127A0,4);
TASK_PP(16'h127A1,4);
TASK_PP(16'h127A2,4);
TASK_PP(16'h127A3,4);
TASK_PP(16'h127A4,4);
TASK_PP(16'h127A5,4);
TASK_PP(16'h127A6,4);
TASK_PP(16'h127A7,4);
TASK_PP(16'h127A8,4);
TASK_PP(16'h127A9,4);
TASK_PP(16'h127AA,4);
TASK_PP(16'h127AB,4);
TASK_PP(16'h127AC,4);
TASK_PP(16'h127AD,4);
TASK_PP(16'h127AE,4);
TASK_PP(16'h127AF,4);
TASK_PP(16'h127B0,4);
TASK_PP(16'h127B1,4);
TASK_PP(16'h127B2,4);
TASK_PP(16'h127B3,4);
TASK_PP(16'h127B4,4);
TASK_PP(16'h127B5,4);
TASK_PP(16'h127B6,4);
TASK_PP(16'h127B7,4);
TASK_PP(16'h127B8,4);
TASK_PP(16'h127B9,4);
TASK_PP(16'h127BA,4);
TASK_PP(16'h127BB,4);
TASK_PP(16'h127BC,4);
TASK_PP(16'h127BD,4);
TASK_PP(16'h127BE,4);
TASK_PP(16'h127BF,4);
TASK_PP(16'h127C0,4);
TASK_PP(16'h127C1,4);
TASK_PP(16'h127C2,4);
TASK_PP(16'h127C3,4);
TASK_PP(16'h127C4,4);
TASK_PP(16'h127C5,4);
TASK_PP(16'h127C6,4);
TASK_PP(16'h127C7,4);
TASK_PP(16'h127C8,4);
TASK_PP(16'h127C9,4);
TASK_PP(16'h127CA,4);
TASK_PP(16'h127CB,4);
TASK_PP(16'h127CC,4);
TASK_PP(16'h127CD,4);
TASK_PP(16'h127CE,4);
TASK_PP(16'h127CF,4);
TASK_PP(16'h127D0,4);
TASK_PP(16'h127D1,4);
TASK_PP(16'h127D2,4);
TASK_PP(16'h127D3,4);
TASK_PP(16'h127D4,4);
TASK_PP(16'h127D5,4);
TASK_PP(16'h127D6,4);
TASK_PP(16'h127D7,4);
TASK_PP(16'h127D8,4);
TASK_PP(16'h127D9,4);
TASK_PP(16'h127DA,4);
TASK_PP(16'h127DB,4);
TASK_PP(16'h127DC,4);
TASK_PP(16'h127DD,4);
TASK_PP(16'h127DE,4);
TASK_PP(16'h127DF,4);
TASK_PP(16'h127E0,4);
TASK_PP(16'h127E1,4);
TASK_PP(16'h127E2,4);
TASK_PP(16'h127E3,4);
TASK_PP(16'h127E4,4);
TASK_PP(16'h127E5,4);
TASK_PP(16'h127E6,4);
TASK_PP(16'h127E7,4);
TASK_PP(16'h127E8,4);
TASK_PP(16'h127E9,4);
TASK_PP(16'h127EA,4);
TASK_PP(16'h127EB,4);
TASK_PP(16'h127EC,4);
TASK_PP(16'h127ED,4);
TASK_PP(16'h127EE,4);
TASK_PP(16'h127EF,4);
TASK_PP(16'h127F0,4);
TASK_PP(16'h127F1,4);
TASK_PP(16'h127F2,4);
TASK_PP(16'h127F3,4);
TASK_PP(16'h127F4,4);
TASK_PP(16'h127F5,4);
TASK_PP(16'h127F6,4);
TASK_PP(16'h127F7,4);
TASK_PP(16'h127F8,4);
TASK_PP(16'h127F9,4);
TASK_PP(16'h127FA,4);
TASK_PP(16'h127FB,4);
TASK_PP(16'h127FC,4);
TASK_PP(16'h127FD,4);
TASK_PP(16'h127FE,4);
TASK_PP(16'h127FF,4);
TASK_PP(16'h12800,4);
TASK_PP(16'h12801,4);
TASK_PP(16'h12802,4);
TASK_PP(16'h12803,4);
TASK_PP(16'h12804,4);
TASK_PP(16'h12805,4);
TASK_PP(16'h12806,4);
TASK_PP(16'h12807,4);
TASK_PP(16'h12808,4);
TASK_PP(16'h12809,4);
TASK_PP(16'h1280A,4);
TASK_PP(16'h1280B,4);
TASK_PP(16'h1280C,4);
TASK_PP(16'h1280D,4);
TASK_PP(16'h1280E,4);
TASK_PP(16'h1280F,4);
TASK_PP(16'h12810,4);
TASK_PP(16'h12811,4);
TASK_PP(16'h12812,4);
TASK_PP(16'h12813,4);
TASK_PP(16'h12814,4);
TASK_PP(16'h12815,4);
TASK_PP(16'h12816,4);
TASK_PP(16'h12817,4);
TASK_PP(16'h12818,4);
TASK_PP(16'h12819,4);
TASK_PP(16'h1281A,4);
TASK_PP(16'h1281B,4);
TASK_PP(16'h1281C,4);
TASK_PP(16'h1281D,4);
TASK_PP(16'h1281E,4);
TASK_PP(16'h1281F,4);
TASK_PP(16'h12820,4);
TASK_PP(16'h12821,4);
TASK_PP(16'h12822,4);
TASK_PP(16'h12823,4);
TASK_PP(16'h12824,4);
TASK_PP(16'h12825,4);
TASK_PP(16'h12826,4);
TASK_PP(16'h12827,4);
TASK_PP(16'h12828,4);
TASK_PP(16'h12829,4);
TASK_PP(16'h1282A,4);
TASK_PP(16'h1282B,4);
TASK_PP(16'h1282C,4);
TASK_PP(16'h1282D,4);
TASK_PP(16'h1282E,4);
TASK_PP(16'h1282F,4);
TASK_PP(16'h12830,4);
TASK_PP(16'h12831,4);
TASK_PP(16'h12832,4);
TASK_PP(16'h12833,4);
TASK_PP(16'h12834,4);
TASK_PP(16'h12835,4);
TASK_PP(16'h12836,4);
TASK_PP(16'h12837,4);
TASK_PP(16'h12838,4);
TASK_PP(16'h12839,4);
TASK_PP(16'h1283A,4);
TASK_PP(16'h1283B,4);
TASK_PP(16'h1283C,4);
TASK_PP(16'h1283D,4);
TASK_PP(16'h1283E,4);
TASK_PP(16'h1283F,4);
TASK_PP(16'h12840,4);
TASK_PP(16'h12841,4);
TASK_PP(16'h12842,4);
TASK_PP(16'h12843,4);
TASK_PP(16'h12844,4);
TASK_PP(16'h12845,4);
TASK_PP(16'h12846,4);
TASK_PP(16'h12847,4);
TASK_PP(16'h12848,4);
TASK_PP(16'h12849,4);
TASK_PP(16'h1284A,4);
TASK_PP(16'h1284B,4);
TASK_PP(16'h1284C,4);
TASK_PP(16'h1284D,4);
TASK_PP(16'h1284E,4);
TASK_PP(16'h1284F,4);
TASK_PP(16'h12850,4);
TASK_PP(16'h12851,4);
TASK_PP(16'h12852,4);
TASK_PP(16'h12853,4);
TASK_PP(16'h12854,4);
TASK_PP(16'h12855,4);
TASK_PP(16'h12856,4);
TASK_PP(16'h12857,4);
TASK_PP(16'h12858,4);
TASK_PP(16'h12859,4);
TASK_PP(16'h1285A,4);
TASK_PP(16'h1285B,4);
TASK_PP(16'h1285C,4);
TASK_PP(16'h1285D,4);
TASK_PP(16'h1285E,4);
TASK_PP(16'h1285F,4);
TASK_PP(16'h12860,4);
TASK_PP(16'h12861,4);
TASK_PP(16'h12862,4);
TASK_PP(16'h12863,4);
TASK_PP(16'h12864,4);
TASK_PP(16'h12865,4);
TASK_PP(16'h12866,4);
TASK_PP(16'h12867,4);
TASK_PP(16'h12868,4);
TASK_PP(16'h12869,4);
TASK_PP(16'h1286A,4);
TASK_PP(16'h1286B,4);
TASK_PP(16'h1286C,4);
TASK_PP(16'h1286D,4);
TASK_PP(16'h1286E,4);
TASK_PP(16'h1286F,4);
TASK_PP(16'h12870,4);
TASK_PP(16'h12871,4);
TASK_PP(16'h12872,4);
TASK_PP(16'h12873,4);
TASK_PP(16'h12874,4);
TASK_PP(16'h12875,4);
TASK_PP(16'h12876,4);
TASK_PP(16'h12877,4);
TASK_PP(16'h12878,4);
TASK_PP(16'h12879,4);
TASK_PP(16'h1287A,4);
TASK_PP(16'h1287B,4);
TASK_PP(16'h1287C,4);
TASK_PP(16'h1287D,4);
TASK_PP(16'h1287E,4);
TASK_PP(16'h1287F,4);
TASK_PP(16'h12880,4);
TASK_PP(16'h12881,4);
TASK_PP(16'h12882,4);
TASK_PP(16'h12883,4);
TASK_PP(16'h12884,4);
TASK_PP(16'h12885,4);
TASK_PP(16'h12886,4);
TASK_PP(16'h12887,4);
TASK_PP(16'h12888,4);
TASK_PP(16'h12889,4);
TASK_PP(16'h1288A,4);
TASK_PP(16'h1288B,4);
TASK_PP(16'h1288C,4);
TASK_PP(16'h1288D,4);
TASK_PP(16'h1288E,4);
TASK_PP(16'h1288F,4);
TASK_PP(16'h12890,4);
TASK_PP(16'h12891,4);
TASK_PP(16'h12892,4);
TASK_PP(16'h12893,4);
TASK_PP(16'h12894,4);
TASK_PP(16'h12895,4);
TASK_PP(16'h12896,4);
TASK_PP(16'h12897,4);
TASK_PP(16'h12898,4);
TASK_PP(16'h12899,4);
TASK_PP(16'h1289A,4);
TASK_PP(16'h1289B,4);
TASK_PP(16'h1289C,4);
TASK_PP(16'h1289D,4);
TASK_PP(16'h1289E,4);
TASK_PP(16'h1289F,4);
TASK_PP(16'h128A0,4);
TASK_PP(16'h128A1,4);
TASK_PP(16'h128A2,4);
TASK_PP(16'h128A3,4);
TASK_PP(16'h128A4,4);
TASK_PP(16'h128A5,4);
TASK_PP(16'h128A6,4);
TASK_PP(16'h128A7,4);
TASK_PP(16'h128A8,4);
TASK_PP(16'h128A9,4);
TASK_PP(16'h128AA,4);
TASK_PP(16'h128AB,4);
TASK_PP(16'h128AC,4);
TASK_PP(16'h128AD,4);
TASK_PP(16'h128AE,4);
TASK_PP(16'h128AF,4);
TASK_PP(16'h128B0,4);
TASK_PP(16'h128B1,4);
TASK_PP(16'h128B2,4);
TASK_PP(16'h128B3,4);
TASK_PP(16'h128B4,4);
TASK_PP(16'h128B5,4);
TASK_PP(16'h128B6,4);
TASK_PP(16'h128B7,4);
TASK_PP(16'h128B8,4);
TASK_PP(16'h128B9,4);
TASK_PP(16'h128BA,4);
TASK_PP(16'h128BB,4);
TASK_PP(16'h128BC,4);
TASK_PP(16'h128BD,4);
TASK_PP(16'h128BE,4);
TASK_PP(16'h128BF,4);
TASK_PP(16'h128C0,4);
TASK_PP(16'h128C1,4);
TASK_PP(16'h128C2,4);
TASK_PP(16'h128C3,4);
TASK_PP(16'h128C4,4);
TASK_PP(16'h128C5,4);
TASK_PP(16'h128C6,4);
TASK_PP(16'h128C7,4);
TASK_PP(16'h128C8,4);
TASK_PP(16'h128C9,4);
TASK_PP(16'h128CA,4);
TASK_PP(16'h128CB,4);
TASK_PP(16'h128CC,4);
TASK_PP(16'h128CD,4);
TASK_PP(16'h128CE,4);
TASK_PP(16'h128CF,4);
TASK_PP(16'h128D0,4);
TASK_PP(16'h128D1,4);
TASK_PP(16'h128D2,4);
TASK_PP(16'h128D3,4);
TASK_PP(16'h128D4,4);
TASK_PP(16'h128D5,4);
TASK_PP(16'h128D6,4);
TASK_PP(16'h128D7,4);
TASK_PP(16'h128D8,4);
TASK_PP(16'h128D9,4);
TASK_PP(16'h128DA,4);
TASK_PP(16'h128DB,4);
TASK_PP(16'h128DC,4);
TASK_PP(16'h128DD,4);
TASK_PP(16'h128DE,4);
TASK_PP(16'h128DF,4);
TASK_PP(16'h128E0,4);
TASK_PP(16'h128E1,4);
TASK_PP(16'h128E2,4);
TASK_PP(16'h128E3,4);
TASK_PP(16'h128E4,4);
TASK_PP(16'h128E5,4);
TASK_PP(16'h128E6,4);
TASK_PP(16'h128E7,4);
TASK_PP(16'h128E8,4);
TASK_PP(16'h128E9,4);
TASK_PP(16'h128EA,4);
TASK_PP(16'h128EB,4);
TASK_PP(16'h128EC,4);
TASK_PP(16'h128ED,4);
TASK_PP(16'h128EE,4);
TASK_PP(16'h128EF,4);
TASK_PP(16'h128F0,4);
TASK_PP(16'h128F1,4);
TASK_PP(16'h128F2,4);
TASK_PP(16'h128F3,4);
TASK_PP(16'h128F4,4);
TASK_PP(16'h128F5,4);
TASK_PP(16'h128F6,4);
TASK_PP(16'h128F7,4);
TASK_PP(16'h128F8,4);
TASK_PP(16'h128F9,4);
TASK_PP(16'h128FA,4);
TASK_PP(16'h128FB,4);
TASK_PP(16'h128FC,4);
TASK_PP(16'h128FD,4);
TASK_PP(16'h128FE,4);
TASK_PP(16'h128FF,4);
TASK_PP(16'h12900,4);
TASK_PP(16'h12901,4);
TASK_PP(16'h12902,4);
TASK_PP(16'h12903,4);
TASK_PP(16'h12904,4);
TASK_PP(16'h12905,4);
TASK_PP(16'h12906,4);
TASK_PP(16'h12907,4);
TASK_PP(16'h12908,4);
TASK_PP(16'h12909,4);
TASK_PP(16'h1290A,4);
TASK_PP(16'h1290B,4);
TASK_PP(16'h1290C,4);
TASK_PP(16'h1290D,4);
TASK_PP(16'h1290E,4);
TASK_PP(16'h1290F,4);
TASK_PP(16'h12910,4);
TASK_PP(16'h12911,4);
TASK_PP(16'h12912,4);
TASK_PP(16'h12913,4);
TASK_PP(16'h12914,4);
TASK_PP(16'h12915,4);
TASK_PP(16'h12916,4);
TASK_PP(16'h12917,4);
TASK_PP(16'h12918,4);
TASK_PP(16'h12919,4);
TASK_PP(16'h1291A,4);
TASK_PP(16'h1291B,4);
TASK_PP(16'h1291C,4);
TASK_PP(16'h1291D,4);
TASK_PP(16'h1291E,4);
TASK_PP(16'h1291F,4);
TASK_PP(16'h12920,4);
TASK_PP(16'h12921,4);
TASK_PP(16'h12922,4);
TASK_PP(16'h12923,4);
TASK_PP(16'h12924,4);
TASK_PP(16'h12925,4);
TASK_PP(16'h12926,4);
TASK_PP(16'h12927,4);
TASK_PP(16'h12928,4);
TASK_PP(16'h12929,4);
TASK_PP(16'h1292A,4);
TASK_PP(16'h1292B,4);
TASK_PP(16'h1292C,4);
TASK_PP(16'h1292D,4);
TASK_PP(16'h1292E,4);
TASK_PP(16'h1292F,4);
TASK_PP(16'h12930,4);
TASK_PP(16'h12931,4);
TASK_PP(16'h12932,4);
TASK_PP(16'h12933,4);
TASK_PP(16'h12934,4);
TASK_PP(16'h12935,4);
TASK_PP(16'h12936,4);
TASK_PP(16'h12937,4);
TASK_PP(16'h12938,4);
TASK_PP(16'h12939,4);
TASK_PP(16'h1293A,4);
TASK_PP(16'h1293B,4);
TASK_PP(16'h1293C,4);
TASK_PP(16'h1293D,4);
TASK_PP(16'h1293E,4);
TASK_PP(16'h1293F,4);
TASK_PP(16'h12940,4);
TASK_PP(16'h12941,4);
TASK_PP(16'h12942,4);
TASK_PP(16'h12943,4);
TASK_PP(16'h12944,4);
TASK_PP(16'h12945,4);
TASK_PP(16'h12946,4);
TASK_PP(16'h12947,4);
TASK_PP(16'h12948,4);
TASK_PP(16'h12949,4);
TASK_PP(16'h1294A,4);
TASK_PP(16'h1294B,4);
TASK_PP(16'h1294C,4);
TASK_PP(16'h1294D,4);
TASK_PP(16'h1294E,4);
TASK_PP(16'h1294F,4);
TASK_PP(16'h12950,4);
TASK_PP(16'h12951,4);
TASK_PP(16'h12952,4);
TASK_PP(16'h12953,4);
TASK_PP(16'h12954,4);
TASK_PP(16'h12955,4);
TASK_PP(16'h12956,4);
TASK_PP(16'h12957,4);
TASK_PP(16'h12958,4);
TASK_PP(16'h12959,4);
TASK_PP(16'h1295A,4);
TASK_PP(16'h1295B,4);
TASK_PP(16'h1295C,4);
TASK_PP(16'h1295D,4);
TASK_PP(16'h1295E,4);
TASK_PP(16'h1295F,4);
TASK_PP(16'h12960,4);
TASK_PP(16'h12961,4);
TASK_PP(16'h12962,4);
TASK_PP(16'h12963,4);
TASK_PP(16'h12964,4);
TASK_PP(16'h12965,4);
TASK_PP(16'h12966,4);
TASK_PP(16'h12967,4);
TASK_PP(16'h12968,4);
TASK_PP(16'h12969,4);
TASK_PP(16'h1296A,4);
TASK_PP(16'h1296B,4);
TASK_PP(16'h1296C,4);
TASK_PP(16'h1296D,4);
TASK_PP(16'h1296E,4);
TASK_PP(16'h1296F,4);
TASK_PP(16'h12970,4);
TASK_PP(16'h12971,4);
TASK_PP(16'h12972,4);
TASK_PP(16'h12973,4);
TASK_PP(16'h12974,4);
TASK_PP(16'h12975,4);
TASK_PP(16'h12976,4);
TASK_PP(16'h12977,4);
TASK_PP(16'h12978,4);
TASK_PP(16'h12979,4);
TASK_PP(16'h1297A,4);
TASK_PP(16'h1297B,4);
TASK_PP(16'h1297C,4);
TASK_PP(16'h1297D,4);
TASK_PP(16'h1297E,4);
TASK_PP(16'h1297F,4);
TASK_PP(16'h12980,4);
TASK_PP(16'h12981,4);
TASK_PP(16'h12982,4);
TASK_PP(16'h12983,4);
TASK_PP(16'h12984,4);
TASK_PP(16'h12985,4);
TASK_PP(16'h12986,4);
TASK_PP(16'h12987,4);
TASK_PP(16'h12988,4);
TASK_PP(16'h12989,4);
TASK_PP(16'h1298A,4);
TASK_PP(16'h1298B,4);
TASK_PP(16'h1298C,4);
TASK_PP(16'h1298D,4);
TASK_PP(16'h1298E,4);
TASK_PP(16'h1298F,4);
TASK_PP(16'h12990,4);
TASK_PP(16'h12991,4);
TASK_PP(16'h12992,4);
TASK_PP(16'h12993,4);
TASK_PP(16'h12994,4);
TASK_PP(16'h12995,4);
TASK_PP(16'h12996,4);
TASK_PP(16'h12997,4);
TASK_PP(16'h12998,4);
TASK_PP(16'h12999,4);
TASK_PP(16'h1299A,4);
TASK_PP(16'h1299B,4);
TASK_PP(16'h1299C,4);
TASK_PP(16'h1299D,4);
TASK_PP(16'h1299E,4);
TASK_PP(16'h1299F,4);
TASK_PP(16'h129A0,4);
TASK_PP(16'h129A1,4);
TASK_PP(16'h129A2,4);
TASK_PP(16'h129A3,4);
TASK_PP(16'h129A4,4);
TASK_PP(16'h129A5,4);
TASK_PP(16'h129A6,4);
TASK_PP(16'h129A7,4);
TASK_PP(16'h129A8,4);
TASK_PP(16'h129A9,4);
TASK_PP(16'h129AA,4);
TASK_PP(16'h129AB,4);
TASK_PP(16'h129AC,4);
TASK_PP(16'h129AD,4);
TASK_PP(16'h129AE,4);
TASK_PP(16'h129AF,4);
TASK_PP(16'h129B0,4);
TASK_PP(16'h129B1,4);
TASK_PP(16'h129B2,4);
TASK_PP(16'h129B3,4);
TASK_PP(16'h129B4,4);
TASK_PP(16'h129B5,4);
TASK_PP(16'h129B6,4);
TASK_PP(16'h129B7,4);
TASK_PP(16'h129B8,4);
TASK_PP(16'h129B9,4);
TASK_PP(16'h129BA,4);
TASK_PP(16'h129BB,4);
TASK_PP(16'h129BC,4);
TASK_PP(16'h129BD,4);
TASK_PP(16'h129BE,4);
TASK_PP(16'h129BF,4);
TASK_PP(16'h129C0,4);
TASK_PP(16'h129C1,4);
TASK_PP(16'h129C2,4);
TASK_PP(16'h129C3,4);
TASK_PP(16'h129C4,4);
TASK_PP(16'h129C5,4);
TASK_PP(16'h129C6,4);
TASK_PP(16'h129C7,4);
TASK_PP(16'h129C8,4);
TASK_PP(16'h129C9,4);
TASK_PP(16'h129CA,4);
TASK_PP(16'h129CB,4);
TASK_PP(16'h129CC,4);
TASK_PP(16'h129CD,4);
TASK_PP(16'h129CE,4);
TASK_PP(16'h129CF,4);
TASK_PP(16'h129D0,4);
TASK_PP(16'h129D1,4);
TASK_PP(16'h129D2,4);
TASK_PP(16'h129D3,4);
TASK_PP(16'h129D4,4);
TASK_PP(16'h129D5,4);
TASK_PP(16'h129D6,4);
TASK_PP(16'h129D7,4);
TASK_PP(16'h129D8,4);
TASK_PP(16'h129D9,4);
TASK_PP(16'h129DA,4);
TASK_PP(16'h129DB,4);
TASK_PP(16'h129DC,4);
TASK_PP(16'h129DD,4);
TASK_PP(16'h129DE,4);
TASK_PP(16'h129DF,4);
TASK_PP(16'h129E0,4);
TASK_PP(16'h129E1,4);
TASK_PP(16'h129E2,4);
TASK_PP(16'h129E3,4);
TASK_PP(16'h129E4,4);
TASK_PP(16'h129E5,4);
TASK_PP(16'h129E6,4);
TASK_PP(16'h129E7,4);
TASK_PP(16'h129E8,4);
TASK_PP(16'h129E9,4);
TASK_PP(16'h129EA,4);
TASK_PP(16'h129EB,4);
TASK_PP(16'h129EC,4);
TASK_PP(16'h129ED,4);
TASK_PP(16'h129EE,4);
TASK_PP(16'h129EF,4);
TASK_PP(16'h129F0,4);
TASK_PP(16'h129F1,4);
TASK_PP(16'h129F2,4);
TASK_PP(16'h129F3,4);
TASK_PP(16'h129F4,4);
TASK_PP(16'h129F5,4);
TASK_PP(16'h129F6,4);
TASK_PP(16'h129F7,4);
TASK_PP(16'h129F8,4);
TASK_PP(16'h129F9,4);
TASK_PP(16'h129FA,4);
TASK_PP(16'h129FB,4);
TASK_PP(16'h129FC,4);
TASK_PP(16'h129FD,4);
TASK_PP(16'h129FE,4);
TASK_PP(16'h129FF,4);
TASK_PP(16'h12A00,4);
TASK_PP(16'h12A01,4);
TASK_PP(16'h12A02,4);
TASK_PP(16'h12A03,4);
TASK_PP(16'h12A04,4);
TASK_PP(16'h12A05,4);
TASK_PP(16'h12A06,4);
TASK_PP(16'h12A07,4);
TASK_PP(16'h12A08,4);
TASK_PP(16'h12A09,4);
TASK_PP(16'h12A0A,4);
TASK_PP(16'h12A0B,4);
TASK_PP(16'h12A0C,4);
TASK_PP(16'h12A0D,4);
TASK_PP(16'h12A0E,4);
TASK_PP(16'h12A0F,4);
TASK_PP(16'h12A10,4);
TASK_PP(16'h12A11,4);
TASK_PP(16'h12A12,4);
TASK_PP(16'h12A13,4);
TASK_PP(16'h12A14,4);
TASK_PP(16'h12A15,4);
TASK_PP(16'h12A16,4);
TASK_PP(16'h12A17,4);
TASK_PP(16'h12A18,4);
TASK_PP(16'h12A19,4);
TASK_PP(16'h12A1A,4);
TASK_PP(16'h12A1B,4);
TASK_PP(16'h12A1C,4);
TASK_PP(16'h12A1D,4);
TASK_PP(16'h12A1E,4);
TASK_PP(16'h12A1F,4);
TASK_PP(16'h12A20,4);
TASK_PP(16'h12A21,4);
TASK_PP(16'h12A22,4);
TASK_PP(16'h12A23,4);
TASK_PP(16'h12A24,4);
TASK_PP(16'h12A25,4);
TASK_PP(16'h12A26,4);
TASK_PP(16'h12A27,4);
TASK_PP(16'h12A28,4);
TASK_PP(16'h12A29,4);
TASK_PP(16'h12A2A,4);
TASK_PP(16'h12A2B,4);
TASK_PP(16'h12A2C,4);
TASK_PP(16'h12A2D,4);
TASK_PP(16'h12A2E,4);
TASK_PP(16'h12A2F,4);
TASK_PP(16'h12A30,4);
TASK_PP(16'h12A31,4);
TASK_PP(16'h12A32,4);
TASK_PP(16'h12A33,4);
TASK_PP(16'h12A34,4);
TASK_PP(16'h12A35,4);
TASK_PP(16'h12A36,4);
TASK_PP(16'h12A37,4);
TASK_PP(16'h12A38,4);
TASK_PP(16'h12A39,4);
TASK_PP(16'h12A3A,4);
TASK_PP(16'h12A3B,4);
TASK_PP(16'h12A3C,4);
TASK_PP(16'h12A3D,4);
TASK_PP(16'h12A3E,4);
TASK_PP(16'h12A3F,4);
TASK_PP(16'h12A40,4);
TASK_PP(16'h12A41,4);
TASK_PP(16'h12A42,4);
TASK_PP(16'h12A43,4);
TASK_PP(16'h12A44,4);
TASK_PP(16'h12A45,4);
TASK_PP(16'h12A46,4);
TASK_PP(16'h12A47,4);
TASK_PP(16'h12A48,4);
TASK_PP(16'h12A49,4);
TASK_PP(16'h12A4A,4);
TASK_PP(16'h12A4B,4);
TASK_PP(16'h12A4C,4);
TASK_PP(16'h12A4D,4);
TASK_PP(16'h12A4E,4);
TASK_PP(16'h12A4F,4);
TASK_PP(16'h12A50,4);
TASK_PP(16'h12A51,4);
TASK_PP(16'h12A52,4);
TASK_PP(16'h12A53,4);
TASK_PP(16'h12A54,4);
TASK_PP(16'h12A55,4);
TASK_PP(16'h12A56,4);
TASK_PP(16'h12A57,4);
TASK_PP(16'h12A58,4);
TASK_PP(16'h12A59,4);
TASK_PP(16'h12A5A,4);
TASK_PP(16'h12A5B,4);
TASK_PP(16'h12A5C,4);
TASK_PP(16'h12A5D,4);
TASK_PP(16'h12A5E,4);
TASK_PP(16'h12A5F,4);
TASK_PP(16'h12A60,4);
TASK_PP(16'h12A61,4);
TASK_PP(16'h12A62,4);
TASK_PP(16'h12A63,4);
TASK_PP(16'h12A64,4);
TASK_PP(16'h12A65,4);
TASK_PP(16'h12A66,4);
TASK_PP(16'h12A67,4);
TASK_PP(16'h12A68,4);
TASK_PP(16'h12A69,4);
TASK_PP(16'h12A6A,4);
TASK_PP(16'h12A6B,4);
TASK_PP(16'h12A6C,4);
TASK_PP(16'h12A6D,4);
TASK_PP(16'h12A6E,4);
TASK_PP(16'h12A6F,4);
TASK_PP(16'h12A70,4);
TASK_PP(16'h12A71,4);
TASK_PP(16'h12A72,4);
TASK_PP(16'h12A73,4);
TASK_PP(16'h12A74,4);
TASK_PP(16'h12A75,4);
TASK_PP(16'h12A76,4);
TASK_PP(16'h12A77,4);
TASK_PP(16'h12A78,4);
TASK_PP(16'h12A79,4);
TASK_PP(16'h12A7A,4);
TASK_PP(16'h12A7B,4);
TASK_PP(16'h12A7C,4);
TASK_PP(16'h12A7D,4);
TASK_PP(16'h12A7E,4);
TASK_PP(16'h12A7F,4);
TASK_PP(16'h12A80,4);
TASK_PP(16'h12A81,4);
TASK_PP(16'h12A82,4);
TASK_PP(16'h12A83,4);
TASK_PP(16'h12A84,4);
TASK_PP(16'h12A85,4);
TASK_PP(16'h12A86,4);
TASK_PP(16'h12A87,4);
TASK_PP(16'h12A88,4);
TASK_PP(16'h12A89,4);
TASK_PP(16'h12A8A,4);
TASK_PP(16'h12A8B,4);
TASK_PP(16'h12A8C,4);
TASK_PP(16'h12A8D,4);
TASK_PP(16'h12A8E,4);
TASK_PP(16'h12A8F,4);
TASK_PP(16'h12A90,4);
TASK_PP(16'h12A91,4);
TASK_PP(16'h12A92,4);
TASK_PP(16'h12A93,4);
TASK_PP(16'h12A94,4);
TASK_PP(16'h12A95,4);
TASK_PP(16'h12A96,4);
TASK_PP(16'h12A97,4);
TASK_PP(16'h12A98,4);
TASK_PP(16'h12A99,4);
TASK_PP(16'h12A9A,4);
TASK_PP(16'h12A9B,4);
TASK_PP(16'h12A9C,4);
TASK_PP(16'h12A9D,4);
TASK_PP(16'h12A9E,4);
TASK_PP(16'h12A9F,4);
TASK_PP(16'h12AA0,4);
TASK_PP(16'h12AA1,4);
TASK_PP(16'h12AA2,4);
TASK_PP(16'h12AA3,4);
TASK_PP(16'h12AA4,4);
TASK_PP(16'h12AA5,4);
TASK_PP(16'h12AA6,4);
TASK_PP(16'h12AA7,4);
TASK_PP(16'h12AA8,4);
TASK_PP(16'h12AA9,4);
TASK_PP(16'h12AAA,4);
TASK_PP(16'h12AAB,4);
TASK_PP(16'h12AAC,4);
TASK_PP(16'h12AAD,4);
TASK_PP(16'h12AAE,4);
TASK_PP(16'h12AAF,4);
TASK_PP(16'h12AB0,4);
TASK_PP(16'h12AB1,4);
TASK_PP(16'h12AB2,4);
TASK_PP(16'h12AB3,4);
TASK_PP(16'h12AB4,4);
TASK_PP(16'h12AB5,4);
TASK_PP(16'h12AB6,4);
TASK_PP(16'h12AB7,4);
TASK_PP(16'h12AB8,4);
TASK_PP(16'h12AB9,4);
TASK_PP(16'h12ABA,4);
TASK_PP(16'h12ABB,4);
TASK_PP(16'h12ABC,4);
TASK_PP(16'h12ABD,4);
TASK_PP(16'h12ABE,4);
TASK_PP(16'h12ABF,4);
TASK_PP(16'h12AC0,4);
TASK_PP(16'h12AC1,4);
TASK_PP(16'h12AC2,4);
TASK_PP(16'h12AC3,4);
TASK_PP(16'h12AC4,4);
TASK_PP(16'h12AC5,4);
TASK_PP(16'h12AC6,4);
TASK_PP(16'h12AC7,4);
TASK_PP(16'h12AC8,4);
TASK_PP(16'h12AC9,4);
TASK_PP(16'h12ACA,4);
TASK_PP(16'h12ACB,4);
TASK_PP(16'h12ACC,4);
TASK_PP(16'h12ACD,4);
TASK_PP(16'h12ACE,4);
TASK_PP(16'h12ACF,4);
TASK_PP(16'h12AD0,4);
TASK_PP(16'h12AD1,4);
TASK_PP(16'h12AD2,4);
TASK_PP(16'h12AD3,4);
TASK_PP(16'h12AD4,4);
TASK_PP(16'h12AD5,4);
TASK_PP(16'h12AD6,4);
TASK_PP(16'h12AD7,4);
TASK_PP(16'h12AD8,4);
TASK_PP(16'h12AD9,4);
TASK_PP(16'h12ADA,4);
TASK_PP(16'h12ADB,4);
TASK_PP(16'h12ADC,4);
TASK_PP(16'h12ADD,4);
TASK_PP(16'h12ADE,4);
TASK_PP(16'h12ADF,4);
TASK_PP(16'h12AE0,4);
TASK_PP(16'h12AE1,4);
TASK_PP(16'h12AE2,4);
TASK_PP(16'h12AE3,4);
TASK_PP(16'h12AE4,4);
TASK_PP(16'h12AE5,4);
TASK_PP(16'h12AE6,4);
TASK_PP(16'h12AE7,4);
TASK_PP(16'h12AE8,4);
TASK_PP(16'h12AE9,4);
TASK_PP(16'h12AEA,4);
TASK_PP(16'h12AEB,4);
TASK_PP(16'h12AEC,4);
TASK_PP(16'h12AED,4);
TASK_PP(16'h12AEE,4);
TASK_PP(16'h12AEF,4);
TASK_PP(16'h12AF0,4);
TASK_PP(16'h12AF1,4);
TASK_PP(16'h12AF2,4);
TASK_PP(16'h12AF3,4);
TASK_PP(16'h12AF4,4);
TASK_PP(16'h12AF5,4);
TASK_PP(16'h12AF6,4);
TASK_PP(16'h12AF7,4);
TASK_PP(16'h12AF8,4);
TASK_PP(16'h12AF9,4);
TASK_PP(16'h12AFA,4);
TASK_PP(16'h12AFB,4);
TASK_PP(16'h12AFC,4);
TASK_PP(16'h12AFD,4);
TASK_PP(16'h12AFE,4);
TASK_PP(16'h12AFF,4);
TASK_PP(16'h12B00,4);
TASK_PP(16'h12B01,4);
TASK_PP(16'h12B02,4);
TASK_PP(16'h12B03,4);
TASK_PP(16'h12B04,4);
TASK_PP(16'h12B05,4);
TASK_PP(16'h12B06,4);
TASK_PP(16'h12B07,4);
TASK_PP(16'h12B08,4);
TASK_PP(16'h12B09,4);
TASK_PP(16'h12B0A,4);
TASK_PP(16'h12B0B,4);
TASK_PP(16'h12B0C,4);
TASK_PP(16'h12B0D,4);
TASK_PP(16'h12B0E,4);
TASK_PP(16'h12B0F,4);
TASK_PP(16'h12B10,4);
TASK_PP(16'h12B11,4);
TASK_PP(16'h12B12,4);
TASK_PP(16'h12B13,4);
TASK_PP(16'h12B14,4);
TASK_PP(16'h12B15,4);
TASK_PP(16'h12B16,4);
TASK_PP(16'h12B17,4);
TASK_PP(16'h12B18,4);
TASK_PP(16'h12B19,4);
TASK_PP(16'h12B1A,4);
TASK_PP(16'h12B1B,4);
TASK_PP(16'h12B1C,4);
TASK_PP(16'h12B1D,4);
TASK_PP(16'h12B1E,4);
TASK_PP(16'h12B1F,4);
TASK_PP(16'h12B20,4);
TASK_PP(16'h12B21,4);
TASK_PP(16'h12B22,4);
TASK_PP(16'h12B23,4);
TASK_PP(16'h12B24,4);
TASK_PP(16'h12B25,4);
TASK_PP(16'h12B26,4);
TASK_PP(16'h12B27,4);
TASK_PP(16'h12B28,4);
TASK_PP(16'h12B29,4);
TASK_PP(16'h12B2A,4);
TASK_PP(16'h12B2B,4);
TASK_PP(16'h12B2C,4);
TASK_PP(16'h12B2D,4);
TASK_PP(16'h12B2E,4);
TASK_PP(16'h12B2F,4);
TASK_PP(16'h12B30,4);
TASK_PP(16'h12B31,4);
TASK_PP(16'h12B32,4);
TASK_PP(16'h12B33,4);
TASK_PP(16'h12B34,4);
TASK_PP(16'h12B35,4);
TASK_PP(16'h12B36,4);
TASK_PP(16'h12B37,4);
TASK_PP(16'h12B38,4);
TASK_PP(16'h12B39,4);
TASK_PP(16'h12B3A,4);
TASK_PP(16'h12B3B,4);
TASK_PP(16'h12B3C,4);
TASK_PP(16'h12B3D,4);
TASK_PP(16'h12B3E,4);
TASK_PP(16'h12B3F,4);
TASK_PP(16'h12B40,4);
TASK_PP(16'h12B41,4);
TASK_PP(16'h12B42,4);
TASK_PP(16'h12B43,4);
TASK_PP(16'h12B44,4);
TASK_PP(16'h12B45,4);
TASK_PP(16'h12B46,4);
TASK_PP(16'h12B47,4);
TASK_PP(16'h12B48,4);
TASK_PP(16'h12B49,4);
TASK_PP(16'h12B4A,4);
TASK_PP(16'h12B4B,4);
TASK_PP(16'h12B4C,4);
TASK_PP(16'h12B4D,4);
TASK_PP(16'h12B4E,4);
TASK_PP(16'h12B4F,4);
TASK_PP(16'h12B50,4);
TASK_PP(16'h12B51,4);
TASK_PP(16'h12B52,4);
TASK_PP(16'h12B53,4);
TASK_PP(16'h12B54,4);
TASK_PP(16'h12B55,4);
TASK_PP(16'h12B56,4);
TASK_PP(16'h12B57,4);
TASK_PP(16'h12B58,4);
TASK_PP(16'h12B59,4);
TASK_PP(16'h12B5A,4);
TASK_PP(16'h12B5B,4);
TASK_PP(16'h12B5C,4);
TASK_PP(16'h12B5D,4);
TASK_PP(16'h12B5E,4);
TASK_PP(16'h12B5F,4);
TASK_PP(16'h12B60,4);
TASK_PP(16'h12B61,4);
TASK_PP(16'h12B62,4);
TASK_PP(16'h12B63,4);
TASK_PP(16'h12B64,4);
TASK_PP(16'h12B65,4);
TASK_PP(16'h12B66,4);
TASK_PP(16'h12B67,4);
TASK_PP(16'h12B68,4);
TASK_PP(16'h12B69,4);
TASK_PP(16'h12B6A,4);
TASK_PP(16'h12B6B,4);
TASK_PP(16'h12B6C,4);
TASK_PP(16'h12B6D,4);
TASK_PP(16'h12B6E,4);
TASK_PP(16'h12B6F,4);
TASK_PP(16'h12B70,4);
TASK_PP(16'h12B71,4);
TASK_PP(16'h12B72,4);
TASK_PP(16'h12B73,4);
TASK_PP(16'h12B74,4);
TASK_PP(16'h12B75,4);
TASK_PP(16'h12B76,4);
TASK_PP(16'h12B77,4);
TASK_PP(16'h12B78,4);
TASK_PP(16'h12B79,4);
TASK_PP(16'h12B7A,4);
TASK_PP(16'h12B7B,4);
TASK_PP(16'h12B7C,4);
TASK_PP(16'h12B7D,4);
TASK_PP(16'h12B7E,4);
TASK_PP(16'h12B7F,4);
TASK_PP(16'h12B80,4);
TASK_PP(16'h12B81,4);
TASK_PP(16'h12B82,4);
TASK_PP(16'h12B83,4);
TASK_PP(16'h12B84,4);
TASK_PP(16'h12B85,4);
TASK_PP(16'h12B86,4);
TASK_PP(16'h12B87,4);
TASK_PP(16'h12B88,4);
TASK_PP(16'h12B89,4);
TASK_PP(16'h12B8A,4);
TASK_PP(16'h12B8B,4);
TASK_PP(16'h12B8C,4);
TASK_PP(16'h12B8D,4);
TASK_PP(16'h12B8E,4);
TASK_PP(16'h12B8F,4);
TASK_PP(16'h12B90,4);
TASK_PP(16'h12B91,4);
TASK_PP(16'h12B92,4);
TASK_PP(16'h12B93,4);
TASK_PP(16'h12B94,4);
TASK_PP(16'h12B95,4);
TASK_PP(16'h12B96,4);
TASK_PP(16'h12B97,4);
TASK_PP(16'h12B98,4);
TASK_PP(16'h12B99,4);
TASK_PP(16'h12B9A,4);
TASK_PP(16'h12B9B,4);
TASK_PP(16'h12B9C,4);
TASK_PP(16'h12B9D,4);
TASK_PP(16'h12B9E,4);
TASK_PP(16'h12B9F,4);
TASK_PP(16'h12BA0,4);
TASK_PP(16'h12BA1,4);
TASK_PP(16'h12BA2,4);
TASK_PP(16'h12BA3,4);
TASK_PP(16'h12BA4,4);
TASK_PP(16'h12BA5,4);
TASK_PP(16'h12BA6,4);
TASK_PP(16'h12BA7,4);
TASK_PP(16'h12BA8,4);
TASK_PP(16'h12BA9,4);
TASK_PP(16'h12BAA,4);
TASK_PP(16'h12BAB,4);
TASK_PP(16'h12BAC,4);
TASK_PP(16'h12BAD,4);
TASK_PP(16'h12BAE,4);
TASK_PP(16'h12BAF,4);
TASK_PP(16'h12BB0,4);
TASK_PP(16'h12BB1,4);
TASK_PP(16'h12BB2,4);
TASK_PP(16'h12BB3,4);
TASK_PP(16'h12BB4,4);
TASK_PP(16'h12BB5,4);
TASK_PP(16'h12BB6,4);
TASK_PP(16'h12BB7,4);
TASK_PP(16'h12BB8,4);
TASK_PP(16'h12BB9,4);
TASK_PP(16'h12BBA,4);
TASK_PP(16'h12BBB,4);
TASK_PP(16'h12BBC,4);
TASK_PP(16'h12BBD,4);
TASK_PP(16'h12BBE,4);
TASK_PP(16'h12BBF,4);
TASK_PP(16'h12BC0,4);
TASK_PP(16'h12BC1,4);
TASK_PP(16'h12BC2,4);
TASK_PP(16'h12BC3,4);
TASK_PP(16'h12BC4,4);
TASK_PP(16'h12BC5,4);
TASK_PP(16'h12BC6,4);
TASK_PP(16'h12BC7,4);
TASK_PP(16'h12BC8,4);
TASK_PP(16'h12BC9,4);
TASK_PP(16'h12BCA,4);
TASK_PP(16'h12BCB,4);
TASK_PP(16'h12BCC,4);
TASK_PP(16'h12BCD,4);
TASK_PP(16'h12BCE,4);
TASK_PP(16'h12BCF,4);
TASK_PP(16'h12BD0,4);
TASK_PP(16'h12BD1,4);
TASK_PP(16'h12BD2,4);
TASK_PP(16'h12BD3,4);
TASK_PP(16'h12BD4,4);
TASK_PP(16'h12BD5,4);
TASK_PP(16'h12BD6,4);
TASK_PP(16'h12BD7,4);
TASK_PP(16'h12BD8,4);
TASK_PP(16'h12BD9,4);
TASK_PP(16'h12BDA,4);
TASK_PP(16'h12BDB,4);
TASK_PP(16'h12BDC,4);
TASK_PP(16'h12BDD,4);
TASK_PP(16'h12BDE,4);
TASK_PP(16'h12BDF,4);
TASK_PP(16'h12BE0,4);
TASK_PP(16'h12BE1,4);
TASK_PP(16'h12BE2,4);
TASK_PP(16'h12BE3,4);
TASK_PP(16'h12BE4,4);
TASK_PP(16'h12BE5,4);
TASK_PP(16'h12BE6,4);
TASK_PP(16'h12BE7,4);
TASK_PP(16'h12BE8,4);
TASK_PP(16'h12BE9,4);
TASK_PP(16'h12BEA,4);
TASK_PP(16'h12BEB,4);
TASK_PP(16'h12BEC,4);
TASK_PP(16'h12BED,4);
TASK_PP(16'h12BEE,4);
TASK_PP(16'h12BEF,4);
TASK_PP(16'h12BF0,4);
TASK_PP(16'h12BF1,4);
TASK_PP(16'h12BF2,4);
TASK_PP(16'h12BF3,4);
TASK_PP(16'h12BF4,4);
TASK_PP(16'h12BF5,4);
TASK_PP(16'h12BF6,4);
TASK_PP(16'h12BF7,4);
TASK_PP(16'h12BF8,4);
TASK_PP(16'h12BF9,4);
TASK_PP(16'h12BFA,4);
TASK_PP(16'h12BFB,4);
TASK_PP(16'h12BFC,4);
TASK_PP(16'h12BFD,4);
TASK_PP(16'h12BFE,4);
TASK_PP(16'h12BFF,4);
TASK_PP(16'h12C00,4);
TASK_PP(16'h12C01,4);
TASK_PP(16'h12C02,4);
TASK_PP(16'h12C03,4);
TASK_PP(16'h12C04,4);
TASK_PP(16'h12C05,4);
TASK_PP(16'h12C06,4);
TASK_PP(16'h12C07,4);
TASK_PP(16'h12C08,4);
TASK_PP(16'h12C09,4);
TASK_PP(16'h12C0A,4);
TASK_PP(16'h12C0B,4);
TASK_PP(16'h12C0C,4);
TASK_PP(16'h12C0D,4);
TASK_PP(16'h12C0E,4);
TASK_PP(16'h12C0F,4);
TASK_PP(16'h12C10,4);
TASK_PP(16'h12C11,4);
TASK_PP(16'h12C12,4);
TASK_PP(16'h12C13,4);
TASK_PP(16'h12C14,4);
TASK_PP(16'h12C15,4);
TASK_PP(16'h12C16,4);
TASK_PP(16'h12C17,4);
TASK_PP(16'h12C18,4);
TASK_PP(16'h12C19,4);
TASK_PP(16'h12C1A,4);
TASK_PP(16'h12C1B,4);
TASK_PP(16'h12C1C,4);
TASK_PP(16'h12C1D,4);
TASK_PP(16'h12C1E,4);
TASK_PP(16'h12C1F,4);
TASK_PP(16'h12C20,4);
TASK_PP(16'h12C21,4);
TASK_PP(16'h12C22,4);
TASK_PP(16'h12C23,4);
TASK_PP(16'h12C24,4);
TASK_PP(16'h12C25,4);
TASK_PP(16'h12C26,4);
TASK_PP(16'h12C27,4);
TASK_PP(16'h12C28,4);
TASK_PP(16'h12C29,4);
TASK_PP(16'h12C2A,4);
TASK_PP(16'h12C2B,4);
TASK_PP(16'h12C2C,4);
TASK_PP(16'h12C2D,4);
TASK_PP(16'h12C2E,4);
TASK_PP(16'h12C2F,4);
TASK_PP(16'h12C30,4);
TASK_PP(16'h12C31,4);
TASK_PP(16'h12C32,4);
TASK_PP(16'h12C33,4);
TASK_PP(16'h12C34,4);
TASK_PP(16'h12C35,4);
TASK_PP(16'h12C36,4);
TASK_PP(16'h12C37,4);
TASK_PP(16'h12C38,4);
TASK_PP(16'h12C39,4);
TASK_PP(16'h12C3A,4);
TASK_PP(16'h12C3B,4);
TASK_PP(16'h12C3C,4);
TASK_PP(16'h12C3D,4);
TASK_PP(16'h12C3E,4);
TASK_PP(16'h12C3F,4);
TASK_PP(16'h12C40,4);
TASK_PP(16'h12C41,4);
TASK_PP(16'h12C42,4);
TASK_PP(16'h12C43,4);
TASK_PP(16'h12C44,4);
TASK_PP(16'h12C45,4);
TASK_PP(16'h12C46,4);
TASK_PP(16'h12C47,4);
TASK_PP(16'h12C48,4);
TASK_PP(16'h12C49,4);
TASK_PP(16'h12C4A,4);
TASK_PP(16'h12C4B,4);
TASK_PP(16'h12C4C,4);
TASK_PP(16'h12C4D,4);
TASK_PP(16'h12C4E,4);
TASK_PP(16'h12C4F,4);
TASK_PP(16'h12C50,4);
TASK_PP(16'h12C51,4);
TASK_PP(16'h12C52,4);
TASK_PP(16'h12C53,4);
TASK_PP(16'h12C54,4);
TASK_PP(16'h12C55,4);
TASK_PP(16'h12C56,4);
TASK_PP(16'h12C57,4);
TASK_PP(16'h12C58,4);
TASK_PP(16'h12C59,4);
TASK_PP(16'h12C5A,4);
TASK_PP(16'h12C5B,4);
TASK_PP(16'h12C5C,4);
TASK_PP(16'h12C5D,4);
TASK_PP(16'h12C5E,4);
TASK_PP(16'h12C5F,4);
TASK_PP(16'h12C60,4);
TASK_PP(16'h12C61,4);
TASK_PP(16'h12C62,4);
TASK_PP(16'h12C63,4);
TASK_PP(16'h12C64,4);
TASK_PP(16'h12C65,4);
TASK_PP(16'h12C66,4);
TASK_PP(16'h12C67,4);
TASK_PP(16'h12C68,4);
TASK_PP(16'h12C69,4);
TASK_PP(16'h12C6A,4);
TASK_PP(16'h12C6B,4);
TASK_PP(16'h12C6C,4);
TASK_PP(16'h12C6D,4);
TASK_PP(16'h12C6E,4);
TASK_PP(16'h12C6F,4);
TASK_PP(16'h12C70,4);
TASK_PP(16'h12C71,4);
TASK_PP(16'h12C72,4);
TASK_PP(16'h12C73,4);
TASK_PP(16'h12C74,4);
TASK_PP(16'h12C75,4);
TASK_PP(16'h12C76,4);
TASK_PP(16'h12C77,4);
TASK_PP(16'h12C78,4);
TASK_PP(16'h12C79,4);
TASK_PP(16'h12C7A,4);
TASK_PP(16'h12C7B,4);
TASK_PP(16'h12C7C,4);
TASK_PP(16'h12C7D,4);
TASK_PP(16'h12C7E,4);
TASK_PP(16'h12C7F,4);
TASK_PP(16'h12C80,4);
TASK_PP(16'h12C81,4);
TASK_PP(16'h12C82,4);
TASK_PP(16'h12C83,4);
TASK_PP(16'h12C84,4);
TASK_PP(16'h12C85,4);
TASK_PP(16'h12C86,4);
TASK_PP(16'h12C87,4);
TASK_PP(16'h12C88,4);
TASK_PP(16'h12C89,4);
TASK_PP(16'h12C8A,4);
TASK_PP(16'h12C8B,4);
TASK_PP(16'h12C8C,4);
TASK_PP(16'h12C8D,4);
TASK_PP(16'h12C8E,4);
TASK_PP(16'h12C8F,4);
TASK_PP(16'h12C90,4);
TASK_PP(16'h12C91,4);
TASK_PP(16'h12C92,4);
TASK_PP(16'h12C93,4);
TASK_PP(16'h12C94,4);
TASK_PP(16'h12C95,4);
TASK_PP(16'h12C96,4);
TASK_PP(16'h12C97,4);
TASK_PP(16'h12C98,4);
TASK_PP(16'h12C99,4);
TASK_PP(16'h12C9A,4);
TASK_PP(16'h12C9B,4);
TASK_PP(16'h12C9C,4);
TASK_PP(16'h12C9D,4);
TASK_PP(16'h12C9E,4);
TASK_PP(16'h12C9F,4);
TASK_PP(16'h12CA0,4);
TASK_PP(16'h12CA1,4);
TASK_PP(16'h12CA2,4);
TASK_PP(16'h12CA3,4);
TASK_PP(16'h12CA4,4);
TASK_PP(16'h12CA5,4);
TASK_PP(16'h12CA6,4);
TASK_PP(16'h12CA7,4);
TASK_PP(16'h12CA8,4);
TASK_PP(16'h12CA9,4);
TASK_PP(16'h12CAA,4);
TASK_PP(16'h12CAB,4);
TASK_PP(16'h12CAC,4);
TASK_PP(16'h12CAD,4);
TASK_PP(16'h12CAE,4);
TASK_PP(16'h12CAF,4);
TASK_PP(16'h12CB0,4);
TASK_PP(16'h12CB1,4);
TASK_PP(16'h12CB2,4);
TASK_PP(16'h12CB3,4);
TASK_PP(16'h12CB4,4);
TASK_PP(16'h12CB5,4);
TASK_PP(16'h12CB6,4);
TASK_PP(16'h12CB7,4);
TASK_PP(16'h12CB8,4);
TASK_PP(16'h12CB9,4);
TASK_PP(16'h12CBA,4);
TASK_PP(16'h12CBB,4);
TASK_PP(16'h12CBC,4);
TASK_PP(16'h12CBD,4);
TASK_PP(16'h12CBE,4);
TASK_PP(16'h12CBF,4);
TASK_PP(16'h12CC0,4);
TASK_PP(16'h12CC1,4);
TASK_PP(16'h12CC2,4);
TASK_PP(16'h12CC3,4);
TASK_PP(16'h12CC4,4);
TASK_PP(16'h12CC5,4);
TASK_PP(16'h12CC6,4);
TASK_PP(16'h12CC7,4);
TASK_PP(16'h12CC8,4);
TASK_PP(16'h12CC9,4);
TASK_PP(16'h12CCA,4);
TASK_PP(16'h12CCB,4);
TASK_PP(16'h12CCC,4);
TASK_PP(16'h12CCD,4);
TASK_PP(16'h12CCE,4);
TASK_PP(16'h12CCF,4);
TASK_PP(16'h12CD0,4);
TASK_PP(16'h12CD1,4);
TASK_PP(16'h12CD2,4);
TASK_PP(16'h12CD3,4);
TASK_PP(16'h12CD4,4);
TASK_PP(16'h12CD5,4);
TASK_PP(16'h12CD6,4);
TASK_PP(16'h12CD7,4);
TASK_PP(16'h12CD8,4);
TASK_PP(16'h12CD9,4);
TASK_PP(16'h12CDA,4);
TASK_PP(16'h12CDB,4);
TASK_PP(16'h12CDC,4);
TASK_PP(16'h12CDD,4);
TASK_PP(16'h12CDE,4);
TASK_PP(16'h12CDF,4);
TASK_PP(16'h12CE0,4);
TASK_PP(16'h12CE1,4);
TASK_PP(16'h12CE2,4);
TASK_PP(16'h12CE3,4);
TASK_PP(16'h12CE4,4);
TASK_PP(16'h12CE5,4);
TASK_PP(16'h12CE6,4);
TASK_PP(16'h12CE7,4);
TASK_PP(16'h12CE8,4);
TASK_PP(16'h12CE9,4);
TASK_PP(16'h12CEA,4);
TASK_PP(16'h12CEB,4);
TASK_PP(16'h12CEC,4);
TASK_PP(16'h12CED,4);
TASK_PP(16'h12CEE,4);
TASK_PP(16'h12CEF,4);
TASK_PP(16'h12CF0,4);
TASK_PP(16'h12CF1,4);
TASK_PP(16'h12CF2,4);
TASK_PP(16'h12CF3,4);
TASK_PP(16'h12CF4,4);
TASK_PP(16'h12CF5,4);
TASK_PP(16'h12CF6,4);
TASK_PP(16'h12CF7,4);
TASK_PP(16'h12CF8,4);
TASK_PP(16'h12CF9,4);
TASK_PP(16'h12CFA,4);
TASK_PP(16'h12CFB,4);
TASK_PP(16'h12CFC,4);
TASK_PP(16'h12CFD,4);
TASK_PP(16'h12CFE,4);
TASK_PP(16'h12CFF,4);
TASK_PP(16'h12D00,4);
TASK_PP(16'h12D01,4);
TASK_PP(16'h12D02,4);
TASK_PP(16'h12D03,4);
TASK_PP(16'h12D04,4);
TASK_PP(16'h12D05,4);
TASK_PP(16'h12D06,4);
TASK_PP(16'h12D07,4);
TASK_PP(16'h12D08,4);
TASK_PP(16'h12D09,4);
TASK_PP(16'h12D0A,4);
TASK_PP(16'h12D0B,4);
TASK_PP(16'h12D0C,4);
TASK_PP(16'h12D0D,4);
TASK_PP(16'h12D0E,4);
TASK_PP(16'h12D0F,4);
TASK_PP(16'h12D10,4);
TASK_PP(16'h12D11,4);
TASK_PP(16'h12D12,4);
TASK_PP(16'h12D13,4);
TASK_PP(16'h12D14,4);
TASK_PP(16'h12D15,4);
TASK_PP(16'h12D16,4);
TASK_PP(16'h12D17,4);
TASK_PP(16'h12D18,4);
TASK_PP(16'h12D19,4);
TASK_PP(16'h12D1A,4);
TASK_PP(16'h12D1B,4);
TASK_PP(16'h12D1C,4);
TASK_PP(16'h12D1D,4);
TASK_PP(16'h12D1E,4);
TASK_PP(16'h12D1F,4);
TASK_PP(16'h12D20,4);
TASK_PP(16'h12D21,4);
TASK_PP(16'h12D22,4);
TASK_PP(16'h12D23,4);
TASK_PP(16'h12D24,4);
TASK_PP(16'h12D25,4);
TASK_PP(16'h12D26,4);
TASK_PP(16'h12D27,4);
TASK_PP(16'h12D28,4);
TASK_PP(16'h12D29,4);
TASK_PP(16'h12D2A,4);
TASK_PP(16'h12D2B,4);
TASK_PP(16'h12D2C,4);
TASK_PP(16'h12D2D,4);
TASK_PP(16'h12D2E,4);
TASK_PP(16'h12D2F,4);
TASK_PP(16'h12D30,4);
TASK_PP(16'h12D31,4);
TASK_PP(16'h12D32,4);
TASK_PP(16'h12D33,4);
TASK_PP(16'h12D34,4);
TASK_PP(16'h12D35,4);
TASK_PP(16'h12D36,4);
TASK_PP(16'h12D37,4);
TASK_PP(16'h12D38,4);
TASK_PP(16'h12D39,4);
TASK_PP(16'h12D3A,4);
TASK_PP(16'h12D3B,4);
TASK_PP(16'h12D3C,4);
TASK_PP(16'h12D3D,4);
TASK_PP(16'h12D3E,4);
TASK_PP(16'h12D3F,4);
TASK_PP(16'h12D40,4);
TASK_PP(16'h12D41,4);
TASK_PP(16'h12D42,4);
TASK_PP(16'h12D43,4);
TASK_PP(16'h12D44,4);
TASK_PP(16'h12D45,4);
TASK_PP(16'h12D46,4);
TASK_PP(16'h12D47,4);
TASK_PP(16'h12D48,4);
TASK_PP(16'h12D49,4);
TASK_PP(16'h12D4A,4);
TASK_PP(16'h12D4B,4);
TASK_PP(16'h12D4C,4);
TASK_PP(16'h12D4D,4);
TASK_PP(16'h12D4E,4);
TASK_PP(16'h12D4F,4);
TASK_PP(16'h12D50,4);
TASK_PP(16'h12D51,4);
TASK_PP(16'h12D52,4);
TASK_PP(16'h12D53,4);
TASK_PP(16'h12D54,4);
TASK_PP(16'h12D55,4);
TASK_PP(16'h12D56,4);
TASK_PP(16'h12D57,4);
TASK_PP(16'h12D58,4);
TASK_PP(16'h12D59,4);
TASK_PP(16'h12D5A,4);
TASK_PP(16'h12D5B,4);
TASK_PP(16'h12D5C,4);
TASK_PP(16'h12D5D,4);
TASK_PP(16'h12D5E,4);
TASK_PP(16'h12D5F,4);
TASK_PP(16'h12D60,4);
TASK_PP(16'h12D61,4);
TASK_PP(16'h12D62,4);
TASK_PP(16'h12D63,4);
TASK_PP(16'h12D64,4);
TASK_PP(16'h12D65,4);
TASK_PP(16'h12D66,4);
TASK_PP(16'h12D67,4);
TASK_PP(16'h12D68,4);
TASK_PP(16'h12D69,4);
TASK_PP(16'h12D6A,4);
TASK_PP(16'h12D6B,4);
TASK_PP(16'h12D6C,4);
TASK_PP(16'h12D6D,4);
TASK_PP(16'h12D6E,4);
TASK_PP(16'h12D6F,4);
TASK_PP(16'h12D70,4);
TASK_PP(16'h12D71,4);
TASK_PP(16'h12D72,4);
TASK_PP(16'h12D73,4);
TASK_PP(16'h12D74,4);
TASK_PP(16'h12D75,4);
TASK_PP(16'h12D76,4);
TASK_PP(16'h12D77,4);
TASK_PP(16'h12D78,4);
TASK_PP(16'h12D79,4);
TASK_PP(16'h12D7A,4);
TASK_PP(16'h12D7B,4);
TASK_PP(16'h12D7C,4);
TASK_PP(16'h12D7D,4);
TASK_PP(16'h12D7E,4);
TASK_PP(16'h12D7F,4);
TASK_PP(16'h12D80,4);
TASK_PP(16'h12D81,4);
TASK_PP(16'h12D82,4);
TASK_PP(16'h12D83,4);
TASK_PP(16'h12D84,4);
TASK_PP(16'h12D85,4);
TASK_PP(16'h12D86,4);
TASK_PP(16'h12D87,4);
TASK_PP(16'h12D88,4);
TASK_PP(16'h12D89,4);
TASK_PP(16'h12D8A,4);
TASK_PP(16'h12D8B,4);
TASK_PP(16'h12D8C,4);
TASK_PP(16'h12D8D,4);
TASK_PP(16'h12D8E,4);
TASK_PP(16'h12D8F,4);
TASK_PP(16'h12D90,4);
TASK_PP(16'h12D91,4);
TASK_PP(16'h12D92,4);
TASK_PP(16'h12D93,4);
TASK_PP(16'h12D94,4);
TASK_PP(16'h12D95,4);
TASK_PP(16'h12D96,4);
TASK_PP(16'h12D97,4);
TASK_PP(16'h12D98,4);
TASK_PP(16'h12D99,4);
TASK_PP(16'h12D9A,4);
TASK_PP(16'h12D9B,4);
TASK_PP(16'h12D9C,4);
TASK_PP(16'h12D9D,4);
TASK_PP(16'h12D9E,4);
TASK_PP(16'h12D9F,4);
TASK_PP(16'h12DA0,4);
TASK_PP(16'h12DA1,4);
TASK_PP(16'h12DA2,4);
TASK_PP(16'h12DA3,4);
TASK_PP(16'h12DA4,4);
TASK_PP(16'h12DA5,4);
TASK_PP(16'h12DA6,4);
TASK_PP(16'h12DA7,4);
TASK_PP(16'h12DA8,4);
TASK_PP(16'h12DA9,4);
TASK_PP(16'h12DAA,4);
TASK_PP(16'h12DAB,4);
TASK_PP(16'h12DAC,4);
TASK_PP(16'h12DAD,4);
TASK_PP(16'h12DAE,4);
TASK_PP(16'h12DAF,4);
TASK_PP(16'h12DB0,4);
TASK_PP(16'h12DB1,4);
TASK_PP(16'h12DB2,4);
TASK_PP(16'h12DB3,4);
TASK_PP(16'h12DB4,4);
TASK_PP(16'h12DB5,4);
TASK_PP(16'h12DB6,4);
TASK_PP(16'h12DB7,4);
TASK_PP(16'h12DB8,4);
TASK_PP(16'h12DB9,4);
TASK_PP(16'h12DBA,4);
TASK_PP(16'h12DBB,4);
TASK_PP(16'h12DBC,4);
TASK_PP(16'h12DBD,4);
TASK_PP(16'h12DBE,4);
TASK_PP(16'h12DBF,4);
TASK_PP(16'h12DC0,4);
TASK_PP(16'h12DC1,4);
TASK_PP(16'h12DC2,4);
TASK_PP(16'h12DC3,4);
TASK_PP(16'h12DC4,4);
TASK_PP(16'h12DC5,4);
TASK_PP(16'h12DC6,4);
TASK_PP(16'h12DC7,4);
TASK_PP(16'h12DC8,4);
TASK_PP(16'h12DC9,4);
TASK_PP(16'h12DCA,4);
TASK_PP(16'h12DCB,4);
TASK_PP(16'h12DCC,4);
TASK_PP(16'h12DCD,4);
TASK_PP(16'h12DCE,4);
TASK_PP(16'h12DCF,4);
TASK_PP(16'h12DD0,4);
TASK_PP(16'h12DD1,4);
TASK_PP(16'h12DD2,4);
TASK_PP(16'h12DD3,4);
TASK_PP(16'h12DD4,4);
TASK_PP(16'h12DD5,4);
TASK_PP(16'h12DD6,4);
TASK_PP(16'h12DD7,4);
TASK_PP(16'h12DD8,4);
TASK_PP(16'h12DD9,4);
TASK_PP(16'h12DDA,4);
TASK_PP(16'h12DDB,4);
TASK_PP(16'h12DDC,4);
TASK_PP(16'h12DDD,4);
TASK_PP(16'h12DDE,4);
TASK_PP(16'h12DDF,4);
TASK_PP(16'h12DE0,4);
TASK_PP(16'h12DE1,4);
TASK_PP(16'h12DE2,4);
TASK_PP(16'h12DE3,4);
TASK_PP(16'h12DE4,4);
TASK_PP(16'h12DE5,4);
TASK_PP(16'h12DE6,4);
TASK_PP(16'h12DE7,4);
TASK_PP(16'h12DE8,4);
TASK_PP(16'h12DE9,4);
TASK_PP(16'h12DEA,4);
TASK_PP(16'h12DEB,4);
TASK_PP(16'h12DEC,4);
TASK_PP(16'h12DED,4);
TASK_PP(16'h12DEE,4);
TASK_PP(16'h12DEF,4);
TASK_PP(16'h12DF0,4);
TASK_PP(16'h12DF1,4);
TASK_PP(16'h12DF2,4);
TASK_PP(16'h12DF3,4);
TASK_PP(16'h12DF4,4);
TASK_PP(16'h12DF5,4);
TASK_PP(16'h12DF6,4);
TASK_PP(16'h12DF7,4);
TASK_PP(16'h12DF8,4);
TASK_PP(16'h12DF9,4);
TASK_PP(16'h12DFA,4);
TASK_PP(16'h12DFB,4);
TASK_PP(16'h12DFC,4);
TASK_PP(16'h12DFD,4);
TASK_PP(16'h12DFE,4);
TASK_PP(16'h12DFF,4);
TASK_PP(16'h12E00,4);
TASK_PP(16'h12E01,4);
TASK_PP(16'h12E02,4);
TASK_PP(16'h12E03,4);
TASK_PP(16'h12E04,4);
TASK_PP(16'h12E05,4);
TASK_PP(16'h12E06,4);
TASK_PP(16'h12E07,4);
TASK_PP(16'h12E08,4);
TASK_PP(16'h12E09,4);
TASK_PP(16'h12E0A,4);
TASK_PP(16'h12E0B,4);
TASK_PP(16'h12E0C,4);
TASK_PP(16'h12E0D,4);
TASK_PP(16'h12E0E,4);
TASK_PP(16'h12E0F,4);
TASK_PP(16'h12E10,4);
TASK_PP(16'h12E11,4);
TASK_PP(16'h12E12,4);
TASK_PP(16'h12E13,4);
TASK_PP(16'h12E14,4);
TASK_PP(16'h12E15,4);
TASK_PP(16'h12E16,4);
TASK_PP(16'h12E17,4);
TASK_PP(16'h12E18,4);
TASK_PP(16'h12E19,4);
TASK_PP(16'h12E1A,4);
TASK_PP(16'h12E1B,4);
TASK_PP(16'h12E1C,4);
TASK_PP(16'h12E1D,4);
TASK_PP(16'h12E1E,4);
TASK_PP(16'h12E1F,4);
TASK_PP(16'h12E20,4);
TASK_PP(16'h12E21,4);
TASK_PP(16'h12E22,4);
TASK_PP(16'h12E23,4);
TASK_PP(16'h12E24,4);
TASK_PP(16'h12E25,4);
TASK_PP(16'h12E26,4);
TASK_PP(16'h12E27,4);
TASK_PP(16'h12E28,4);
TASK_PP(16'h12E29,4);
TASK_PP(16'h12E2A,4);
TASK_PP(16'h12E2B,4);
TASK_PP(16'h12E2C,4);
TASK_PP(16'h12E2D,4);
TASK_PP(16'h12E2E,4);
TASK_PP(16'h12E2F,4);
TASK_PP(16'h12E30,4);
TASK_PP(16'h12E31,4);
TASK_PP(16'h12E32,4);
TASK_PP(16'h12E33,4);
TASK_PP(16'h12E34,4);
TASK_PP(16'h12E35,4);
TASK_PP(16'h12E36,4);
TASK_PP(16'h12E37,4);
TASK_PP(16'h12E38,4);
TASK_PP(16'h12E39,4);
TASK_PP(16'h12E3A,4);
TASK_PP(16'h12E3B,4);
TASK_PP(16'h12E3C,4);
TASK_PP(16'h12E3D,4);
TASK_PP(16'h12E3E,4);
TASK_PP(16'h12E3F,4);
TASK_PP(16'h12E40,4);
TASK_PP(16'h12E41,4);
TASK_PP(16'h12E42,4);
TASK_PP(16'h12E43,4);
TASK_PP(16'h12E44,4);
TASK_PP(16'h12E45,4);
TASK_PP(16'h12E46,4);
TASK_PP(16'h12E47,4);
TASK_PP(16'h12E48,4);
TASK_PP(16'h12E49,4);
TASK_PP(16'h12E4A,4);
TASK_PP(16'h12E4B,4);
TASK_PP(16'h12E4C,4);
TASK_PP(16'h12E4D,4);
TASK_PP(16'h12E4E,4);
TASK_PP(16'h12E4F,4);
TASK_PP(16'h12E50,4);
TASK_PP(16'h12E51,4);
TASK_PP(16'h12E52,4);
TASK_PP(16'h12E53,4);
TASK_PP(16'h12E54,4);
TASK_PP(16'h12E55,4);
TASK_PP(16'h12E56,4);
TASK_PP(16'h12E57,4);
TASK_PP(16'h12E58,4);
TASK_PP(16'h12E59,4);
TASK_PP(16'h12E5A,4);
TASK_PP(16'h12E5B,4);
TASK_PP(16'h12E5C,4);
TASK_PP(16'h12E5D,4);
TASK_PP(16'h12E5E,4);
TASK_PP(16'h12E5F,4);
TASK_PP(16'h12E60,4);
TASK_PP(16'h12E61,4);
TASK_PP(16'h12E62,4);
TASK_PP(16'h12E63,4);
TASK_PP(16'h12E64,4);
TASK_PP(16'h12E65,4);
TASK_PP(16'h12E66,4);
TASK_PP(16'h12E67,4);
TASK_PP(16'h12E68,4);
TASK_PP(16'h12E69,4);
TASK_PP(16'h12E6A,4);
TASK_PP(16'h12E6B,4);
TASK_PP(16'h12E6C,4);
TASK_PP(16'h12E6D,4);
TASK_PP(16'h12E6E,4);
TASK_PP(16'h12E6F,4);
TASK_PP(16'h12E70,4);
TASK_PP(16'h12E71,4);
TASK_PP(16'h12E72,4);
TASK_PP(16'h12E73,4);
TASK_PP(16'h12E74,4);
TASK_PP(16'h12E75,4);
TASK_PP(16'h12E76,4);
TASK_PP(16'h12E77,4);
TASK_PP(16'h12E78,4);
TASK_PP(16'h12E79,4);
TASK_PP(16'h12E7A,4);
TASK_PP(16'h12E7B,4);
TASK_PP(16'h12E7C,4);
TASK_PP(16'h12E7D,4);
TASK_PP(16'h12E7E,4);
TASK_PP(16'h12E7F,4);
TASK_PP(16'h12E80,4);
TASK_PP(16'h12E81,4);
TASK_PP(16'h12E82,4);
TASK_PP(16'h12E83,4);
TASK_PP(16'h12E84,4);
TASK_PP(16'h12E85,4);
TASK_PP(16'h12E86,4);
TASK_PP(16'h12E87,4);
TASK_PP(16'h12E88,4);
TASK_PP(16'h12E89,4);
TASK_PP(16'h12E8A,4);
TASK_PP(16'h12E8B,4);
TASK_PP(16'h12E8C,4);
TASK_PP(16'h12E8D,4);
TASK_PP(16'h12E8E,4);
TASK_PP(16'h12E8F,4);
TASK_PP(16'h12E90,4);
TASK_PP(16'h12E91,4);
TASK_PP(16'h12E92,4);
TASK_PP(16'h12E93,4);
TASK_PP(16'h12E94,4);
TASK_PP(16'h12E95,4);
TASK_PP(16'h12E96,4);
TASK_PP(16'h12E97,4);
TASK_PP(16'h12E98,4);
TASK_PP(16'h12E99,4);
TASK_PP(16'h12E9A,4);
TASK_PP(16'h12E9B,4);
TASK_PP(16'h12E9C,4);
TASK_PP(16'h12E9D,4);
TASK_PP(16'h12E9E,4);
TASK_PP(16'h12E9F,4);
TASK_PP(16'h12EA0,4);
TASK_PP(16'h12EA1,4);
TASK_PP(16'h12EA2,4);
TASK_PP(16'h12EA3,4);
TASK_PP(16'h12EA4,4);
TASK_PP(16'h12EA5,4);
TASK_PP(16'h12EA6,4);
TASK_PP(16'h12EA7,4);
TASK_PP(16'h12EA8,4);
TASK_PP(16'h12EA9,4);
TASK_PP(16'h12EAA,4);
TASK_PP(16'h12EAB,4);
TASK_PP(16'h12EAC,4);
TASK_PP(16'h12EAD,4);
TASK_PP(16'h12EAE,4);
TASK_PP(16'h12EAF,4);
TASK_PP(16'h12EB0,4);
TASK_PP(16'h12EB1,4);
TASK_PP(16'h12EB2,4);
TASK_PP(16'h12EB3,4);
TASK_PP(16'h12EB4,4);
TASK_PP(16'h12EB5,4);
TASK_PP(16'h12EB6,4);
TASK_PP(16'h12EB7,4);
TASK_PP(16'h12EB8,4);
TASK_PP(16'h12EB9,4);
TASK_PP(16'h12EBA,4);
TASK_PP(16'h12EBB,4);
TASK_PP(16'h12EBC,4);
TASK_PP(16'h12EBD,4);
TASK_PP(16'h12EBE,4);
TASK_PP(16'h12EBF,4);
TASK_PP(16'h12EC0,4);
TASK_PP(16'h12EC1,4);
TASK_PP(16'h12EC2,4);
TASK_PP(16'h12EC3,4);
TASK_PP(16'h12EC4,4);
TASK_PP(16'h12EC5,4);
TASK_PP(16'h12EC6,4);
TASK_PP(16'h12EC7,4);
TASK_PP(16'h12EC8,4);
TASK_PP(16'h12EC9,4);
TASK_PP(16'h12ECA,4);
TASK_PP(16'h12ECB,4);
TASK_PP(16'h12ECC,4);
TASK_PP(16'h12ECD,4);
TASK_PP(16'h12ECE,4);
TASK_PP(16'h12ECF,4);
TASK_PP(16'h12ED0,4);
TASK_PP(16'h12ED1,4);
TASK_PP(16'h12ED2,4);
TASK_PP(16'h12ED3,4);
TASK_PP(16'h12ED4,4);
TASK_PP(16'h12ED5,4);
TASK_PP(16'h12ED6,4);
TASK_PP(16'h12ED7,4);
TASK_PP(16'h12ED8,4);
TASK_PP(16'h12ED9,4);
TASK_PP(16'h12EDA,4);
TASK_PP(16'h12EDB,4);
TASK_PP(16'h12EDC,4);
TASK_PP(16'h12EDD,4);
TASK_PP(16'h12EDE,4);
TASK_PP(16'h12EDF,4);
TASK_PP(16'h12EE0,4);
TASK_PP(16'h12EE1,4);
TASK_PP(16'h12EE2,4);
TASK_PP(16'h12EE3,4);
TASK_PP(16'h12EE4,4);
TASK_PP(16'h12EE5,4);
TASK_PP(16'h12EE6,4);
TASK_PP(16'h12EE7,4);
TASK_PP(16'h12EE8,4);
TASK_PP(16'h12EE9,4);
TASK_PP(16'h12EEA,4);
TASK_PP(16'h12EEB,4);
TASK_PP(16'h12EEC,4);
TASK_PP(16'h12EED,4);
TASK_PP(16'h12EEE,4);
TASK_PP(16'h12EEF,4);
TASK_PP(16'h12EF0,4);
TASK_PP(16'h12EF1,4);
TASK_PP(16'h12EF2,4);
TASK_PP(16'h12EF3,4);
TASK_PP(16'h12EF4,4);
TASK_PP(16'h12EF5,4);
TASK_PP(16'h12EF6,4);
TASK_PP(16'h12EF7,4);
TASK_PP(16'h12EF8,4);
TASK_PP(16'h12EF9,4);
TASK_PP(16'h12EFA,4);
TASK_PP(16'h12EFB,4);
TASK_PP(16'h12EFC,4);
TASK_PP(16'h12EFD,4);
TASK_PP(16'h12EFE,4);
TASK_PP(16'h12EFF,4);
TASK_PP(16'h12F00,4);
TASK_PP(16'h12F01,4);
TASK_PP(16'h12F02,4);
TASK_PP(16'h12F03,4);
TASK_PP(16'h12F04,4);
TASK_PP(16'h12F05,4);
TASK_PP(16'h12F06,4);
TASK_PP(16'h12F07,4);
TASK_PP(16'h12F08,4);
TASK_PP(16'h12F09,4);
TASK_PP(16'h12F0A,4);
TASK_PP(16'h12F0B,4);
TASK_PP(16'h12F0C,4);
TASK_PP(16'h12F0D,4);
TASK_PP(16'h12F0E,4);
TASK_PP(16'h12F0F,4);
TASK_PP(16'h12F10,4);
TASK_PP(16'h12F11,4);
TASK_PP(16'h12F12,4);
TASK_PP(16'h12F13,4);
TASK_PP(16'h12F14,4);
TASK_PP(16'h12F15,4);
TASK_PP(16'h12F16,4);
TASK_PP(16'h12F17,4);
TASK_PP(16'h12F18,4);
TASK_PP(16'h12F19,4);
TASK_PP(16'h12F1A,4);
TASK_PP(16'h12F1B,4);
TASK_PP(16'h12F1C,4);
TASK_PP(16'h12F1D,4);
TASK_PP(16'h12F1E,4);
TASK_PP(16'h12F1F,4);
TASK_PP(16'h12F20,4);
TASK_PP(16'h12F21,4);
TASK_PP(16'h12F22,4);
TASK_PP(16'h12F23,4);
TASK_PP(16'h12F24,4);
TASK_PP(16'h12F25,4);
TASK_PP(16'h12F26,4);
TASK_PP(16'h12F27,4);
TASK_PP(16'h12F28,4);
TASK_PP(16'h12F29,4);
TASK_PP(16'h12F2A,4);
TASK_PP(16'h12F2B,4);
TASK_PP(16'h12F2C,4);
TASK_PP(16'h12F2D,4);
TASK_PP(16'h12F2E,4);
TASK_PP(16'h12F2F,4);
TASK_PP(16'h12F30,4);
TASK_PP(16'h12F31,4);
TASK_PP(16'h12F32,4);
TASK_PP(16'h12F33,4);
TASK_PP(16'h12F34,4);
TASK_PP(16'h12F35,4);
TASK_PP(16'h12F36,4);
TASK_PP(16'h12F37,4);
TASK_PP(16'h12F38,4);
TASK_PP(16'h12F39,4);
TASK_PP(16'h12F3A,4);
TASK_PP(16'h12F3B,4);
TASK_PP(16'h12F3C,4);
TASK_PP(16'h12F3D,4);
TASK_PP(16'h12F3E,4);
TASK_PP(16'h12F3F,4);
TASK_PP(16'h12F40,4);
TASK_PP(16'h12F41,4);
TASK_PP(16'h12F42,4);
TASK_PP(16'h12F43,4);
TASK_PP(16'h12F44,4);
TASK_PP(16'h12F45,4);
TASK_PP(16'h12F46,4);
TASK_PP(16'h12F47,4);
TASK_PP(16'h12F48,4);
TASK_PP(16'h12F49,4);
TASK_PP(16'h12F4A,4);
TASK_PP(16'h12F4B,4);
TASK_PP(16'h12F4C,4);
TASK_PP(16'h12F4D,4);
TASK_PP(16'h12F4E,4);
TASK_PP(16'h12F4F,4);
TASK_PP(16'h12F50,4);
TASK_PP(16'h12F51,4);
TASK_PP(16'h12F52,4);
TASK_PP(16'h12F53,4);
TASK_PP(16'h12F54,4);
TASK_PP(16'h12F55,4);
TASK_PP(16'h12F56,4);
TASK_PP(16'h12F57,4);
TASK_PP(16'h12F58,4);
TASK_PP(16'h12F59,4);
TASK_PP(16'h12F5A,4);
TASK_PP(16'h12F5B,4);
TASK_PP(16'h12F5C,4);
TASK_PP(16'h12F5D,4);
TASK_PP(16'h12F5E,4);
TASK_PP(16'h12F5F,4);
TASK_PP(16'h12F60,4);
TASK_PP(16'h12F61,4);
TASK_PP(16'h12F62,4);
TASK_PP(16'h12F63,4);
TASK_PP(16'h12F64,4);
TASK_PP(16'h12F65,4);
TASK_PP(16'h12F66,4);
TASK_PP(16'h12F67,4);
TASK_PP(16'h12F68,4);
TASK_PP(16'h12F69,4);
TASK_PP(16'h12F6A,4);
TASK_PP(16'h12F6B,4);
TASK_PP(16'h12F6C,4);
TASK_PP(16'h12F6D,4);
TASK_PP(16'h12F6E,4);
TASK_PP(16'h12F6F,4);
TASK_PP(16'h12F70,4);
TASK_PP(16'h12F71,4);
TASK_PP(16'h12F72,4);
TASK_PP(16'h12F73,4);
TASK_PP(16'h12F74,4);
TASK_PP(16'h12F75,4);
TASK_PP(16'h12F76,4);
TASK_PP(16'h12F77,4);
TASK_PP(16'h12F78,4);
TASK_PP(16'h12F79,4);
TASK_PP(16'h12F7A,4);
TASK_PP(16'h12F7B,4);
TASK_PP(16'h12F7C,4);
TASK_PP(16'h12F7D,4);
TASK_PP(16'h12F7E,4);
TASK_PP(16'h12F7F,4);
TASK_PP(16'h12F80,4);
TASK_PP(16'h12F81,4);
TASK_PP(16'h12F82,4);
TASK_PP(16'h12F83,4);
TASK_PP(16'h12F84,4);
TASK_PP(16'h12F85,4);
TASK_PP(16'h12F86,4);
TASK_PP(16'h12F87,4);
TASK_PP(16'h12F88,4);
TASK_PP(16'h12F89,4);
TASK_PP(16'h12F8A,4);
TASK_PP(16'h12F8B,4);
TASK_PP(16'h12F8C,4);
TASK_PP(16'h12F8D,4);
TASK_PP(16'h12F8E,4);
TASK_PP(16'h12F8F,4);
TASK_PP(16'h12F90,4);
TASK_PP(16'h12F91,4);
TASK_PP(16'h12F92,4);
TASK_PP(16'h12F93,4);
TASK_PP(16'h12F94,4);
TASK_PP(16'h12F95,4);
TASK_PP(16'h12F96,4);
TASK_PP(16'h12F97,4);
TASK_PP(16'h12F98,4);
TASK_PP(16'h12F99,4);
TASK_PP(16'h12F9A,4);
TASK_PP(16'h12F9B,4);
TASK_PP(16'h12F9C,4);
TASK_PP(16'h12F9D,4);
TASK_PP(16'h12F9E,4);
TASK_PP(16'h12F9F,4);
TASK_PP(16'h12FA0,4);
TASK_PP(16'h12FA1,4);
TASK_PP(16'h12FA2,4);
TASK_PP(16'h12FA3,4);
TASK_PP(16'h12FA4,4);
TASK_PP(16'h12FA5,4);
TASK_PP(16'h12FA6,4);
TASK_PP(16'h12FA7,4);
TASK_PP(16'h12FA8,4);
TASK_PP(16'h12FA9,4);
TASK_PP(16'h12FAA,4);
TASK_PP(16'h12FAB,4);
TASK_PP(16'h12FAC,4);
TASK_PP(16'h12FAD,4);
TASK_PP(16'h12FAE,4);
TASK_PP(16'h12FAF,4);
TASK_PP(16'h12FB0,4);
TASK_PP(16'h12FB1,4);
TASK_PP(16'h12FB2,4);
TASK_PP(16'h12FB3,4);
TASK_PP(16'h12FB4,4);
TASK_PP(16'h12FB5,4);
TASK_PP(16'h12FB6,4);
TASK_PP(16'h12FB7,4);
TASK_PP(16'h12FB8,4);
TASK_PP(16'h12FB9,4);
TASK_PP(16'h12FBA,4);
TASK_PP(16'h12FBB,4);
TASK_PP(16'h12FBC,4);
TASK_PP(16'h12FBD,4);
TASK_PP(16'h12FBE,4);
TASK_PP(16'h12FBF,4);
TASK_PP(16'h12FC0,4);
TASK_PP(16'h12FC1,4);
TASK_PP(16'h12FC2,4);
TASK_PP(16'h12FC3,4);
TASK_PP(16'h12FC4,4);
TASK_PP(16'h12FC5,4);
TASK_PP(16'h12FC6,4);
TASK_PP(16'h12FC7,4);
TASK_PP(16'h12FC8,4);
TASK_PP(16'h12FC9,4);
TASK_PP(16'h12FCA,4);
TASK_PP(16'h12FCB,4);
TASK_PP(16'h12FCC,4);
TASK_PP(16'h12FCD,4);
TASK_PP(16'h12FCE,4);
TASK_PP(16'h12FCF,4);
TASK_PP(16'h12FD0,4);
TASK_PP(16'h12FD1,4);
TASK_PP(16'h12FD2,4);
TASK_PP(16'h12FD3,4);
TASK_PP(16'h12FD4,4);
TASK_PP(16'h12FD5,4);
TASK_PP(16'h12FD6,4);
TASK_PP(16'h12FD7,4);
TASK_PP(16'h12FD8,4);
TASK_PP(16'h12FD9,4);
TASK_PP(16'h12FDA,4);
TASK_PP(16'h12FDB,4);
TASK_PP(16'h12FDC,4);
TASK_PP(16'h12FDD,4);
TASK_PP(16'h12FDE,4);
TASK_PP(16'h12FDF,4);
TASK_PP(16'h12FE0,4);
TASK_PP(16'h12FE1,4);
TASK_PP(16'h12FE2,4);
TASK_PP(16'h12FE3,4);
TASK_PP(16'h12FE4,4);
TASK_PP(16'h12FE5,4);
TASK_PP(16'h12FE6,4);
TASK_PP(16'h12FE7,4);
TASK_PP(16'h12FE8,4);
TASK_PP(16'h12FE9,4);
TASK_PP(16'h12FEA,4);
TASK_PP(16'h12FEB,4);
TASK_PP(16'h12FEC,4);
TASK_PP(16'h12FED,4);
TASK_PP(16'h12FEE,4);
TASK_PP(16'h12FEF,4);
TASK_PP(16'h12FF0,4);
TASK_PP(16'h12FF1,4);
TASK_PP(16'h12FF2,4);
TASK_PP(16'h12FF3,4);
TASK_PP(16'h12FF4,4);
TASK_PP(16'h12FF5,4);
TASK_PP(16'h12FF6,4);
TASK_PP(16'h12FF7,4);
TASK_PP(16'h12FF8,4);
TASK_PP(16'h12FF9,4);
TASK_PP(16'h12FFA,4);
TASK_PP(16'h12FFB,4);
TASK_PP(16'h12FFC,4);
TASK_PP(16'h12FFD,4);
TASK_PP(16'h12FFE,4);
TASK_PP(16'h12FFF,4);
TASK_PP(16'h13000,4);
TASK_PP(16'h13001,4);
TASK_PP(16'h13002,4);
TASK_PP(16'h13003,4);
TASK_PP(16'h13004,4);
TASK_PP(16'h13005,4);
TASK_PP(16'h13006,4);
TASK_PP(16'h13007,4);
TASK_PP(16'h13008,4);
TASK_PP(16'h13009,4);
TASK_PP(16'h1300A,4);
TASK_PP(16'h1300B,4);
TASK_PP(16'h1300C,4);
TASK_PP(16'h1300D,4);
TASK_PP(16'h1300E,4);
TASK_PP(16'h1300F,4);
TASK_PP(16'h13010,4);
TASK_PP(16'h13011,4);
TASK_PP(16'h13012,4);
TASK_PP(16'h13013,4);
TASK_PP(16'h13014,4);
TASK_PP(16'h13015,4);
TASK_PP(16'h13016,4);
TASK_PP(16'h13017,4);
TASK_PP(16'h13018,4);
TASK_PP(16'h13019,4);
TASK_PP(16'h1301A,4);
TASK_PP(16'h1301B,4);
TASK_PP(16'h1301C,4);
TASK_PP(16'h1301D,4);
TASK_PP(16'h1301E,4);
TASK_PP(16'h1301F,4);
TASK_PP(16'h13020,4);
TASK_PP(16'h13021,4);
TASK_PP(16'h13022,4);
TASK_PP(16'h13023,4);
TASK_PP(16'h13024,4);
TASK_PP(16'h13025,4);
TASK_PP(16'h13026,4);
TASK_PP(16'h13027,4);
TASK_PP(16'h13028,4);
TASK_PP(16'h13029,4);
TASK_PP(16'h1302A,4);
TASK_PP(16'h1302B,4);
TASK_PP(16'h1302C,4);
TASK_PP(16'h1302D,4);
TASK_PP(16'h1302E,4);
TASK_PP(16'h1302F,4);
TASK_PP(16'h13030,4);
TASK_PP(16'h13031,4);
TASK_PP(16'h13032,4);
TASK_PP(16'h13033,4);
TASK_PP(16'h13034,4);
TASK_PP(16'h13035,4);
TASK_PP(16'h13036,4);
TASK_PP(16'h13037,4);
TASK_PP(16'h13038,4);
TASK_PP(16'h13039,4);
TASK_PP(16'h1303A,4);
TASK_PP(16'h1303B,4);
TASK_PP(16'h1303C,4);
TASK_PP(16'h1303D,4);
TASK_PP(16'h1303E,4);
TASK_PP(16'h1303F,4);
TASK_PP(16'h13040,4);
TASK_PP(16'h13041,4);
TASK_PP(16'h13042,4);
TASK_PP(16'h13043,4);
TASK_PP(16'h13044,4);
TASK_PP(16'h13045,4);
TASK_PP(16'h13046,4);
TASK_PP(16'h13047,4);
TASK_PP(16'h13048,4);
TASK_PP(16'h13049,4);
TASK_PP(16'h1304A,4);
TASK_PP(16'h1304B,4);
TASK_PP(16'h1304C,4);
TASK_PP(16'h1304D,4);
TASK_PP(16'h1304E,4);
TASK_PP(16'h1304F,4);
TASK_PP(16'h13050,4);
TASK_PP(16'h13051,4);
TASK_PP(16'h13052,4);
TASK_PP(16'h13053,4);
TASK_PP(16'h13054,4);
TASK_PP(16'h13055,4);
TASK_PP(16'h13056,4);
TASK_PP(16'h13057,4);
TASK_PP(16'h13058,4);
TASK_PP(16'h13059,4);
TASK_PP(16'h1305A,4);
TASK_PP(16'h1305B,4);
TASK_PP(16'h1305C,4);
TASK_PP(16'h1305D,4);
TASK_PP(16'h1305E,4);
TASK_PP(16'h1305F,4);
TASK_PP(16'h13060,4);
TASK_PP(16'h13061,4);
TASK_PP(16'h13062,4);
TASK_PP(16'h13063,4);
TASK_PP(16'h13064,4);
TASK_PP(16'h13065,4);
TASK_PP(16'h13066,4);
TASK_PP(16'h13067,4);
TASK_PP(16'h13068,4);
TASK_PP(16'h13069,4);
TASK_PP(16'h1306A,4);
TASK_PP(16'h1306B,4);
TASK_PP(16'h1306C,4);
TASK_PP(16'h1306D,4);
TASK_PP(16'h1306E,4);
TASK_PP(16'h1306F,4);
TASK_PP(16'h13070,4);
TASK_PP(16'h13071,4);
TASK_PP(16'h13072,4);
TASK_PP(16'h13073,4);
TASK_PP(16'h13074,4);
TASK_PP(16'h13075,4);
TASK_PP(16'h13076,4);
TASK_PP(16'h13077,4);
TASK_PP(16'h13078,4);
TASK_PP(16'h13079,4);
TASK_PP(16'h1307A,4);
TASK_PP(16'h1307B,4);
TASK_PP(16'h1307C,4);
TASK_PP(16'h1307D,4);
TASK_PP(16'h1307E,4);
TASK_PP(16'h1307F,4);
TASK_PP(16'h13080,4);
TASK_PP(16'h13081,4);
TASK_PP(16'h13082,4);
TASK_PP(16'h13083,4);
TASK_PP(16'h13084,4);
TASK_PP(16'h13085,4);
TASK_PP(16'h13086,4);
TASK_PP(16'h13087,4);
TASK_PP(16'h13088,4);
TASK_PP(16'h13089,4);
TASK_PP(16'h1308A,4);
TASK_PP(16'h1308B,4);
TASK_PP(16'h1308C,4);
TASK_PP(16'h1308D,4);
TASK_PP(16'h1308E,4);
TASK_PP(16'h1308F,4);
TASK_PP(16'h13090,4);
TASK_PP(16'h13091,4);
TASK_PP(16'h13092,4);
TASK_PP(16'h13093,4);
TASK_PP(16'h13094,4);
TASK_PP(16'h13095,4);
TASK_PP(16'h13096,4);
TASK_PP(16'h13097,4);
TASK_PP(16'h13098,4);
TASK_PP(16'h13099,4);
TASK_PP(16'h1309A,4);
TASK_PP(16'h1309B,4);
TASK_PP(16'h1309C,4);
TASK_PP(16'h1309D,4);
TASK_PP(16'h1309E,4);
TASK_PP(16'h1309F,4);
TASK_PP(16'h130A0,4);
TASK_PP(16'h130A1,4);
TASK_PP(16'h130A2,4);
TASK_PP(16'h130A3,4);
TASK_PP(16'h130A4,4);
TASK_PP(16'h130A5,4);
TASK_PP(16'h130A6,4);
TASK_PP(16'h130A7,4);
TASK_PP(16'h130A8,4);
TASK_PP(16'h130A9,4);
TASK_PP(16'h130AA,4);
TASK_PP(16'h130AB,4);
TASK_PP(16'h130AC,4);
TASK_PP(16'h130AD,4);
TASK_PP(16'h130AE,4);
TASK_PP(16'h130AF,4);
TASK_PP(16'h130B0,4);
TASK_PP(16'h130B1,4);
TASK_PP(16'h130B2,4);
TASK_PP(16'h130B3,4);
TASK_PP(16'h130B4,4);
TASK_PP(16'h130B5,4);
TASK_PP(16'h130B6,4);
TASK_PP(16'h130B7,4);
TASK_PP(16'h130B8,4);
TASK_PP(16'h130B9,4);
TASK_PP(16'h130BA,4);
TASK_PP(16'h130BB,4);
TASK_PP(16'h130BC,4);
TASK_PP(16'h130BD,4);
TASK_PP(16'h130BE,4);
TASK_PP(16'h130BF,4);
TASK_PP(16'h130C0,4);
TASK_PP(16'h130C1,4);
TASK_PP(16'h130C2,4);
TASK_PP(16'h130C3,4);
TASK_PP(16'h130C4,4);
TASK_PP(16'h130C5,4);
TASK_PP(16'h130C6,4);
TASK_PP(16'h130C7,4);
TASK_PP(16'h130C8,4);
TASK_PP(16'h130C9,4);
TASK_PP(16'h130CA,4);
TASK_PP(16'h130CB,4);
TASK_PP(16'h130CC,4);
TASK_PP(16'h130CD,4);
TASK_PP(16'h130CE,4);
TASK_PP(16'h130CF,4);
TASK_PP(16'h130D0,4);
TASK_PP(16'h130D1,4);
TASK_PP(16'h130D2,4);
TASK_PP(16'h130D3,4);
TASK_PP(16'h130D4,4);
TASK_PP(16'h130D5,4);
TASK_PP(16'h130D6,4);
TASK_PP(16'h130D7,4);
TASK_PP(16'h130D8,4);
TASK_PP(16'h130D9,4);
TASK_PP(16'h130DA,4);
TASK_PP(16'h130DB,4);
TASK_PP(16'h130DC,4);
TASK_PP(16'h130DD,4);
TASK_PP(16'h130DE,4);
TASK_PP(16'h130DF,4);
TASK_PP(16'h130E0,4);
TASK_PP(16'h130E1,4);
TASK_PP(16'h130E2,4);
TASK_PP(16'h130E3,4);
TASK_PP(16'h130E4,4);
TASK_PP(16'h130E5,4);
TASK_PP(16'h130E6,4);
TASK_PP(16'h130E7,4);
TASK_PP(16'h130E8,4);
TASK_PP(16'h130E9,4);
TASK_PP(16'h130EA,4);
TASK_PP(16'h130EB,4);
TASK_PP(16'h130EC,4);
TASK_PP(16'h130ED,4);
TASK_PP(16'h130EE,4);
TASK_PP(16'h130EF,4);
TASK_PP(16'h130F0,4);
TASK_PP(16'h130F1,4);
TASK_PP(16'h130F2,4);
TASK_PP(16'h130F3,4);
TASK_PP(16'h130F4,4);
TASK_PP(16'h130F5,4);
TASK_PP(16'h130F6,4);
TASK_PP(16'h130F7,4);
TASK_PP(16'h130F8,4);
TASK_PP(16'h130F9,4);
TASK_PP(16'h130FA,4);
TASK_PP(16'h130FB,4);
TASK_PP(16'h130FC,4);
TASK_PP(16'h130FD,4);
TASK_PP(16'h130FE,4);
TASK_PP(16'h130FF,4);
TASK_PP(16'h13100,4);
TASK_PP(16'h13101,4);
TASK_PP(16'h13102,4);
TASK_PP(16'h13103,4);
TASK_PP(16'h13104,4);
TASK_PP(16'h13105,4);
TASK_PP(16'h13106,4);
TASK_PP(16'h13107,4);
TASK_PP(16'h13108,4);
TASK_PP(16'h13109,4);
TASK_PP(16'h1310A,4);
TASK_PP(16'h1310B,4);
TASK_PP(16'h1310C,4);
TASK_PP(16'h1310D,4);
TASK_PP(16'h1310E,4);
TASK_PP(16'h1310F,4);
TASK_PP(16'h13110,4);
TASK_PP(16'h13111,4);
TASK_PP(16'h13112,4);
TASK_PP(16'h13113,4);
TASK_PP(16'h13114,4);
TASK_PP(16'h13115,4);
TASK_PP(16'h13116,4);
TASK_PP(16'h13117,4);
TASK_PP(16'h13118,4);
TASK_PP(16'h13119,4);
TASK_PP(16'h1311A,4);
TASK_PP(16'h1311B,4);
TASK_PP(16'h1311C,4);
TASK_PP(16'h1311D,4);
TASK_PP(16'h1311E,4);
TASK_PP(16'h1311F,4);
TASK_PP(16'h13120,4);
TASK_PP(16'h13121,4);
TASK_PP(16'h13122,4);
TASK_PP(16'h13123,4);
TASK_PP(16'h13124,4);
TASK_PP(16'h13125,4);
TASK_PP(16'h13126,4);
TASK_PP(16'h13127,4);
TASK_PP(16'h13128,4);
TASK_PP(16'h13129,4);
TASK_PP(16'h1312A,4);
TASK_PP(16'h1312B,4);
TASK_PP(16'h1312C,4);
TASK_PP(16'h1312D,4);
TASK_PP(16'h1312E,4);
TASK_PP(16'h1312F,4);
TASK_PP(16'h13130,4);
TASK_PP(16'h13131,4);
TASK_PP(16'h13132,4);
TASK_PP(16'h13133,4);
TASK_PP(16'h13134,4);
TASK_PP(16'h13135,4);
TASK_PP(16'h13136,4);
TASK_PP(16'h13137,4);
TASK_PP(16'h13138,4);
TASK_PP(16'h13139,4);
TASK_PP(16'h1313A,4);
TASK_PP(16'h1313B,4);
TASK_PP(16'h1313C,4);
TASK_PP(16'h1313D,4);
TASK_PP(16'h1313E,4);
TASK_PP(16'h1313F,4);
TASK_PP(16'h13140,4);
TASK_PP(16'h13141,4);
TASK_PP(16'h13142,4);
TASK_PP(16'h13143,4);
TASK_PP(16'h13144,4);
TASK_PP(16'h13145,4);
TASK_PP(16'h13146,4);
TASK_PP(16'h13147,4);
TASK_PP(16'h13148,4);
TASK_PP(16'h13149,4);
TASK_PP(16'h1314A,4);
TASK_PP(16'h1314B,4);
TASK_PP(16'h1314C,4);
TASK_PP(16'h1314D,4);
TASK_PP(16'h1314E,4);
TASK_PP(16'h1314F,4);
TASK_PP(16'h13150,4);
TASK_PP(16'h13151,4);
TASK_PP(16'h13152,4);
TASK_PP(16'h13153,4);
TASK_PP(16'h13154,4);
TASK_PP(16'h13155,4);
TASK_PP(16'h13156,4);
TASK_PP(16'h13157,4);
TASK_PP(16'h13158,4);
TASK_PP(16'h13159,4);
TASK_PP(16'h1315A,4);
TASK_PP(16'h1315B,4);
TASK_PP(16'h1315C,4);
TASK_PP(16'h1315D,4);
TASK_PP(16'h1315E,4);
TASK_PP(16'h1315F,4);
TASK_PP(16'h13160,4);
TASK_PP(16'h13161,4);
TASK_PP(16'h13162,4);
TASK_PP(16'h13163,4);
TASK_PP(16'h13164,4);
TASK_PP(16'h13165,4);
TASK_PP(16'h13166,4);
TASK_PP(16'h13167,4);
TASK_PP(16'h13168,4);
TASK_PP(16'h13169,4);
TASK_PP(16'h1316A,4);
TASK_PP(16'h1316B,4);
TASK_PP(16'h1316C,4);
TASK_PP(16'h1316D,4);
TASK_PP(16'h1316E,4);
TASK_PP(16'h1316F,4);
TASK_PP(16'h13170,4);
TASK_PP(16'h13171,4);
TASK_PP(16'h13172,4);
TASK_PP(16'h13173,4);
TASK_PP(16'h13174,4);
TASK_PP(16'h13175,4);
TASK_PP(16'h13176,4);
TASK_PP(16'h13177,4);
TASK_PP(16'h13178,4);
TASK_PP(16'h13179,4);
TASK_PP(16'h1317A,4);
TASK_PP(16'h1317B,4);
TASK_PP(16'h1317C,4);
TASK_PP(16'h1317D,4);
TASK_PP(16'h1317E,4);
TASK_PP(16'h1317F,4);
TASK_PP(16'h13180,4);
TASK_PP(16'h13181,4);
TASK_PP(16'h13182,4);
TASK_PP(16'h13183,4);
TASK_PP(16'h13184,4);
TASK_PP(16'h13185,4);
TASK_PP(16'h13186,4);
TASK_PP(16'h13187,4);
TASK_PP(16'h13188,4);
TASK_PP(16'h13189,4);
TASK_PP(16'h1318A,4);
TASK_PP(16'h1318B,4);
TASK_PP(16'h1318C,4);
TASK_PP(16'h1318D,4);
TASK_PP(16'h1318E,4);
TASK_PP(16'h1318F,4);
TASK_PP(16'h13190,4);
TASK_PP(16'h13191,4);
TASK_PP(16'h13192,4);
TASK_PP(16'h13193,4);
TASK_PP(16'h13194,4);
TASK_PP(16'h13195,4);
TASK_PP(16'h13196,4);
TASK_PP(16'h13197,4);
TASK_PP(16'h13198,4);
TASK_PP(16'h13199,4);
TASK_PP(16'h1319A,4);
TASK_PP(16'h1319B,4);
TASK_PP(16'h1319C,4);
TASK_PP(16'h1319D,4);
TASK_PP(16'h1319E,4);
TASK_PP(16'h1319F,4);
TASK_PP(16'h131A0,4);
TASK_PP(16'h131A1,4);
TASK_PP(16'h131A2,4);
TASK_PP(16'h131A3,4);
TASK_PP(16'h131A4,4);
TASK_PP(16'h131A5,4);
TASK_PP(16'h131A6,4);
TASK_PP(16'h131A7,4);
TASK_PP(16'h131A8,4);
TASK_PP(16'h131A9,4);
TASK_PP(16'h131AA,4);
TASK_PP(16'h131AB,4);
TASK_PP(16'h131AC,4);
TASK_PP(16'h131AD,4);
TASK_PP(16'h131AE,4);
TASK_PP(16'h131AF,4);
TASK_PP(16'h131B0,4);
TASK_PP(16'h131B1,4);
TASK_PP(16'h131B2,4);
TASK_PP(16'h131B3,4);
TASK_PP(16'h131B4,4);
TASK_PP(16'h131B5,4);
TASK_PP(16'h131B6,4);
TASK_PP(16'h131B7,4);
TASK_PP(16'h131B8,4);
TASK_PP(16'h131B9,4);
TASK_PP(16'h131BA,4);
TASK_PP(16'h131BB,4);
TASK_PP(16'h131BC,4);
TASK_PP(16'h131BD,4);
TASK_PP(16'h131BE,4);
TASK_PP(16'h131BF,4);
TASK_PP(16'h131C0,4);
TASK_PP(16'h131C1,4);
TASK_PP(16'h131C2,4);
TASK_PP(16'h131C3,4);
TASK_PP(16'h131C4,4);
TASK_PP(16'h131C5,4);
TASK_PP(16'h131C6,4);
TASK_PP(16'h131C7,4);
TASK_PP(16'h131C8,4);
TASK_PP(16'h131C9,4);
TASK_PP(16'h131CA,4);
TASK_PP(16'h131CB,4);
TASK_PP(16'h131CC,4);
TASK_PP(16'h131CD,4);
TASK_PP(16'h131CE,4);
TASK_PP(16'h131CF,4);
TASK_PP(16'h131D0,4);
TASK_PP(16'h131D1,4);
TASK_PP(16'h131D2,4);
TASK_PP(16'h131D3,4);
TASK_PP(16'h131D4,4);
TASK_PP(16'h131D5,4);
TASK_PP(16'h131D6,4);
TASK_PP(16'h131D7,4);
TASK_PP(16'h131D8,4);
TASK_PP(16'h131D9,4);
TASK_PP(16'h131DA,4);
TASK_PP(16'h131DB,4);
TASK_PP(16'h131DC,4);
TASK_PP(16'h131DD,4);
TASK_PP(16'h131DE,4);
TASK_PP(16'h131DF,4);
TASK_PP(16'h131E0,4);
TASK_PP(16'h131E1,4);
TASK_PP(16'h131E2,4);
TASK_PP(16'h131E3,4);
TASK_PP(16'h131E4,4);
TASK_PP(16'h131E5,4);
TASK_PP(16'h131E6,4);
TASK_PP(16'h131E7,4);
TASK_PP(16'h131E8,4);
TASK_PP(16'h131E9,4);
TASK_PP(16'h131EA,4);
TASK_PP(16'h131EB,4);
TASK_PP(16'h131EC,4);
TASK_PP(16'h131ED,4);
TASK_PP(16'h131EE,4);
TASK_PP(16'h131EF,4);
TASK_PP(16'h131F0,4);
TASK_PP(16'h131F1,4);
TASK_PP(16'h131F2,4);
TASK_PP(16'h131F3,4);
TASK_PP(16'h131F4,4);
TASK_PP(16'h131F5,4);
TASK_PP(16'h131F6,4);
TASK_PP(16'h131F7,4);
TASK_PP(16'h131F8,4);
TASK_PP(16'h131F9,4);
TASK_PP(16'h131FA,4);
TASK_PP(16'h131FB,4);
TASK_PP(16'h131FC,4);
TASK_PP(16'h131FD,4);
TASK_PP(16'h131FE,4);
TASK_PP(16'h131FF,4);
TASK_PP(16'h13200,4);
TASK_PP(16'h13201,4);
TASK_PP(16'h13202,4);
TASK_PP(16'h13203,4);
TASK_PP(16'h13204,4);
TASK_PP(16'h13205,4);
TASK_PP(16'h13206,4);
TASK_PP(16'h13207,4);
TASK_PP(16'h13208,4);
TASK_PP(16'h13209,4);
TASK_PP(16'h1320A,4);
TASK_PP(16'h1320B,4);
TASK_PP(16'h1320C,4);
TASK_PP(16'h1320D,4);
TASK_PP(16'h1320E,4);
TASK_PP(16'h1320F,4);
TASK_PP(16'h13210,4);
TASK_PP(16'h13211,4);
TASK_PP(16'h13212,4);
TASK_PP(16'h13213,4);
TASK_PP(16'h13214,4);
TASK_PP(16'h13215,4);
TASK_PP(16'h13216,4);
TASK_PP(16'h13217,4);
TASK_PP(16'h13218,4);
TASK_PP(16'h13219,4);
TASK_PP(16'h1321A,4);
TASK_PP(16'h1321B,4);
TASK_PP(16'h1321C,4);
TASK_PP(16'h1321D,4);
TASK_PP(16'h1321E,4);
TASK_PP(16'h1321F,4);
TASK_PP(16'h13220,4);
TASK_PP(16'h13221,4);
TASK_PP(16'h13222,4);
TASK_PP(16'h13223,4);
TASK_PP(16'h13224,4);
TASK_PP(16'h13225,4);
TASK_PP(16'h13226,4);
TASK_PP(16'h13227,4);
TASK_PP(16'h13228,4);
TASK_PP(16'h13229,4);
TASK_PP(16'h1322A,4);
TASK_PP(16'h1322B,4);
TASK_PP(16'h1322C,4);
TASK_PP(16'h1322D,4);
TASK_PP(16'h1322E,4);
TASK_PP(16'h1322F,4);
TASK_PP(16'h13230,4);
TASK_PP(16'h13231,4);
TASK_PP(16'h13232,4);
TASK_PP(16'h13233,4);
TASK_PP(16'h13234,4);
TASK_PP(16'h13235,4);
TASK_PP(16'h13236,4);
TASK_PP(16'h13237,4);
TASK_PP(16'h13238,4);
TASK_PP(16'h13239,4);
TASK_PP(16'h1323A,4);
TASK_PP(16'h1323B,4);
TASK_PP(16'h1323C,4);
TASK_PP(16'h1323D,4);
TASK_PP(16'h1323E,4);
TASK_PP(16'h1323F,4);
TASK_PP(16'h13240,4);
TASK_PP(16'h13241,4);
TASK_PP(16'h13242,4);
TASK_PP(16'h13243,4);
TASK_PP(16'h13244,4);
TASK_PP(16'h13245,4);
TASK_PP(16'h13246,4);
TASK_PP(16'h13247,4);
TASK_PP(16'h13248,4);
TASK_PP(16'h13249,4);
TASK_PP(16'h1324A,4);
TASK_PP(16'h1324B,4);
TASK_PP(16'h1324C,4);
TASK_PP(16'h1324D,4);
TASK_PP(16'h1324E,4);
TASK_PP(16'h1324F,4);
TASK_PP(16'h13250,4);
TASK_PP(16'h13251,4);
TASK_PP(16'h13252,4);
TASK_PP(16'h13253,4);
TASK_PP(16'h13254,4);
TASK_PP(16'h13255,4);
TASK_PP(16'h13256,4);
TASK_PP(16'h13257,4);
TASK_PP(16'h13258,4);
TASK_PP(16'h13259,4);
TASK_PP(16'h1325A,4);
TASK_PP(16'h1325B,4);
TASK_PP(16'h1325C,4);
TASK_PP(16'h1325D,4);
TASK_PP(16'h1325E,4);
TASK_PP(16'h1325F,4);
TASK_PP(16'h13260,4);
TASK_PP(16'h13261,4);
TASK_PP(16'h13262,4);
TASK_PP(16'h13263,4);
TASK_PP(16'h13264,4);
TASK_PP(16'h13265,4);
TASK_PP(16'h13266,4);
TASK_PP(16'h13267,4);
TASK_PP(16'h13268,4);
TASK_PP(16'h13269,4);
TASK_PP(16'h1326A,4);
TASK_PP(16'h1326B,4);
TASK_PP(16'h1326C,4);
TASK_PP(16'h1326D,4);
TASK_PP(16'h1326E,4);
TASK_PP(16'h1326F,4);
TASK_PP(16'h13270,4);
TASK_PP(16'h13271,4);
TASK_PP(16'h13272,4);
TASK_PP(16'h13273,4);
TASK_PP(16'h13274,4);
TASK_PP(16'h13275,4);
TASK_PP(16'h13276,4);
TASK_PP(16'h13277,4);
TASK_PP(16'h13278,4);
TASK_PP(16'h13279,4);
TASK_PP(16'h1327A,4);
TASK_PP(16'h1327B,4);
TASK_PP(16'h1327C,4);
TASK_PP(16'h1327D,4);
TASK_PP(16'h1327E,4);
TASK_PP(16'h1327F,4);
TASK_PP(16'h13280,4);
TASK_PP(16'h13281,4);
TASK_PP(16'h13282,4);
TASK_PP(16'h13283,4);
TASK_PP(16'h13284,4);
TASK_PP(16'h13285,4);
TASK_PP(16'h13286,4);
TASK_PP(16'h13287,4);
TASK_PP(16'h13288,4);
TASK_PP(16'h13289,4);
TASK_PP(16'h1328A,4);
TASK_PP(16'h1328B,4);
TASK_PP(16'h1328C,4);
TASK_PP(16'h1328D,4);
TASK_PP(16'h1328E,4);
TASK_PP(16'h1328F,4);
TASK_PP(16'h13290,4);
TASK_PP(16'h13291,4);
TASK_PP(16'h13292,4);
TASK_PP(16'h13293,4);
TASK_PP(16'h13294,4);
TASK_PP(16'h13295,4);
TASK_PP(16'h13296,4);
TASK_PP(16'h13297,4);
TASK_PP(16'h13298,4);
TASK_PP(16'h13299,4);
TASK_PP(16'h1329A,4);
TASK_PP(16'h1329B,4);
TASK_PP(16'h1329C,4);
TASK_PP(16'h1329D,4);
TASK_PP(16'h1329E,4);
TASK_PP(16'h1329F,4);
TASK_PP(16'h132A0,4);
TASK_PP(16'h132A1,4);
TASK_PP(16'h132A2,4);
TASK_PP(16'h132A3,4);
TASK_PP(16'h132A4,4);
TASK_PP(16'h132A5,4);
TASK_PP(16'h132A6,4);
TASK_PP(16'h132A7,4);
TASK_PP(16'h132A8,4);
TASK_PP(16'h132A9,4);
TASK_PP(16'h132AA,4);
TASK_PP(16'h132AB,4);
TASK_PP(16'h132AC,4);
TASK_PP(16'h132AD,4);
TASK_PP(16'h132AE,4);
TASK_PP(16'h132AF,4);
TASK_PP(16'h132B0,4);
TASK_PP(16'h132B1,4);
TASK_PP(16'h132B2,4);
TASK_PP(16'h132B3,4);
TASK_PP(16'h132B4,4);
TASK_PP(16'h132B5,4);
TASK_PP(16'h132B6,4);
TASK_PP(16'h132B7,4);
TASK_PP(16'h132B8,4);
TASK_PP(16'h132B9,4);
TASK_PP(16'h132BA,4);
TASK_PP(16'h132BB,4);
TASK_PP(16'h132BC,4);
TASK_PP(16'h132BD,4);
TASK_PP(16'h132BE,4);
TASK_PP(16'h132BF,4);
TASK_PP(16'h132C0,4);
TASK_PP(16'h132C1,4);
TASK_PP(16'h132C2,4);
TASK_PP(16'h132C3,4);
TASK_PP(16'h132C4,4);
TASK_PP(16'h132C5,4);
TASK_PP(16'h132C6,4);
TASK_PP(16'h132C7,4);
TASK_PP(16'h132C8,4);
TASK_PP(16'h132C9,4);
TASK_PP(16'h132CA,4);
TASK_PP(16'h132CB,4);
TASK_PP(16'h132CC,4);
TASK_PP(16'h132CD,4);
TASK_PP(16'h132CE,4);
TASK_PP(16'h132CF,4);
TASK_PP(16'h132D0,4);
TASK_PP(16'h132D1,4);
TASK_PP(16'h132D2,4);
TASK_PP(16'h132D3,4);
TASK_PP(16'h132D4,4);
TASK_PP(16'h132D5,4);
TASK_PP(16'h132D6,4);
TASK_PP(16'h132D7,4);
TASK_PP(16'h132D8,4);
TASK_PP(16'h132D9,4);
TASK_PP(16'h132DA,4);
TASK_PP(16'h132DB,4);
TASK_PP(16'h132DC,4);
TASK_PP(16'h132DD,4);
TASK_PP(16'h132DE,4);
TASK_PP(16'h132DF,4);
TASK_PP(16'h132E0,4);
TASK_PP(16'h132E1,4);
TASK_PP(16'h132E2,4);
TASK_PP(16'h132E3,4);
TASK_PP(16'h132E4,4);
TASK_PP(16'h132E5,4);
TASK_PP(16'h132E6,4);
TASK_PP(16'h132E7,4);
TASK_PP(16'h132E8,4);
TASK_PP(16'h132E9,4);
TASK_PP(16'h132EA,4);
TASK_PP(16'h132EB,4);
TASK_PP(16'h132EC,4);
TASK_PP(16'h132ED,4);
TASK_PP(16'h132EE,4);
TASK_PP(16'h132EF,4);
TASK_PP(16'h132F0,4);
TASK_PP(16'h132F1,4);
TASK_PP(16'h132F2,4);
TASK_PP(16'h132F3,4);
TASK_PP(16'h132F4,4);
TASK_PP(16'h132F5,4);
TASK_PP(16'h132F6,4);
TASK_PP(16'h132F7,4);
TASK_PP(16'h132F8,4);
TASK_PP(16'h132F9,4);
TASK_PP(16'h132FA,4);
TASK_PP(16'h132FB,4);
TASK_PP(16'h132FC,4);
TASK_PP(16'h132FD,4);
TASK_PP(16'h132FE,4);
TASK_PP(16'h132FF,4);
TASK_PP(16'h13300,4);
TASK_PP(16'h13301,4);
TASK_PP(16'h13302,4);
TASK_PP(16'h13303,4);
TASK_PP(16'h13304,4);
TASK_PP(16'h13305,4);
TASK_PP(16'h13306,4);
TASK_PP(16'h13307,4);
TASK_PP(16'h13308,4);
TASK_PP(16'h13309,4);
TASK_PP(16'h1330A,4);
TASK_PP(16'h1330B,4);
TASK_PP(16'h1330C,4);
TASK_PP(16'h1330D,4);
TASK_PP(16'h1330E,4);
TASK_PP(16'h1330F,4);
TASK_PP(16'h13310,4);
TASK_PP(16'h13311,4);
TASK_PP(16'h13312,4);
TASK_PP(16'h13313,4);
TASK_PP(16'h13314,4);
TASK_PP(16'h13315,4);
TASK_PP(16'h13316,4);
TASK_PP(16'h13317,4);
TASK_PP(16'h13318,4);
TASK_PP(16'h13319,4);
TASK_PP(16'h1331A,4);
TASK_PP(16'h1331B,4);
TASK_PP(16'h1331C,4);
TASK_PP(16'h1331D,4);
TASK_PP(16'h1331E,4);
TASK_PP(16'h1331F,4);
TASK_PP(16'h13320,4);
TASK_PP(16'h13321,4);
TASK_PP(16'h13322,4);
TASK_PP(16'h13323,4);
TASK_PP(16'h13324,4);
TASK_PP(16'h13325,4);
TASK_PP(16'h13326,4);
TASK_PP(16'h13327,4);
TASK_PP(16'h13328,4);
TASK_PP(16'h13329,4);
TASK_PP(16'h1332A,4);
TASK_PP(16'h1332B,4);
TASK_PP(16'h1332C,4);
TASK_PP(16'h1332D,4);
TASK_PP(16'h1332E,4);
TASK_PP(16'h1332F,4);
TASK_PP(16'h13330,4);
TASK_PP(16'h13331,4);
TASK_PP(16'h13332,4);
TASK_PP(16'h13333,4);
TASK_PP(16'h13334,4);
TASK_PP(16'h13335,4);
TASK_PP(16'h13336,4);
TASK_PP(16'h13337,4);
TASK_PP(16'h13338,4);
TASK_PP(16'h13339,4);
TASK_PP(16'h1333A,4);
TASK_PP(16'h1333B,4);
TASK_PP(16'h1333C,4);
TASK_PP(16'h1333D,4);
TASK_PP(16'h1333E,4);
TASK_PP(16'h1333F,4);
TASK_PP(16'h13340,4);
TASK_PP(16'h13341,4);
TASK_PP(16'h13342,4);
TASK_PP(16'h13343,4);
TASK_PP(16'h13344,4);
TASK_PP(16'h13345,4);
TASK_PP(16'h13346,4);
TASK_PP(16'h13347,4);
TASK_PP(16'h13348,4);
TASK_PP(16'h13349,4);
TASK_PP(16'h1334A,4);
TASK_PP(16'h1334B,4);
TASK_PP(16'h1334C,4);
TASK_PP(16'h1334D,4);
TASK_PP(16'h1334E,4);
TASK_PP(16'h1334F,4);
TASK_PP(16'h13350,4);
TASK_PP(16'h13351,4);
TASK_PP(16'h13352,4);
TASK_PP(16'h13353,4);
TASK_PP(16'h13354,4);
TASK_PP(16'h13355,4);
TASK_PP(16'h13356,4);
TASK_PP(16'h13357,4);
TASK_PP(16'h13358,4);
TASK_PP(16'h13359,4);
TASK_PP(16'h1335A,4);
TASK_PP(16'h1335B,4);
TASK_PP(16'h1335C,4);
TASK_PP(16'h1335D,4);
TASK_PP(16'h1335E,4);
TASK_PP(16'h1335F,4);
TASK_PP(16'h13360,4);
TASK_PP(16'h13361,4);
TASK_PP(16'h13362,4);
TASK_PP(16'h13363,4);
TASK_PP(16'h13364,4);
TASK_PP(16'h13365,4);
TASK_PP(16'h13366,4);
TASK_PP(16'h13367,4);
TASK_PP(16'h13368,4);
TASK_PP(16'h13369,4);
TASK_PP(16'h1336A,4);
TASK_PP(16'h1336B,4);
TASK_PP(16'h1336C,4);
TASK_PP(16'h1336D,4);
TASK_PP(16'h1336E,4);
TASK_PP(16'h1336F,4);
TASK_PP(16'h13370,4);
TASK_PP(16'h13371,4);
TASK_PP(16'h13372,4);
TASK_PP(16'h13373,4);
TASK_PP(16'h13374,4);
TASK_PP(16'h13375,4);
TASK_PP(16'h13376,4);
TASK_PP(16'h13377,4);
TASK_PP(16'h13378,4);
TASK_PP(16'h13379,4);
TASK_PP(16'h1337A,4);
TASK_PP(16'h1337B,4);
TASK_PP(16'h1337C,4);
TASK_PP(16'h1337D,4);
TASK_PP(16'h1337E,4);
TASK_PP(16'h1337F,4);
TASK_PP(16'h13380,4);
TASK_PP(16'h13381,4);
TASK_PP(16'h13382,4);
TASK_PP(16'h13383,4);
TASK_PP(16'h13384,4);
TASK_PP(16'h13385,4);
TASK_PP(16'h13386,4);
TASK_PP(16'h13387,4);
TASK_PP(16'h13388,4);
TASK_PP(16'h13389,4);
TASK_PP(16'h1338A,4);
TASK_PP(16'h1338B,4);
TASK_PP(16'h1338C,4);
TASK_PP(16'h1338D,4);
TASK_PP(16'h1338E,4);
TASK_PP(16'h1338F,4);
TASK_PP(16'h13390,4);
TASK_PP(16'h13391,4);
TASK_PP(16'h13392,4);
TASK_PP(16'h13393,4);
TASK_PP(16'h13394,4);
TASK_PP(16'h13395,4);
TASK_PP(16'h13396,4);
TASK_PP(16'h13397,4);
TASK_PP(16'h13398,4);
TASK_PP(16'h13399,4);
TASK_PP(16'h1339A,4);
TASK_PP(16'h1339B,4);
TASK_PP(16'h1339C,4);
TASK_PP(16'h1339D,4);
TASK_PP(16'h1339E,4);
TASK_PP(16'h1339F,4);
TASK_PP(16'h133A0,4);
TASK_PP(16'h133A1,4);
TASK_PP(16'h133A2,4);
TASK_PP(16'h133A3,4);
TASK_PP(16'h133A4,4);
TASK_PP(16'h133A5,4);
TASK_PP(16'h133A6,4);
TASK_PP(16'h133A7,4);
TASK_PP(16'h133A8,4);
TASK_PP(16'h133A9,4);
TASK_PP(16'h133AA,4);
TASK_PP(16'h133AB,4);
TASK_PP(16'h133AC,4);
TASK_PP(16'h133AD,4);
TASK_PP(16'h133AE,4);
TASK_PP(16'h133AF,4);
TASK_PP(16'h133B0,4);
TASK_PP(16'h133B1,4);
TASK_PP(16'h133B2,4);
TASK_PP(16'h133B3,4);
TASK_PP(16'h133B4,4);
TASK_PP(16'h133B5,4);
TASK_PP(16'h133B6,4);
TASK_PP(16'h133B7,4);
TASK_PP(16'h133B8,4);
TASK_PP(16'h133B9,4);
TASK_PP(16'h133BA,4);
TASK_PP(16'h133BB,4);
TASK_PP(16'h133BC,4);
TASK_PP(16'h133BD,4);
TASK_PP(16'h133BE,4);
TASK_PP(16'h133BF,4);
TASK_PP(16'h133C0,4);
TASK_PP(16'h133C1,4);
TASK_PP(16'h133C2,4);
TASK_PP(16'h133C3,4);
TASK_PP(16'h133C4,4);
TASK_PP(16'h133C5,4);
TASK_PP(16'h133C6,4);
TASK_PP(16'h133C7,4);
TASK_PP(16'h133C8,4);
TASK_PP(16'h133C9,4);
TASK_PP(16'h133CA,4);
TASK_PP(16'h133CB,4);
TASK_PP(16'h133CC,4);
TASK_PP(16'h133CD,4);
TASK_PP(16'h133CE,4);
TASK_PP(16'h133CF,4);
TASK_PP(16'h133D0,4);
TASK_PP(16'h133D1,4);
TASK_PP(16'h133D2,4);
TASK_PP(16'h133D3,4);
TASK_PP(16'h133D4,4);
TASK_PP(16'h133D5,4);
TASK_PP(16'h133D6,4);
TASK_PP(16'h133D7,4);
TASK_PP(16'h133D8,4);
TASK_PP(16'h133D9,4);
TASK_PP(16'h133DA,4);
TASK_PP(16'h133DB,4);
TASK_PP(16'h133DC,4);
TASK_PP(16'h133DD,4);
TASK_PP(16'h133DE,4);
TASK_PP(16'h133DF,4);
TASK_PP(16'h133E0,4);
TASK_PP(16'h133E1,4);
TASK_PP(16'h133E2,4);
TASK_PP(16'h133E3,4);
TASK_PP(16'h133E4,4);
TASK_PP(16'h133E5,4);
TASK_PP(16'h133E6,4);
TASK_PP(16'h133E7,4);
TASK_PP(16'h133E8,4);
TASK_PP(16'h133E9,4);
TASK_PP(16'h133EA,4);
TASK_PP(16'h133EB,4);
TASK_PP(16'h133EC,4);
TASK_PP(16'h133ED,4);
TASK_PP(16'h133EE,4);
TASK_PP(16'h133EF,4);
TASK_PP(16'h133F0,4);
TASK_PP(16'h133F1,4);
TASK_PP(16'h133F2,4);
TASK_PP(16'h133F3,4);
TASK_PP(16'h133F4,4);
TASK_PP(16'h133F5,4);
TASK_PP(16'h133F6,4);
TASK_PP(16'h133F7,4);
TASK_PP(16'h133F8,4);
TASK_PP(16'h133F9,4);
TASK_PP(16'h133FA,4);
TASK_PP(16'h133FB,4);
TASK_PP(16'h133FC,4);
TASK_PP(16'h133FD,4);
TASK_PP(16'h133FE,4);
TASK_PP(16'h133FF,4);
TASK_PP(16'h13400,4);
TASK_PP(16'h13401,4);
TASK_PP(16'h13402,4);
TASK_PP(16'h13403,4);
TASK_PP(16'h13404,4);
TASK_PP(16'h13405,4);
TASK_PP(16'h13406,4);
TASK_PP(16'h13407,4);
TASK_PP(16'h13408,4);
TASK_PP(16'h13409,4);
TASK_PP(16'h1340A,4);
TASK_PP(16'h1340B,4);
TASK_PP(16'h1340C,4);
TASK_PP(16'h1340D,4);
TASK_PP(16'h1340E,4);
TASK_PP(16'h1340F,4);
TASK_PP(16'h13410,4);
TASK_PP(16'h13411,4);
TASK_PP(16'h13412,4);
TASK_PP(16'h13413,4);
TASK_PP(16'h13414,4);
TASK_PP(16'h13415,4);
TASK_PP(16'h13416,4);
TASK_PP(16'h13417,4);
TASK_PP(16'h13418,4);
TASK_PP(16'h13419,4);
TASK_PP(16'h1341A,4);
TASK_PP(16'h1341B,4);
TASK_PP(16'h1341C,4);
TASK_PP(16'h1341D,4);
TASK_PP(16'h1341E,4);
TASK_PP(16'h1341F,4);
TASK_PP(16'h13420,4);
TASK_PP(16'h13421,4);
TASK_PP(16'h13422,4);
TASK_PP(16'h13423,4);
TASK_PP(16'h13424,4);
TASK_PP(16'h13425,4);
TASK_PP(16'h13426,4);
TASK_PP(16'h13427,4);
TASK_PP(16'h13428,4);
TASK_PP(16'h13429,4);
TASK_PP(16'h1342A,4);
TASK_PP(16'h1342B,4);
TASK_PP(16'h1342C,4);
TASK_PP(16'h1342D,4);
TASK_PP(16'h1342E,4);
TASK_PP(16'h1342F,4);
TASK_PP(16'h13430,4);
TASK_PP(16'h13431,4);
TASK_PP(16'h13432,4);
TASK_PP(16'h13433,4);
TASK_PP(16'h13434,4);
TASK_PP(16'h13435,4);
TASK_PP(16'h13436,4);
TASK_PP(16'h13437,4);
TASK_PP(16'h13438,4);
TASK_PP(16'h13439,4);
TASK_PP(16'h1343A,4);
TASK_PP(16'h1343B,4);
TASK_PP(16'h1343C,4);
TASK_PP(16'h1343D,4);
TASK_PP(16'h1343E,4);
TASK_PP(16'h1343F,4);
TASK_PP(16'h13440,4);
TASK_PP(16'h13441,4);
TASK_PP(16'h13442,4);
TASK_PP(16'h13443,4);
TASK_PP(16'h13444,4);
TASK_PP(16'h13445,4);
TASK_PP(16'h13446,4);
TASK_PP(16'h13447,4);
TASK_PP(16'h13448,4);
TASK_PP(16'h13449,4);
TASK_PP(16'h1344A,4);
TASK_PP(16'h1344B,4);
TASK_PP(16'h1344C,4);
TASK_PP(16'h1344D,4);
TASK_PP(16'h1344E,4);
TASK_PP(16'h1344F,4);
TASK_PP(16'h13450,4);
TASK_PP(16'h13451,4);
TASK_PP(16'h13452,4);
TASK_PP(16'h13453,4);
TASK_PP(16'h13454,4);
TASK_PP(16'h13455,4);
TASK_PP(16'h13456,4);
TASK_PP(16'h13457,4);
TASK_PP(16'h13458,4);
TASK_PP(16'h13459,4);
TASK_PP(16'h1345A,4);
TASK_PP(16'h1345B,4);
TASK_PP(16'h1345C,4);
TASK_PP(16'h1345D,4);
TASK_PP(16'h1345E,4);
TASK_PP(16'h1345F,4);
TASK_PP(16'h13460,4);
TASK_PP(16'h13461,4);
TASK_PP(16'h13462,4);
TASK_PP(16'h13463,4);
TASK_PP(16'h13464,4);
TASK_PP(16'h13465,4);
TASK_PP(16'h13466,4);
TASK_PP(16'h13467,4);
TASK_PP(16'h13468,4);
TASK_PP(16'h13469,4);
TASK_PP(16'h1346A,4);
TASK_PP(16'h1346B,4);
TASK_PP(16'h1346C,4);
TASK_PP(16'h1346D,4);
TASK_PP(16'h1346E,4);
TASK_PP(16'h1346F,4);
TASK_PP(16'h13470,4);
TASK_PP(16'h13471,4);
TASK_PP(16'h13472,4);
TASK_PP(16'h13473,4);
TASK_PP(16'h13474,4);
TASK_PP(16'h13475,4);
TASK_PP(16'h13476,4);
TASK_PP(16'h13477,4);
TASK_PP(16'h13478,4);
TASK_PP(16'h13479,4);
TASK_PP(16'h1347A,4);
TASK_PP(16'h1347B,4);
TASK_PP(16'h1347C,4);
TASK_PP(16'h1347D,4);
TASK_PP(16'h1347E,4);
TASK_PP(16'h1347F,4);
TASK_PP(16'h13480,4);
TASK_PP(16'h13481,4);
TASK_PP(16'h13482,4);
TASK_PP(16'h13483,4);
TASK_PP(16'h13484,4);
TASK_PP(16'h13485,4);
TASK_PP(16'h13486,4);
TASK_PP(16'h13487,4);
TASK_PP(16'h13488,4);
TASK_PP(16'h13489,4);
TASK_PP(16'h1348A,4);
TASK_PP(16'h1348B,4);
TASK_PP(16'h1348C,4);
TASK_PP(16'h1348D,4);
TASK_PP(16'h1348E,4);
TASK_PP(16'h1348F,4);
TASK_PP(16'h13490,4);
TASK_PP(16'h13491,4);
TASK_PP(16'h13492,4);
TASK_PP(16'h13493,4);
TASK_PP(16'h13494,4);
TASK_PP(16'h13495,4);
TASK_PP(16'h13496,4);
TASK_PP(16'h13497,4);
TASK_PP(16'h13498,4);
TASK_PP(16'h13499,4);
TASK_PP(16'h1349A,4);
TASK_PP(16'h1349B,4);
TASK_PP(16'h1349C,4);
TASK_PP(16'h1349D,4);
TASK_PP(16'h1349E,4);
TASK_PP(16'h1349F,4);
TASK_PP(16'h134A0,4);
TASK_PP(16'h134A1,4);
TASK_PP(16'h134A2,4);
TASK_PP(16'h134A3,4);
TASK_PP(16'h134A4,4);
TASK_PP(16'h134A5,4);
TASK_PP(16'h134A6,4);
TASK_PP(16'h134A7,4);
TASK_PP(16'h134A8,4);
TASK_PP(16'h134A9,4);
TASK_PP(16'h134AA,4);
TASK_PP(16'h134AB,4);
TASK_PP(16'h134AC,4);
TASK_PP(16'h134AD,4);
TASK_PP(16'h134AE,4);
TASK_PP(16'h134AF,4);
TASK_PP(16'h134B0,4);
TASK_PP(16'h134B1,4);
TASK_PP(16'h134B2,4);
TASK_PP(16'h134B3,4);
TASK_PP(16'h134B4,4);
TASK_PP(16'h134B5,4);
TASK_PP(16'h134B6,4);
TASK_PP(16'h134B7,4);
TASK_PP(16'h134B8,4);
TASK_PP(16'h134B9,4);
TASK_PP(16'h134BA,4);
TASK_PP(16'h134BB,4);
TASK_PP(16'h134BC,4);
TASK_PP(16'h134BD,4);
TASK_PP(16'h134BE,4);
TASK_PP(16'h134BF,4);
TASK_PP(16'h134C0,4);
TASK_PP(16'h134C1,4);
TASK_PP(16'h134C2,4);
TASK_PP(16'h134C3,4);
TASK_PP(16'h134C4,4);
TASK_PP(16'h134C5,4);
TASK_PP(16'h134C6,4);
TASK_PP(16'h134C7,4);
TASK_PP(16'h134C8,4);
TASK_PP(16'h134C9,4);
TASK_PP(16'h134CA,4);
TASK_PP(16'h134CB,4);
TASK_PP(16'h134CC,4);
TASK_PP(16'h134CD,4);
TASK_PP(16'h134CE,4);
TASK_PP(16'h134CF,4);
TASK_PP(16'h134D0,4);
TASK_PP(16'h134D1,4);
TASK_PP(16'h134D2,4);
TASK_PP(16'h134D3,4);
TASK_PP(16'h134D4,4);
TASK_PP(16'h134D5,4);
TASK_PP(16'h134D6,4);
TASK_PP(16'h134D7,4);
TASK_PP(16'h134D8,4);
TASK_PP(16'h134D9,4);
TASK_PP(16'h134DA,4);
TASK_PP(16'h134DB,4);
TASK_PP(16'h134DC,4);
TASK_PP(16'h134DD,4);
TASK_PP(16'h134DE,4);
TASK_PP(16'h134DF,4);
TASK_PP(16'h134E0,4);
TASK_PP(16'h134E1,4);
TASK_PP(16'h134E2,4);
TASK_PP(16'h134E3,4);
TASK_PP(16'h134E4,4);
TASK_PP(16'h134E5,4);
TASK_PP(16'h134E6,4);
TASK_PP(16'h134E7,4);
TASK_PP(16'h134E8,4);
TASK_PP(16'h134E9,4);
TASK_PP(16'h134EA,4);
TASK_PP(16'h134EB,4);
TASK_PP(16'h134EC,4);
TASK_PP(16'h134ED,4);
TASK_PP(16'h134EE,4);
TASK_PP(16'h134EF,4);
TASK_PP(16'h134F0,4);
TASK_PP(16'h134F1,4);
TASK_PP(16'h134F2,4);
TASK_PP(16'h134F3,4);
TASK_PP(16'h134F4,4);
TASK_PP(16'h134F5,4);
TASK_PP(16'h134F6,4);
TASK_PP(16'h134F7,4);
TASK_PP(16'h134F8,4);
TASK_PP(16'h134F9,4);
TASK_PP(16'h134FA,4);
TASK_PP(16'h134FB,4);
TASK_PP(16'h134FC,4);
TASK_PP(16'h134FD,4);
TASK_PP(16'h134FE,4);
TASK_PP(16'h134FF,4);
TASK_PP(16'h13500,4);
TASK_PP(16'h13501,4);
TASK_PP(16'h13502,4);
TASK_PP(16'h13503,4);
TASK_PP(16'h13504,4);
TASK_PP(16'h13505,4);
TASK_PP(16'h13506,4);
TASK_PP(16'h13507,4);
TASK_PP(16'h13508,4);
TASK_PP(16'h13509,4);
TASK_PP(16'h1350A,4);
TASK_PP(16'h1350B,4);
TASK_PP(16'h1350C,4);
TASK_PP(16'h1350D,4);
TASK_PP(16'h1350E,4);
TASK_PP(16'h1350F,4);
TASK_PP(16'h13510,4);
TASK_PP(16'h13511,4);
TASK_PP(16'h13512,4);
TASK_PP(16'h13513,4);
TASK_PP(16'h13514,4);
TASK_PP(16'h13515,4);
TASK_PP(16'h13516,4);
TASK_PP(16'h13517,4);
TASK_PP(16'h13518,4);
TASK_PP(16'h13519,4);
TASK_PP(16'h1351A,4);
TASK_PP(16'h1351B,4);
TASK_PP(16'h1351C,4);
TASK_PP(16'h1351D,4);
TASK_PP(16'h1351E,4);
TASK_PP(16'h1351F,4);
TASK_PP(16'h13520,4);
TASK_PP(16'h13521,4);
TASK_PP(16'h13522,4);
TASK_PP(16'h13523,4);
TASK_PP(16'h13524,4);
TASK_PP(16'h13525,4);
TASK_PP(16'h13526,4);
TASK_PP(16'h13527,4);
TASK_PP(16'h13528,4);
TASK_PP(16'h13529,4);
TASK_PP(16'h1352A,4);
TASK_PP(16'h1352B,4);
TASK_PP(16'h1352C,4);
TASK_PP(16'h1352D,4);
TASK_PP(16'h1352E,4);
TASK_PP(16'h1352F,4);
TASK_PP(16'h13530,4);
TASK_PP(16'h13531,4);
TASK_PP(16'h13532,4);
TASK_PP(16'h13533,4);
TASK_PP(16'h13534,4);
TASK_PP(16'h13535,4);
TASK_PP(16'h13536,4);
TASK_PP(16'h13537,4);
TASK_PP(16'h13538,4);
TASK_PP(16'h13539,4);
TASK_PP(16'h1353A,4);
TASK_PP(16'h1353B,4);
TASK_PP(16'h1353C,4);
TASK_PP(16'h1353D,4);
TASK_PP(16'h1353E,4);
TASK_PP(16'h1353F,4);
TASK_PP(16'h13540,4);
TASK_PP(16'h13541,4);
TASK_PP(16'h13542,4);
TASK_PP(16'h13543,4);
TASK_PP(16'h13544,4);
TASK_PP(16'h13545,4);
TASK_PP(16'h13546,4);
TASK_PP(16'h13547,4);
TASK_PP(16'h13548,4);
TASK_PP(16'h13549,4);
TASK_PP(16'h1354A,4);
TASK_PP(16'h1354B,4);
TASK_PP(16'h1354C,4);
TASK_PP(16'h1354D,4);
TASK_PP(16'h1354E,4);
TASK_PP(16'h1354F,4);
TASK_PP(16'h13550,4);
TASK_PP(16'h13551,4);
TASK_PP(16'h13552,4);
TASK_PP(16'h13553,4);
TASK_PP(16'h13554,4);
TASK_PP(16'h13555,4);
TASK_PP(16'h13556,4);
TASK_PP(16'h13557,4);
TASK_PP(16'h13558,4);
TASK_PP(16'h13559,4);
TASK_PP(16'h1355A,4);
TASK_PP(16'h1355B,4);
TASK_PP(16'h1355C,4);
TASK_PP(16'h1355D,4);
TASK_PP(16'h1355E,4);
TASK_PP(16'h1355F,4);
TASK_PP(16'h13560,4);
TASK_PP(16'h13561,4);
TASK_PP(16'h13562,4);
TASK_PP(16'h13563,4);
TASK_PP(16'h13564,4);
TASK_PP(16'h13565,4);
TASK_PP(16'h13566,4);
TASK_PP(16'h13567,4);
TASK_PP(16'h13568,4);
TASK_PP(16'h13569,4);
TASK_PP(16'h1356A,4);
TASK_PP(16'h1356B,4);
TASK_PP(16'h1356C,4);
TASK_PP(16'h1356D,4);
TASK_PP(16'h1356E,4);
TASK_PP(16'h1356F,4);
TASK_PP(16'h13570,4);
TASK_PP(16'h13571,4);
TASK_PP(16'h13572,4);
TASK_PP(16'h13573,4);
TASK_PP(16'h13574,4);
TASK_PP(16'h13575,4);
TASK_PP(16'h13576,4);
TASK_PP(16'h13577,4);
TASK_PP(16'h13578,4);
TASK_PP(16'h13579,4);
TASK_PP(16'h1357A,4);
TASK_PP(16'h1357B,4);
TASK_PP(16'h1357C,4);
TASK_PP(16'h1357D,4);
TASK_PP(16'h1357E,4);
TASK_PP(16'h1357F,4);
TASK_PP(16'h13580,4);
TASK_PP(16'h13581,4);
TASK_PP(16'h13582,4);
TASK_PP(16'h13583,4);
TASK_PP(16'h13584,4);
TASK_PP(16'h13585,4);
TASK_PP(16'h13586,4);
TASK_PP(16'h13587,4);
TASK_PP(16'h13588,4);
TASK_PP(16'h13589,4);
TASK_PP(16'h1358A,4);
TASK_PP(16'h1358B,4);
TASK_PP(16'h1358C,4);
TASK_PP(16'h1358D,4);
TASK_PP(16'h1358E,4);
TASK_PP(16'h1358F,4);
TASK_PP(16'h13590,4);
TASK_PP(16'h13591,4);
TASK_PP(16'h13592,4);
TASK_PP(16'h13593,4);
TASK_PP(16'h13594,4);
TASK_PP(16'h13595,4);
TASK_PP(16'h13596,4);
TASK_PP(16'h13597,4);
TASK_PP(16'h13598,4);
TASK_PP(16'h13599,4);
TASK_PP(16'h1359A,4);
TASK_PP(16'h1359B,4);
TASK_PP(16'h1359C,4);
TASK_PP(16'h1359D,4);
TASK_PP(16'h1359E,4);
TASK_PP(16'h1359F,4);
TASK_PP(16'h135A0,4);
TASK_PP(16'h135A1,4);
TASK_PP(16'h135A2,4);
TASK_PP(16'h135A3,4);
TASK_PP(16'h135A4,4);
TASK_PP(16'h135A5,4);
TASK_PP(16'h135A6,4);
TASK_PP(16'h135A7,4);
TASK_PP(16'h135A8,4);
TASK_PP(16'h135A9,4);
TASK_PP(16'h135AA,4);
TASK_PP(16'h135AB,4);
TASK_PP(16'h135AC,4);
TASK_PP(16'h135AD,4);
TASK_PP(16'h135AE,4);
TASK_PP(16'h135AF,4);
TASK_PP(16'h135B0,4);
TASK_PP(16'h135B1,4);
TASK_PP(16'h135B2,4);
TASK_PP(16'h135B3,4);
TASK_PP(16'h135B4,4);
TASK_PP(16'h135B5,4);
TASK_PP(16'h135B6,4);
TASK_PP(16'h135B7,4);
TASK_PP(16'h135B8,4);
TASK_PP(16'h135B9,4);
TASK_PP(16'h135BA,4);
TASK_PP(16'h135BB,4);
TASK_PP(16'h135BC,4);
TASK_PP(16'h135BD,4);
TASK_PP(16'h135BE,4);
TASK_PP(16'h135BF,4);
TASK_PP(16'h135C0,4);
TASK_PP(16'h135C1,4);
TASK_PP(16'h135C2,4);
TASK_PP(16'h135C3,4);
TASK_PP(16'h135C4,4);
TASK_PP(16'h135C5,4);
TASK_PP(16'h135C6,4);
TASK_PP(16'h135C7,4);
TASK_PP(16'h135C8,4);
TASK_PP(16'h135C9,4);
TASK_PP(16'h135CA,4);
TASK_PP(16'h135CB,4);
TASK_PP(16'h135CC,4);
TASK_PP(16'h135CD,4);
TASK_PP(16'h135CE,4);
TASK_PP(16'h135CF,4);
TASK_PP(16'h135D0,4);
TASK_PP(16'h135D1,4);
TASK_PP(16'h135D2,4);
TASK_PP(16'h135D3,4);
TASK_PP(16'h135D4,4);
TASK_PP(16'h135D5,4);
TASK_PP(16'h135D6,4);
TASK_PP(16'h135D7,4);
TASK_PP(16'h135D8,4);
TASK_PP(16'h135D9,4);
TASK_PP(16'h135DA,4);
TASK_PP(16'h135DB,4);
TASK_PP(16'h135DC,4);
TASK_PP(16'h135DD,4);
TASK_PP(16'h135DE,4);
TASK_PP(16'h135DF,4);
TASK_PP(16'h135E0,4);
TASK_PP(16'h135E1,4);
TASK_PP(16'h135E2,4);
TASK_PP(16'h135E3,4);
TASK_PP(16'h135E4,4);
TASK_PP(16'h135E5,4);
TASK_PP(16'h135E6,4);
TASK_PP(16'h135E7,4);
TASK_PP(16'h135E8,4);
TASK_PP(16'h135E9,4);
TASK_PP(16'h135EA,4);
TASK_PP(16'h135EB,4);
TASK_PP(16'h135EC,4);
TASK_PP(16'h135ED,4);
TASK_PP(16'h135EE,4);
TASK_PP(16'h135EF,4);
TASK_PP(16'h135F0,4);
TASK_PP(16'h135F1,4);
TASK_PP(16'h135F2,4);
TASK_PP(16'h135F3,4);
TASK_PP(16'h135F4,4);
TASK_PP(16'h135F5,4);
TASK_PP(16'h135F6,4);
TASK_PP(16'h135F7,4);
TASK_PP(16'h135F8,4);
TASK_PP(16'h135F9,4);
TASK_PP(16'h135FA,4);
TASK_PP(16'h135FB,4);
TASK_PP(16'h135FC,4);
TASK_PP(16'h135FD,4);
TASK_PP(16'h135FE,4);
TASK_PP(16'h135FF,4);
TASK_PP(16'h13600,4);
TASK_PP(16'h13601,4);
TASK_PP(16'h13602,4);
TASK_PP(16'h13603,4);
TASK_PP(16'h13604,4);
TASK_PP(16'h13605,4);
TASK_PP(16'h13606,4);
TASK_PP(16'h13607,4);
TASK_PP(16'h13608,4);
TASK_PP(16'h13609,4);
TASK_PP(16'h1360A,4);
TASK_PP(16'h1360B,4);
TASK_PP(16'h1360C,4);
TASK_PP(16'h1360D,4);
TASK_PP(16'h1360E,4);
TASK_PP(16'h1360F,4);
TASK_PP(16'h13610,4);
TASK_PP(16'h13611,4);
TASK_PP(16'h13612,4);
TASK_PP(16'h13613,4);
TASK_PP(16'h13614,4);
TASK_PP(16'h13615,4);
TASK_PP(16'h13616,4);
TASK_PP(16'h13617,4);
TASK_PP(16'h13618,4);
TASK_PP(16'h13619,4);
TASK_PP(16'h1361A,4);
TASK_PP(16'h1361B,4);
TASK_PP(16'h1361C,4);
TASK_PP(16'h1361D,4);
TASK_PP(16'h1361E,4);
TASK_PP(16'h1361F,4);
TASK_PP(16'h13620,4);
TASK_PP(16'h13621,4);
TASK_PP(16'h13622,4);
TASK_PP(16'h13623,4);
TASK_PP(16'h13624,4);
TASK_PP(16'h13625,4);
TASK_PP(16'h13626,4);
TASK_PP(16'h13627,4);
TASK_PP(16'h13628,4);
TASK_PP(16'h13629,4);
TASK_PP(16'h1362A,4);
TASK_PP(16'h1362B,4);
TASK_PP(16'h1362C,4);
TASK_PP(16'h1362D,4);
TASK_PP(16'h1362E,4);
TASK_PP(16'h1362F,4);
TASK_PP(16'h13630,4);
TASK_PP(16'h13631,4);
TASK_PP(16'h13632,4);
TASK_PP(16'h13633,4);
TASK_PP(16'h13634,4);
TASK_PP(16'h13635,4);
TASK_PP(16'h13636,4);
TASK_PP(16'h13637,4);
TASK_PP(16'h13638,4);
TASK_PP(16'h13639,4);
TASK_PP(16'h1363A,4);
TASK_PP(16'h1363B,4);
TASK_PP(16'h1363C,4);
TASK_PP(16'h1363D,4);
TASK_PP(16'h1363E,4);
TASK_PP(16'h1363F,4);
TASK_PP(16'h13640,4);
TASK_PP(16'h13641,4);
TASK_PP(16'h13642,4);
TASK_PP(16'h13643,4);
TASK_PP(16'h13644,4);
TASK_PP(16'h13645,4);
TASK_PP(16'h13646,4);
TASK_PP(16'h13647,4);
TASK_PP(16'h13648,4);
TASK_PP(16'h13649,4);
TASK_PP(16'h1364A,4);
TASK_PP(16'h1364B,4);
TASK_PP(16'h1364C,4);
TASK_PP(16'h1364D,4);
TASK_PP(16'h1364E,4);
TASK_PP(16'h1364F,4);
TASK_PP(16'h13650,4);
TASK_PP(16'h13651,4);
TASK_PP(16'h13652,4);
TASK_PP(16'h13653,4);
TASK_PP(16'h13654,4);
TASK_PP(16'h13655,4);
TASK_PP(16'h13656,4);
TASK_PP(16'h13657,4);
TASK_PP(16'h13658,4);
TASK_PP(16'h13659,4);
TASK_PP(16'h1365A,4);
TASK_PP(16'h1365B,4);
TASK_PP(16'h1365C,4);
TASK_PP(16'h1365D,4);
TASK_PP(16'h1365E,4);
TASK_PP(16'h1365F,4);
TASK_PP(16'h13660,4);
TASK_PP(16'h13661,4);
TASK_PP(16'h13662,4);
TASK_PP(16'h13663,4);
TASK_PP(16'h13664,4);
TASK_PP(16'h13665,4);
TASK_PP(16'h13666,4);
TASK_PP(16'h13667,4);
TASK_PP(16'h13668,4);
TASK_PP(16'h13669,4);
TASK_PP(16'h1366A,4);
TASK_PP(16'h1366B,4);
TASK_PP(16'h1366C,4);
TASK_PP(16'h1366D,4);
TASK_PP(16'h1366E,4);
TASK_PP(16'h1366F,4);
TASK_PP(16'h13670,4);
TASK_PP(16'h13671,4);
TASK_PP(16'h13672,4);
TASK_PP(16'h13673,4);
TASK_PP(16'h13674,4);
TASK_PP(16'h13675,4);
TASK_PP(16'h13676,4);
TASK_PP(16'h13677,4);
TASK_PP(16'h13678,4);
TASK_PP(16'h13679,4);
TASK_PP(16'h1367A,4);
TASK_PP(16'h1367B,4);
TASK_PP(16'h1367C,4);
TASK_PP(16'h1367D,4);
TASK_PP(16'h1367E,4);
TASK_PP(16'h1367F,4);
TASK_PP(16'h13680,4);
TASK_PP(16'h13681,4);
TASK_PP(16'h13682,4);
TASK_PP(16'h13683,4);
TASK_PP(16'h13684,4);
TASK_PP(16'h13685,4);
TASK_PP(16'h13686,4);
TASK_PP(16'h13687,4);
TASK_PP(16'h13688,4);
TASK_PP(16'h13689,4);
TASK_PP(16'h1368A,4);
TASK_PP(16'h1368B,4);
TASK_PP(16'h1368C,4);
TASK_PP(16'h1368D,4);
TASK_PP(16'h1368E,4);
TASK_PP(16'h1368F,4);
TASK_PP(16'h13690,4);
TASK_PP(16'h13691,4);
TASK_PP(16'h13692,4);
TASK_PP(16'h13693,4);
TASK_PP(16'h13694,4);
TASK_PP(16'h13695,4);
TASK_PP(16'h13696,4);
TASK_PP(16'h13697,4);
TASK_PP(16'h13698,4);
TASK_PP(16'h13699,4);
TASK_PP(16'h1369A,4);
TASK_PP(16'h1369B,4);
TASK_PP(16'h1369C,4);
TASK_PP(16'h1369D,4);
TASK_PP(16'h1369E,4);
TASK_PP(16'h1369F,4);
TASK_PP(16'h136A0,4);
TASK_PP(16'h136A1,4);
TASK_PP(16'h136A2,4);
TASK_PP(16'h136A3,4);
TASK_PP(16'h136A4,4);
TASK_PP(16'h136A5,4);
TASK_PP(16'h136A6,4);
TASK_PP(16'h136A7,4);
TASK_PP(16'h136A8,4);
TASK_PP(16'h136A9,4);
TASK_PP(16'h136AA,4);
TASK_PP(16'h136AB,4);
TASK_PP(16'h136AC,4);
TASK_PP(16'h136AD,4);
TASK_PP(16'h136AE,4);
TASK_PP(16'h136AF,4);
TASK_PP(16'h136B0,4);
TASK_PP(16'h136B1,4);
TASK_PP(16'h136B2,4);
TASK_PP(16'h136B3,4);
TASK_PP(16'h136B4,4);
TASK_PP(16'h136B5,4);
TASK_PP(16'h136B6,4);
TASK_PP(16'h136B7,4);
TASK_PP(16'h136B8,4);
TASK_PP(16'h136B9,4);
TASK_PP(16'h136BA,4);
TASK_PP(16'h136BB,4);
TASK_PP(16'h136BC,4);
TASK_PP(16'h136BD,4);
TASK_PP(16'h136BE,4);
TASK_PP(16'h136BF,4);
TASK_PP(16'h136C0,4);
TASK_PP(16'h136C1,4);
TASK_PP(16'h136C2,4);
TASK_PP(16'h136C3,4);
TASK_PP(16'h136C4,4);
TASK_PP(16'h136C5,4);
TASK_PP(16'h136C6,4);
TASK_PP(16'h136C7,4);
TASK_PP(16'h136C8,4);
TASK_PP(16'h136C9,4);
TASK_PP(16'h136CA,4);
TASK_PP(16'h136CB,4);
TASK_PP(16'h136CC,4);
TASK_PP(16'h136CD,4);
TASK_PP(16'h136CE,4);
TASK_PP(16'h136CF,4);
TASK_PP(16'h136D0,4);
TASK_PP(16'h136D1,4);
TASK_PP(16'h136D2,4);
TASK_PP(16'h136D3,4);
TASK_PP(16'h136D4,4);
TASK_PP(16'h136D5,4);
TASK_PP(16'h136D6,4);
TASK_PP(16'h136D7,4);
TASK_PP(16'h136D8,4);
TASK_PP(16'h136D9,4);
TASK_PP(16'h136DA,4);
TASK_PP(16'h136DB,4);
TASK_PP(16'h136DC,4);
TASK_PP(16'h136DD,4);
TASK_PP(16'h136DE,4);
TASK_PP(16'h136DF,4);
TASK_PP(16'h136E0,4);
TASK_PP(16'h136E1,4);
TASK_PP(16'h136E2,4);
TASK_PP(16'h136E3,4);
TASK_PP(16'h136E4,4);
TASK_PP(16'h136E5,4);
TASK_PP(16'h136E6,4);
TASK_PP(16'h136E7,4);
TASK_PP(16'h136E8,4);
TASK_PP(16'h136E9,4);
TASK_PP(16'h136EA,4);
TASK_PP(16'h136EB,4);
TASK_PP(16'h136EC,4);
TASK_PP(16'h136ED,4);
TASK_PP(16'h136EE,4);
TASK_PP(16'h136EF,4);
TASK_PP(16'h136F0,4);
TASK_PP(16'h136F1,4);
TASK_PP(16'h136F2,4);
TASK_PP(16'h136F3,4);
TASK_PP(16'h136F4,4);
TASK_PP(16'h136F5,4);
TASK_PP(16'h136F6,4);
TASK_PP(16'h136F7,4);
TASK_PP(16'h136F8,4);
TASK_PP(16'h136F9,4);
TASK_PP(16'h136FA,4);
TASK_PP(16'h136FB,4);
TASK_PP(16'h136FC,4);
TASK_PP(16'h136FD,4);
TASK_PP(16'h136FE,4);
TASK_PP(16'h136FF,4);
TASK_PP(16'h13700,4);
TASK_PP(16'h13701,4);
TASK_PP(16'h13702,4);
TASK_PP(16'h13703,4);
TASK_PP(16'h13704,4);
TASK_PP(16'h13705,4);
TASK_PP(16'h13706,4);
TASK_PP(16'h13707,4);
TASK_PP(16'h13708,4);
TASK_PP(16'h13709,4);
TASK_PP(16'h1370A,4);
TASK_PP(16'h1370B,4);
TASK_PP(16'h1370C,4);
TASK_PP(16'h1370D,4);
TASK_PP(16'h1370E,4);
TASK_PP(16'h1370F,4);
TASK_PP(16'h13710,4);
TASK_PP(16'h13711,4);
TASK_PP(16'h13712,4);
TASK_PP(16'h13713,4);
TASK_PP(16'h13714,4);
TASK_PP(16'h13715,4);
TASK_PP(16'h13716,4);
TASK_PP(16'h13717,4);
TASK_PP(16'h13718,4);
TASK_PP(16'h13719,4);
TASK_PP(16'h1371A,4);
TASK_PP(16'h1371B,4);
TASK_PP(16'h1371C,4);
TASK_PP(16'h1371D,4);
TASK_PP(16'h1371E,4);
TASK_PP(16'h1371F,4);
TASK_PP(16'h13720,4);
TASK_PP(16'h13721,4);
TASK_PP(16'h13722,4);
TASK_PP(16'h13723,4);
TASK_PP(16'h13724,4);
TASK_PP(16'h13725,4);
TASK_PP(16'h13726,4);
TASK_PP(16'h13727,4);
TASK_PP(16'h13728,4);
TASK_PP(16'h13729,4);
TASK_PP(16'h1372A,4);
TASK_PP(16'h1372B,4);
TASK_PP(16'h1372C,4);
TASK_PP(16'h1372D,4);
TASK_PP(16'h1372E,4);
TASK_PP(16'h1372F,4);
TASK_PP(16'h13730,4);
TASK_PP(16'h13731,4);
TASK_PP(16'h13732,4);
TASK_PP(16'h13733,4);
TASK_PP(16'h13734,4);
TASK_PP(16'h13735,4);
TASK_PP(16'h13736,4);
TASK_PP(16'h13737,4);
TASK_PP(16'h13738,4);
TASK_PP(16'h13739,4);
TASK_PP(16'h1373A,4);
TASK_PP(16'h1373B,4);
TASK_PP(16'h1373C,4);
TASK_PP(16'h1373D,4);
TASK_PP(16'h1373E,4);
TASK_PP(16'h1373F,4);
TASK_PP(16'h13740,4);
TASK_PP(16'h13741,4);
TASK_PP(16'h13742,4);
TASK_PP(16'h13743,4);
TASK_PP(16'h13744,4);
TASK_PP(16'h13745,4);
TASK_PP(16'h13746,4);
TASK_PP(16'h13747,4);
TASK_PP(16'h13748,4);
TASK_PP(16'h13749,4);
TASK_PP(16'h1374A,4);
TASK_PP(16'h1374B,4);
TASK_PP(16'h1374C,4);
TASK_PP(16'h1374D,4);
TASK_PP(16'h1374E,4);
TASK_PP(16'h1374F,4);
TASK_PP(16'h13750,4);
TASK_PP(16'h13751,4);
TASK_PP(16'h13752,4);
TASK_PP(16'h13753,4);
TASK_PP(16'h13754,4);
TASK_PP(16'h13755,4);
TASK_PP(16'h13756,4);
TASK_PP(16'h13757,4);
TASK_PP(16'h13758,4);
TASK_PP(16'h13759,4);
TASK_PP(16'h1375A,4);
TASK_PP(16'h1375B,4);
TASK_PP(16'h1375C,4);
TASK_PP(16'h1375D,4);
TASK_PP(16'h1375E,4);
TASK_PP(16'h1375F,4);
TASK_PP(16'h13760,4);
TASK_PP(16'h13761,4);
TASK_PP(16'h13762,4);
TASK_PP(16'h13763,4);
TASK_PP(16'h13764,4);
TASK_PP(16'h13765,4);
TASK_PP(16'h13766,4);
TASK_PP(16'h13767,4);
TASK_PP(16'h13768,4);
TASK_PP(16'h13769,4);
TASK_PP(16'h1376A,4);
TASK_PP(16'h1376B,4);
TASK_PP(16'h1376C,4);
TASK_PP(16'h1376D,4);
TASK_PP(16'h1376E,4);
TASK_PP(16'h1376F,4);
TASK_PP(16'h13770,4);
TASK_PP(16'h13771,4);
TASK_PP(16'h13772,4);
TASK_PP(16'h13773,4);
TASK_PP(16'h13774,4);
TASK_PP(16'h13775,4);
TASK_PP(16'h13776,4);
TASK_PP(16'h13777,4);
TASK_PP(16'h13778,4);
TASK_PP(16'h13779,4);
TASK_PP(16'h1377A,4);
TASK_PP(16'h1377B,4);
TASK_PP(16'h1377C,4);
TASK_PP(16'h1377D,4);
TASK_PP(16'h1377E,4);
TASK_PP(16'h1377F,4);
TASK_PP(16'h13780,4);
TASK_PP(16'h13781,4);
TASK_PP(16'h13782,4);
TASK_PP(16'h13783,4);
TASK_PP(16'h13784,4);
TASK_PP(16'h13785,4);
TASK_PP(16'h13786,4);
TASK_PP(16'h13787,4);
TASK_PP(16'h13788,4);
TASK_PP(16'h13789,4);
TASK_PP(16'h1378A,4);
TASK_PP(16'h1378B,4);
TASK_PP(16'h1378C,4);
TASK_PP(16'h1378D,4);
TASK_PP(16'h1378E,4);
TASK_PP(16'h1378F,4);
TASK_PP(16'h13790,4);
TASK_PP(16'h13791,4);
TASK_PP(16'h13792,4);
TASK_PP(16'h13793,4);
TASK_PP(16'h13794,4);
TASK_PP(16'h13795,4);
TASK_PP(16'h13796,4);
TASK_PP(16'h13797,4);
TASK_PP(16'h13798,4);
TASK_PP(16'h13799,4);
TASK_PP(16'h1379A,4);
TASK_PP(16'h1379B,4);
TASK_PP(16'h1379C,4);
TASK_PP(16'h1379D,4);
TASK_PP(16'h1379E,4);
TASK_PP(16'h1379F,4);
TASK_PP(16'h137A0,4);
TASK_PP(16'h137A1,4);
TASK_PP(16'h137A2,4);
TASK_PP(16'h137A3,4);
TASK_PP(16'h137A4,4);
TASK_PP(16'h137A5,4);
TASK_PP(16'h137A6,4);
TASK_PP(16'h137A7,4);
TASK_PP(16'h137A8,4);
TASK_PP(16'h137A9,4);
TASK_PP(16'h137AA,4);
TASK_PP(16'h137AB,4);
TASK_PP(16'h137AC,4);
TASK_PP(16'h137AD,4);
TASK_PP(16'h137AE,4);
TASK_PP(16'h137AF,4);
TASK_PP(16'h137B0,4);
TASK_PP(16'h137B1,4);
TASK_PP(16'h137B2,4);
TASK_PP(16'h137B3,4);
TASK_PP(16'h137B4,4);
TASK_PP(16'h137B5,4);
TASK_PP(16'h137B6,4);
TASK_PP(16'h137B7,4);
TASK_PP(16'h137B8,4);
TASK_PP(16'h137B9,4);
TASK_PP(16'h137BA,4);
TASK_PP(16'h137BB,4);
TASK_PP(16'h137BC,4);
TASK_PP(16'h137BD,4);
TASK_PP(16'h137BE,4);
TASK_PP(16'h137BF,4);
TASK_PP(16'h137C0,4);
TASK_PP(16'h137C1,4);
TASK_PP(16'h137C2,4);
TASK_PP(16'h137C3,4);
TASK_PP(16'h137C4,4);
TASK_PP(16'h137C5,4);
TASK_PP(16'h137C6,4);
TASK_PP(16'h137C7,4);
TASK_PP(16'h137C8,4);
TASK_PP(16'h137C9,4);
TASK_PP(16'h137CA,4);
TASK_PP(16'h137CB,4);
TASK_PP(16'h137CC,4);
TASK_PP(16'h137CD,4);
TASK_PP(16'h137CE,4);
TASK_PP(16'h137CF,4);
TASK_PP(16'h137D0,4);
TASK_PP(16'h137D1,4);
TASK_PP(16'h137D2,4);
TASK_PP(16'h137D3,4);
TASK_PP(16'h137D4,4);
TASK_PP(16'h137D5,4);
TASK_PP(16'h137D6,4);
TASK_PP(16'h137D7,4);
TASK_PP(16'h137D8,4);
TASK_PP(16'h137D9,4);
TASK_PP(16'h137DA,4);
TASK_PP(16'h137DB,4);
TASK_PP(16'h137DC,4);
TASK_PP(16'h137DD,4);
TASK_PP(16'h137DE,4);
TASK_PP(16'h137DF,4);
TASK_PP(16'h137E0,4);
TASK_PP(16'h137E1,4);
TASK_PP(16'h137E2,4);
TASK_PP(16'h137E3,4);
TASK_PP(16'h137E4,4);
TASK_PP(16'h137E5,4);
TASK_PP(16'h137E6,4);
TASK_PP(16'h137E7,4);
TASK_PP(16'h137E8,4);
TASK_PP(16'h137E9,4);
TASK_PP(16'h137EA,4);
TASK_PP(16'h137EB,4);
TASK_PP(16'h137EC,4);
TASK_PP(16'h137ED,4);
TASK_PP(16'h137EE,4);
TASK_PP(16'h137EF,4);
TASK_PP(16'h137F0,4);
TASK_PP(16'h137F1,4);
TASK_PP(16'h137F2,4);
TASK_PP(16'h137F3,4);
TASK_PP(16'h137F4,4);
TASK_PP(16'h137F5,4);
TASK_PP(16'h137F6,4);
TASK_PP(16'h137F7,4);
TASK_PP(16'h137F8,4);
TASK_PP(16'h137F9,4);
TASK_PP(16'h137FA,4);
TASK_PP(16'h137FB,4);
TASK_PP(16'h137FC,4);
TASK_PP(16'h137FD,4);
TASK_PP(16'h137FE,4);
TASK_PP(16'h137FF,4);
TASK_PP(16'h13800,4);
TASK_PP(16'h13801,4);
TASK_PP(16'h13802,4);
TASK_PP(16'h13803,4);
TASK_PP(16'h13804,4);
TASK_PP(16'h13805,4);
TASK_PP(16'h13806,4);
TASK_PP(16'h13807,4);
TASK_PP(16'h13808,4);
TASK_PP(16'h13809,4);
TASK_PP(16'h1380A,4);
TASK_PP(16'h1380B,4);
TASK_PP(16'h1380C,4);
TASK_PP(16'h1380D,4);
TASK_PP(16'h1380E,4);
TASK_PP(16'h1380F,4);
TASK_PP(16'h13810,4);
TASK_PP(16'h13811,4);
TASK_PP(16'h13812,4);
TASK_PP(16'h13813,4);
TASK_PP(16'h13814,4);
TASK_PP(16'h13815,4);
TASK_PP(16'h13816,4);
TASK_PP(16'h13817,4);
TASK_PP(16'h13818,4);
TASK_PP(16'h13819,4);
TASK_PP(16'h1381A,4);
TASK_PP(16'h1381B,4);
TASK_PP(16'h1381C,4);
TASK_PP(16'h1381D,4);
TASK_PP(16'h1381E,4);
TASK_PP(16'h1381F,4);
TASK_PP(16'h13820,4);
TASK_PP(16'h13821,4);
TASK_PP(16'h13822,4);
TASK_PP(16'h13823,4);
TASK_PP(16'h13824,4);
TASK_PP(16'h13825,4);
TASK_PP(16'h13826,4);
TASK_PP(16'h13827,4);
TASK_PP(16'h13828,4);
TASK_PP(16'h13829,4);
TASK_PP(16'h1382A,4);
TASK_PP(16'h1382B,4);
TASK_PP(16'h1382C,4);
TASK_PP(16'h1382D,4);
TASK_PP(16'h1382E,4);
TASK_PP(16'h1382F,4);
TASK_PP(16'h13830,4);
TASK_PP(16'h13831,4);
TASK_PP(16'h13832,4);
TASK_PP(16'h13833,4);
TASK_PP(16'h13834,4);
TASK_PP(16'h13835,4);
TASK_PP(16'h13836,4);
TASK_PP(16'h13837,4);
TASK_PP(16'h13838,4);
TASK_PP(16'h13839,4);
TASK_PP(16'h1383A,4);
TASK_PP(16'h1383B,4);
TASK_PP(16'h1383C,4);
TASK_PP(16'h1383D,4);
TASK_PP(16'h1383E,4);
TASK_PP(16'h1383F,4);
TASK_PP(16'h13840,4);
TASK_PP(16'h13841,4);
TASK_PP(16'h13842,4);
TASK_PP(16'h13843,4);
TASK_PP(16'h13844,4);
TASK_PP(16'h13845,4);
TASK_PP(16'h13846,4);
TASK_PP(16'h13847,4);
TASK_PP(16'h13848,4);
TASK_PP(16'h13849,4);
TASK_PP(16'h1384A,4);
TASK_PP(16'h1384B,4);
TASK_PP(16'h1384C,4);
TASK_PP(16'h1384D,4);
TASK_PP(16'h1384E,4);
TASK_PP(16'h1384F,4);
TASK_PP(16'h13850,4);
TASK_PP(16'h13851,4);
TASK_PP(16'h13852,4);
TASK_PP(16'h13853,4);
TASK_PP(16'h13854,4);
TASK_PP(16'h13855,4);
TASK_PP(16'h13856,4);
TASK_PP(16'h13857,4);
TASK_PP(16'h13858,4);
TASK_PP(16'h13859,4);
TASK_PP(16'h1385A,4);
TASK_PP(16'h1385B,4);
TASK_PP(16'h1385C,4);
TASK_PP(16'h1385D,4);
TASK_PP(16'h1385E,4);
TASK_PP(16'h1385F,4);
TASK_PP(16'h13860,4);
TASK_PP(16'h13861,4);
TASK_PP(16'h13862,4);
TASK_PP(16'h13863,4);
TASK_PP(16'h13864,4);
TASK_PP(16'h13865,4);
TASK_PP(16'h13866,4);
TASK_PP(16'h13867,4);
TASK_PP(16'h13868,4);
TASK_PP(16'h13869,4);
TASK_PP(16'h1386A,4);
TASK_PP(16'h1386B,4);
TASK_PP(16'h1386C,4);
TASK_PP(16'h1386D,4);
TASK_PP(16'h1386E,4);
TASK_PP(16'h1386F,4);
TASK_PP(16'h13870,4);
TASK_PP(16'h13871,4);
TASK_PP(16'h13872,4);
TASK_PP(16'h13873,4);
TASK_PP(16'h13874,4);
TASK_PP(16'h13875,4);
TASK_PP(16'h13876,4);
TASK_PP(16'h13877,4);
TASK_PP(16'h13878,4);
TASK_PP(16'h13879,4);
TASK_PP(16'h1387A,4);
TASK_PP(16'h1387B,4);
TASK_PP(16'h1387C,4);
TASK_PP(16'h1387D,4);
TASK_PP(16'h1387E,4);
TASK_PP(16'h1387F,4);
TASK_PP(16'h13880,4);
TASK_PP(16'h13881,4);
TASK_PP(16'h13882,4);
TASK_PP(16'h13883,4);
TASK_PP(16'h13884,4);
TASK_PP(16'h13885,4);
TASK_PP(16'h13886,4);
TASK_PP(16'h13887,4);
TASK_PP(16'h13888,4);
TASK_PP(16'h13889,4);
TASK_PP(16'h1388A,4);
TASK_PP(16'h1388B,4);
TASK_PP(16'h1388C,4);
TASK_PP(16'h1388D,4);
TASK_PP(16'h1388E,4);
TASK_PP(16'h1388F,4);
TASK_PP(16'h13890,4);
TASK_PP(16'h13891,4);
TASK_PP(16'h13892,4);
TASK_PP(16'h13893,4);
TASK_PP(16'h13894,4);
TASK_PP(16'h13895,4);
TASK_PP(16'h13896,4);
TASK_PP(16'h13897,4);
TASK_PP(16'h13898,4);
TASK_PP(16'h13899,4);
TASK_PP(16'h1389A,4);
TASK_PP(16'h1389B,4);
TASK_PP(16'h1389C,4);
TASK_PP(16'h1389D,4);
TASK_PP(16'h1389E,4);
TASK_PP(16'h1389F,4);
TASK_PP(16'h138A0,4);
TASK_PP(16'h138A1,4);
TASK_PP(16'h138A2,4);
TASK_PP(16'h138A3,4);
TASK_PP(16'h138A4,4);
TASK_PP(16'h138A5,4);
TASK_PP(16'h138A6,4);
TASK_PP(16'h138A7,4);
TASK_PP(16'h138A8,4);
TASK_PP(16'h138A9,4);
TASK_PP(16'h138AA,4);
TASK_PP(16'h138AB,4);
TASK_PP(16'h138AC,4);
TASK_PP(16'h138AD,4);
TASK_PP(16'h138AE,4);
TASK_PP(16'h138AF,4);
TASK_PP(16'h138B0,4);
TASK_PP(16'h138B1,4);
TASK_PP(16'h138B2,4);
TASK_PP(16'h138B3,4);
TASK_PP(16'h138B4,4);
TASK_PP(16'h138B5,4);
TASK_PP(16'h138B6,4);
TASK_PP(16'h138B7,4);
TASK_PP(16'h138B8,4);
TASK_PP(16'h138B9,4);
TASK_PP(16'h138BA,4);
TASK_PP(16'h138BB,4);
TASK_PP(16'h138BC,4);
TASK_PP(16'h138BD,4);
TASK_PP(16'h138BE,4);
TASK_PP(16'h138BF,4);
TASK_PP(16'h138C0,4);
TASK_PP(16'h138C1,4);
TASK_PP(16'h138C2,4);
TASK_PP(16'h138C3,4);
TASK_PP(16'h138C4,4);
TASK_PP(16'h138C5,4);
TASK_PP(16'h138C6,4);
TASK_PP(16'h138C7,4);
TASK_PP(16'h138C8,4);
TASK_PP(16'h138C9,4);
TASK_PP(16'h138CA,4);
TASK_PP(16'h138CB,4);
TASK_PP(16'h138CC,4);
TASK_PP(16'h138CD,4);
TASK_PP(16'h138CE,4);
TASK_PP(16'h138CF,4);
TASK_PP(16'h138D0,4);
TASK_PP(16'h138D1,4);
TASK_PP(16'h138D2,4);
TASK_PP(16'h138D3,4);
TASK_PP(16'h138D4,4);
TASK_PP(16'h138D5,4);
TASK_PP(16'h138D6,4);
TASK_PP(16'h138D7,4);
TASK_PP(16'h138D8,4);
TASK_PP(16'h138D9,4);
TASK_PP(16'h138DA,4);
TASK_PP(16'h138DB,4);
TASK_PP(16'h138DC,4);
TASK_PP(16'h138DD,4);
TASK_PP(16'h138DE,4);
TASK_PP(16'h138DF,4);
TASK_PP(16'h138E0,4);
TASK_PP(16'h138E1,4);
TASK_PP(16'h138E2,4);
TASK_PP(16'h138E3,4);
TASK_PP(16'h138E4,4);
TASK_PP(16'h138E5,4);
TASK_PP(16'h138E6,4);
TASK_PP(16'h138E7,4);
TASK_PP(16'h138E8,4);
TASK_PP(16'h138E9,4);
TASK_PP(16'h138EA,4);
TASK_PP(16'h138EB,4);
TASK_PP(16'h138EC,4);
TASK_PP(16'h138ED,4);
TASK_PP(16'h138EE,4);
TASK_PP(16'h138EF,4);
TASK_PP(16'h138F0,4);
TASK_PP(16'h138F1,4);
TASK_PP(16'h138F2,4);
TASK_PP(16'h138F3,4);
TASK_PP(16'h138F4,4);
TASK_PP(16'h138F5,4);
TASK_PP(16'h138F6,4);
TASK_PP(16'h138F7,4);
TASK_PP(16'h138F8,4);
TASK_PP(16'h138F9,4);
TASK_PP(16'h138FA,4);
TASK_PP(16'h138FB,4);
TASK_PP(16'h138FC,4);
TASK_PP(16'h138FD,4);
TASK_PP(16'h138FE,4);
TASK_PP(16'h138FF,4);
TASK_PP(16'h13900,4);
TASK_PP(16'h13901,4);
TASK_PP(16'h13902,4);
TASK_PP(16'h13903,4);
TASK_PP(16'h13904,4);
TASK_PP(16'h13905,4);
TASK_PP(16'h13906,4);
TASK_PP(16'h13907,4);
TASK_PP(16'h13908,4);
TASK_PP(16'h13909,4);
TASK_PP(16'h1390A,4);
TASK_PP(16'h1390B,4);
TASK_PP(16'h1390C,4);
TASK_PP(16'h1390D,4);
TASK_PP(16'h1390E,4);
TASK_PP(16'h1390F,4);
TASK_PP(16'h13910,4);
TASK_PP(16'h13911,4);
TASK_PP(16'h13912,4);
TASK_PP(16'h13913,4);
TASK_PP(16'h13914,4);
TASK_PP(16'h13915,4);
TASK_PP(16'h13916,4);
TASK_PP(16'h13917,4);
TASK_PP(16'h13918,4);
TASK_PP(16'h13919,4);
TASK_PP(16'h1391A,4);
TASK_PP(16'h1391B,4);
TASK_PP(16'h1391C,4);
TASK_PP(16'h1391D,4);
TASK_PP(16'h1391E,4);
TASK_PP(16'h1391F,4);
TASK_PP(16'h13920,4);
TASK_PP(16'h13921,4);
TASK_PP(16'h13922,4);
TASK_PP(16'h13923,4);
TASK_PP(16'h13924,4);
TASK_PP(16'h13925,4);
TASK_PP(16'h13926,4);
TASK_PP(16'h13927,4);
TASK_PP(16'h13928,4);
TASK_PP(16'h13929,4);
TASK_PP(16'h1392A,4);
TASK_PP(16'h1392B,4);
TASK_PP(16'h1392C,4);
TASK_PP(16'h1392D,4);
TASK_PP(16'h1392E,4);
TASK_PP(16'h1392F,4);
TASK_PP(16'h13930,4);
TASK_PP(16'h13931,4);
TASK_PP(16'h13932,4);
TASK_PP(16'h13933,4);
TASK_PP(16'h13934,4);
TASK_PP(16'h13935,4);
TASK_PP(16'h13936,4);
TASK_PP(16'h13937,4);
TASK_PP(16'h13938,4);
TASK_PP(16'h13939,4);
TASK_PP(16'h1393A,4);
TASK_PP(16'h1393B,4);
TASK_PP(16'h1393C,4);
TASK_PP(16'h1393D,4);
TASK_PP(16'h1393E,4);
TASK_PP(16'h1393F,4);
TASK_PP(16'h13940,4);
TASK_PP(16'h13941,4);
TASK_PP(16'h13942,4);
TASK_PP(16'h13943,4);
TASK_PP(16'h13944,4);
TASK_PP(16'h13945,4);
TASK_PP(16'h13946,4);
TASK_PP(16'h13947,4);
TASK_PP(16'h13948,4);
TASK_PP(16'h13949,4);
TASK_PP(16'h1394A,4);
TASK_PP(16'h1394B,4);
TASK_PP(16'h1394C,4);
TASK_PP(16'h1394D,4);
TASK_PP(16'h1394E,4);
TASK_PP(16'h1394F,4);
TASK_PP(16'h13950,4);
TASK_PP(16'h13951,4);
TASK_PP(16'h13952,4);
TASK_PP(16'h13953,4);
TASK_PP(16'h13954,4);
TASK_PP(16'h13955,4);
TASK_PP(16'h13956,4);
TASK_PP(16'h13957,4);
TASK_PP(16'h13958,4);
TASK_PP(16'h13959,4);
TASK_PP(16'h1395A,4);
TASK_PP(16'h1395B,4);
TASK_PP(16'h1395C,4);
TASK_PP(16'h1395D,4);
TASK_PP(16'h1395E,4);
TASK_PP(16'h1395F,4);
TASK_PP(16'h13960,4);
TASK_PP(16'h13961,4);
TASK_PP(16'h13962,4);
TASK_PP(16'h13963,4);
TASK_PP(16'h13964,4);
TASK_PP(16'h13965,4);
TASK_PP(16'h13966,4);
TASK_PP(16'h13967,4);
TASK_PP(16'h13968,4);
TASK_PP(16'h13969,4);
TASK_PP(16'h1396A,4);
TASK_PP(16'h1396B,4);
TASK_PP(16'h1396C,4);
TASK_PP(16'h1396D,4);
TASK_PP(16'h1396E,4);
TASK_PP(16'h1396F,4);
TASK_PP(16'h13970,4);
TASK_PP(16'h13971,4);
TASK_PP(16'h13972,4);
TASK_PP(16'h13973,4);
TASK_PP(16'h13974,4);
TASK_PP(16'h13975,4);
TASK_PP(16'h13976,4);
TASK_PP(16'h13977,4);
TASK_PP(16'h13978,4);
TASK_PP(16'h13979,4);
TASK_PP(16'h1397A,4);
TASK_PP(16'h1397B,4);
TASK_PP(16'h1397C,4);
TASK_PP(16'h1397D,4);
TASK_PP(16'h1397E,4);
TASK_PP(16'h1397F,4);
TASK_PP(16'h13980,4);
TASK_PP(16'h13981,4);
TASK_PP(16'h13982,4);
TASK_PP(16'h13983,4);
TASK_PP(16'h13984,4);
TASK_PP(16'h13985,4);
TASK_PP(16'h13986,4);
TASK_PP(16'h13987,4);
TASK_PP(16'h13988,4);
TASK_PP(16'h13989,4);
TASK_PP(16'h1398A,4);
TASK_PP(16'h1398B,4);
TASK_PP(16'h1398C,4);
TASK_PP(16'h1398D,4);
TASK_PP(16'h1398E,4);
TASK_PP(16'h1398F,4);
TASK_PP(16'h13990,4);
TASK_PP(16'h13991,4);
TASK_PP(16'h13992,4);
TASK_PP(16'h13993,4);
TASK_PP(16'h13994,4);
TASK_PP(16'h13995,4);
TASK_PP(16'h13996,4);
TASK_PP(16'h13997,4);
TASK_PP(16'h13998,4);
TASK_PP(16'h13999,4);
TASK_PP(16'h1399A,4);
TASK_PP(16'h1399B,4);
TASK_PP(16'h1399C,4);
TASK_PP(16'h1399D,4);
TASK_PP(16'h1399E,4);
TASK_PP(16'h1399F,4);
TASK_PP(16'h139A0,4);
TASK_PP(16'h139A1,4);
TASK_PP(16'h139A2,4);
TASK_PP(16'h139A3,4);
TASK_PP(16'h139A4,4);
TASK_PP(16'h139A5,4);
TASK_PP(16'h139A6,4);
TASK_PP(16'h139A7,4);
TASK_PP(16'h139A8,4);
TASK_PP(16'h139A9,4);
TASK_PP(16'h139AA,4);
TASK_PP(16'h139AB,4);
TASK_PP(16'h139AC,4);
TASK_PP(16'h139AD,4);
TASK_PP(16'h139AE,4);
TASK_PP(16'h139AF,4);
TASK_PP(16'h139B0,4);
TASK_PP(16'h139B1,4);
TASK_PP(16'h139B2,4);
TASK_PP(16'h139B3,4);
TASK_PP(16'h139B4,4);
TASK_PP(16'h139B5,4);
TASK_PP(16'h139B6,4);
TASK_PP(16'h139B7,4);
TASK_PP(16'h139B8,4);
TASK_PP(16'h139B9,4);
TASK_PP(16'h139BA,4);
TASK_PP(16'h139BB,4);
TASK_PP(16'h139BC,4);
TASK_PP(16'h139BD,4);
TASK_PP(16'h139BE,4);
TASK_PP(16'h139BF,4);
TASK_PP(16'h139C0,4);
TASK_PP(16'h139C1,4);
TASK_PP(16'h139C2,4);
TASK_PP(16'h139C3,4);
TASK_PP(16'h139C4,4);
TASK_PP(16'h139C5,4);
TASK_PP(16'h139C6,4);
TASK_PP(16'h139C7,4);
TASK_PP(16'h139C8,4);
TASK_PP(16'h139C9,4);
TASK_PP(16'h139CA,4);
TASK_PP(16'h139CB,4);
TASK_PP(16'h139CC,4);
TASK_PP(16'h139CD,4);
TASK_PP(16'h139CE,4);
TASK_PP(16'h139CF,4);
TASK_PP(16'h139D0,4);
TASK_PP(16'h139D1,4);
TASK_PP(16'h139D2,4);
TASK_PP(16'h139D3,4);
TASK_PP(16'h139D4,4);
TASK_PP(16'h139D5,4);
TASK_PP(16'h139D6,4);
TASK_PP(16'h139D7,4);
TASK_PP(16'h139D8,4);
TASK_PP(16'h139D9,4);
TASK_PP(16'h139DA,4);
TASK_PP(16'h139DB,4);
TASK_PP(16'h139DC,4);
TASK_PP(16'h139DD,4);
TASK_PP(16'h139DE,4);
TASK_PP(16'h139DF,4);
TASK_PP(16'h139E0,4);
TASK_PP(16'h139E1,4);
TASK_PP(16'h139E2,4);
TASK_PP(16'h139E3,4);
TASK_PP(16'h139E4,4);
TASK_PP(16'h139E5,4);
TASK_PP(16'h139E6,4);
TASK_PP(16'h139E7,4);
TASK_PP(16'h139E8,4);
TASK_PP(16'h139E9,4);
TASK_PP(16'h139EA,4);
TASK_PP(16'h139EB,4);
TASK_PP(16'h139EC,4);
TASK_PP(16'h139ED,4);
TASK_PP(16'h139EE,4);
TASK_PP(16'h139EF,4);
TASK_PP(16'h139F0,4);
TASK_PP(16'h139F1,4);
TASK_PP(16'h139F2,4);
TASK_PP(16'h139F3,4);
TASK_PP(16'h139F4,4);
TASK_PP(16'h139F5,4);
TASK_PP(16'h139F6,4);
TASK_PP(16'h139F7,4);
TASK_PP(16'h139F8,4);
TASK_PP(16'h139F9,4);
TASK_PP(16'h139FA,4);
TASK_PP(16'h139FB,4);
TASK_PP(16'h139FC,4);
TASK_PP(16'h139FD,4);
TASK_PP(16'h139FE,4);
TASK_PP(16'h139FF,4);
TASK_PP(16'h13A00,4);
TASK_PP(16'h13A01,4);
TASK_PP(16'h13A02,4);
TASK_PP(16'h13A03,4);
TASK_PP(16'h13A04,4);
TASK_PP(16'h13A05,4);
TASK_PP(16'h13A06,4);
TASK_PP(16'h13A07,4);
TASK_PP(16'h13A08,4);
TASK_PP(16'h13A09,4);
TASK_PP(16'h13A0A,4);
TASK_PP(16'h13A0B,4);
TASK_PP(16'h13A0C,4);
TASK_PP(16'h13A0D,4);
TASK_PP(16'h13A0E,4);
TASK_PP(16'h13A0F,4);
TASK_PP(16'h13A10,4);
TASK_PP(16'h13A11,4);
TASK_PP(16'h13A12,4);
TASK_PP(16'h13A13,4);
TASK_PP(16'h13A14,4);
TASK_PP(16'h13A15,4);
TASK_PP(16'h13A16,4);
TASK_PP(16'h13A17,4);
TASK_PP(16'h13A18,4);
TASK_PP(16'h13A19,4);
TASK_PP(16'h13A1A,4);
TASK_PP(16'h13A1B,4);
TASK_PP(16'h13A1C,4);
TASK_PP(16'h13A1D,4);
TASK_PP(16'h13A1E,4);
TASK_PP(16'h13A1F,4);
TASK_PP(16'h13A20,4);
TASK_PP(16'h13A21,4);
TASK_PP(16'h13A22,4);
TASK_PP(16'h13A23,4);
TASK_PP(16'h13A24,4);
TASK_PP(16'h13A25,4);
TASK_PP(16'h13A26,4);
TASK_PP(16'h13A27,4);
TASK_PP(16'h13A28,4);
TASK_PP(16'h13A29,4);
TASK_PP(16'h13A2A,4);
TASK_PP(16'h13A2B,4);
TASK_PP(16'h13A2C,4);
TASK_PP(16'h13A2D,4);
TASK_PP(16'h13A2E,4);
TASK_PP(16'h13A2F,4);
TASK_PP(16'h13A30,4);
TASK_PP(16'h13A31,4);
TASK_PP(16'h13A32,4);
TASK_PP(16'h13A33,4);
TASK_PP(16'h13A34,4);
TASK_PP(16'h13A35,4);
TASK_PP(16'h13A36,4);
TASK_PP(16'h13A37,4);
TASK_PP(16'h13A38,4);
TASK_PP(16'h13A39,4);
TASK_PP(16'h13A3A,4);
TASK_PP(16'h13A3B,4);
TASK_PP(16'h13A3C,4);
TASK_PP(16'h13A3D,4);
TASK_PP(16'h13A3E,4);
TASK_PP(16'h13A3F,4);
TASK_PP(16'h13A40,4);
TASK_PP(16'h13A41,4);
TASK_PP(16'h13A42,4);
TASK_PP(16'h13A43,4);
TASK_PP(16'h13A44,4);
TASK_PP(16'h13A45,4);
TASK_PP(16'h13A46,4);
TASK_PP(16'h13A47,4);
TASK_PP(16'h13A48,4);
TASK_PP(16'h13A49,4);
TASK_PP(16'h13A4A,4);
TASK_PP(16'h13A4B,4);
TASK_PP(16'h13A4C,4);
TASK_PP(16'h13A4D,4);
TASK_PP(16'h13A4E,4);
TASK_PP(16'h13A4F,4);
TASK_PP(16'h13A50,4);
TASK_PP(16'h13A51,4);
TASK_PP(16'h13A52,4);
TASK_PP(16'h13A53,4);
TASK_PP(16'h13A54,4);
TASK_PP(16'h13A55,4);
TASK_PP(16'h13A56,4);
TASK_PP(16'h13A57,4);
TASK_PP(16'h13A58,4);
TASK_PP(16'h13A59,4);
TASK_PP(16'h13A5A,4);
TASK_PP(16'h13A5B,4);
TASK_PP(16'h13A5C,4);
TASK_PP(16'h13A5D,4);
TASK_PP(16'h13A5E,4);
TASK_PP(16'h13A5F,4);
TASK_PP(16'h13A60,4);
TASK_PP(16'h13A61,4);
TASK_PP(16'h13A62,4);
TASK_PP(16'h13A63,4);
TASK_PP(16'h13A64,4);
TASK_PP(16'h13A65,4);
TASK_PP(16'h13A66,4);
TASK_PP(16'h13A67,4);
TASK_PP(16'h13A68,4);
TASK_PP(16'h13A69,4);
TASK_PP(16'h13A6A,4);
TASK_PP(16'h13A6B,4);
TASK_PP(16'h13A6C,4);
TASK_PP(16'h13A6D,4);
TASK_PP(16'h13A6E,4);
TASK_PP(16'h13A6F,4);
TASK_PP(16'h13A70,4);
TASK_PP(16'h13A71,4);
TASK_PP(16'h13A72,4);
TASK_PP(16'h13A73,4);
TASK_PP(16'h13A74,4);
TASK_PP(16'h13A75,4);
TASK_PP(16'h13A76,4);
TASK_PP(16'h13A77,4);
TASK_PP(16'h13A78,4);
TASK_PP(16'h13A79,4);
TASK_PP(16'h13A7A,4);
TASK_PP(16'h13A7B,4);
TASK_PP(16'h13A7C,4);
TASK_PP(16'h13A7D,4);
TASK_PP(16'h13A7E,4);
TASK_PP(16'h13A7F,4);
TASK_PP(16'h13A80,4);
TASK_PP(16'h13A81,4);
TASK_PP(16'h13A82,4);
TASK_PP(16'h13A83,4);
TASK_PP(16'h13A84,4);
TASK_PP(16'h13A85,4);
TASK_PP(16'h13A86,4);
TASK_PP(16'h13A87,4);
TASK_PP(16'h13A88,4);
TASK_PP(16'h13A89,4);
TASK_PP(16'h13A8A,4);
TASK_PP(16'h13A8B,4);
TASK_PP(16'h13A8C,4);
TASK_PP(16'h13A8D,4);
TASK_PP(16'h13A8E,4);
TASK_PP(16'h13A8F,4);
TASK_PP(16'h13A90,4);
TASK_PP(16'h13A91,4);
TASK_PP(16'h13A92,4);
TASK_PP(16'h13A93,4);
TASK_PP(16'h13A94,4);
TASK_PP(16'h13A95,4);
TASK_PP(16'h13A96,4);
TASK_PP(16'h13A97,4);
TASK_PP(16'h13A98,4);
TASK_PP(16'h13A99,4);
TASK_PP(16'h13A9A,4);
TASK_PP(16'h13A9B,4);
TASK_PP(16'h13A9C,4);
TASK_PP(16'h13A9D,4);
TASK_PP(16'h13A9E,4);
TASK_PP(16'h13A9F,4);
TASK_PP(16'h13AA0,4);
TASK_PP(16'h13AA1,4);
TASK_PP(16'h13AA2,4);
TASK_PP(16'h13AA3,4);
TASK_PP(16'h13AA4,4);
TASK_PP(16'h13AA5,4);
TASK_PP(16'h13AA6,4);
TASK_PP(16'h13AA7,4);
TASK_PP(16'h13AA8,4);
TASK_PP(16'h13AA9,4);
TASK_PP(16'h13AAA,4);
TASK_PP(16'h13AAB,4);
TASK_PP(16'h13AAC,4);
TASK_PP(16'h13AAD,4);
TASK_PP(16'h13AAE,4);
TASK_PP(16'h13AAF,4);
TASK_PP(16'h13AB0,4);
TASK_PP(16'h13AB1,4);
TASK_PP(16'h13AB2,4);
TASK_PP(16'h13AB3,4);
TASK_PP(16'h13AB4,4);
TASK_PP(16'h13AB5,4);
TASK_PP(16'h13AB6,4);
TASK_PP(16'h13AB7,4);
TASK_PP(16'h13AB8,4);
TASK_PP(16'h13AB9,4);
TASK_PP(16'h13ABA,4);
TASK_PP(16'h13ABB,4);
TASK_PP(16'h13ABC,4);
TASK_PP(16'h13ABD,4);
TASK_PP(16'h13ABE,4);
TASK_PP(16'h13ABF,4);
TASK_PP(16'h13AC0,4);
TASK_PP(16'h13AC1,4);
TASK_PP(16'h13AC2,4);
TASK_PP(16'h13AC3,4);
TASK_PP(16'h13AC4,4);
TASK_PP(16'h13AC5,4);
TASK_PP(16'h13AC6,4);
TASK_PP(16'h13AC7,4);
TASK_PP(16'h13AC8,4);
TASK_PP(16'h13AC9,4);
TASK_PP(16'h13ACA,4);
TASK_PP(16'h13ACB,4);
TASK_PP(16'h13ACC,4);
TASK_PP(16'h13ACD,4);
TASK_PP(16'h13ACE,4);
TASK_PP(16'h13ACF,4);
TASK_PP(16'h13AD0,4);
TASK_PP(16'h13AD1,4);
TASK_PP(16'h13AD2,4);
TASK_PP(16'h13AD3,4);
TASK_PP(16'h13AD4,4);
TASK_PP(16'h13AD5,4);
TASK_PP(16'h13AD6,4);
TASK_PP(16'h13AD7,4);
TASK_PP(16'h13AD8,4);
TASK_PP(16'h13AD9,4);
TASK_PP(16'h13ADA,4);
TASK_PP(16'h13ADB,4);
TASK_PP(16'h13ADC,4);
TASK_PP(16'h13ADD,4);
TASK_PP(16'h13ADE,4);
TASK_PP(16'h13ADF,4);
TASK_PP(16'h13AE0,4);
TASK_PP(16'h13AE1,4);
TASK_PP(16'h13AE2,4);
TASK_PP(16'h13AE3,4);
TASK_PP(16'h13AE4,4);
TASK_PP(16'h13AE5,4);
TASK_PP(16'h13AE6,4);
TASK_PP(16'h13AE7,4);
TASK_PP(16'h13AE8,4);
TASK_PP(16'h13AE9,4);
TASK_PP(16'h13AEA,4);
TASK_PP(16'h13AEB,4);
TASK_PP(16'h13AEC,4);
TASK_PP(16'h13AED,4);
TASK_PP(16'h13AEE,4);
TASK_PP(16'h13AEF,4);
TASK_PP(16'h13AF0,4);
TASK_PP(16'h13AF1,4);
TASK_PP(16'h13AF2,4);
TASK_PP(16'h13AF3,4);
TASK_PP(16'h13AF4,4);
TASK_PP(16'h13AF5,4);
TASK_PP(16'h13AF6,4);
TASK_PP(16'h13AF7,4);
TASK_PP(16'h13AF8,4);
TASK_PP(16'h13AF9,4);
TASK_PP(16'h13AFA,4);
TASK_PP(16'h13AFB,4);
TASK_PP(16'h13AFC,4);
TASK_PP(16'h13AFD,4);
TASK_PP(16'h13AFE,4);
TASK_PP(16'h13AFF,4);
TASK_PP(16'h13B00,4);
TASK_PP(16'h13B01,4);
TASK_PP(16'h13B02,4);
TASK_PP(16'h13B03,4);
TASK_PP(16'h13B04,4);
TASK_PP(16'h13B05,4);
TASK_PP(16'h13B06,4);
TASK_PP(16'h13B07,4);
TASK_PP(16'h13B08,4);
TASK_PP(16'h13B09,4);
TASK_PP(16'h13B0A,4);
TASK_PP(16'h13B0B,4);
TASK_PP(16'h13B0C,4);
TASK_PP(16'h13B0D,4);
TASK_PP(16'h13B0E,4);
TASK_PP(16'h13B0F,4);
TASK_PP(16'h13B10,4);
TASK_PP(16'h13B11,4);
TASK_PP(16'h13B12,4);
TASK_PP(16'h13B13,4);
TASK_PP(16'h13B14,4);
TASK_PP(16'h13B15,4);
TASK_PP(16'h13B16,4);
TASK_PP(16'h13B17,4);
TASK_PP(16'h13B18,4);
TASK_PP(16'h13B19,4);
TASK_PP(16'h13B1A,4);
TASK_PP(16'h13B1B,4);
TASK_PP(16'h13B1C,4);
TASK_PP(16'h13B1D,4);
TASK_PP(16'h13B1E,4);
TASK_PP(16'h13B1F,4);
TASK_PP(16'h13B20,4);
TASK_PP(16'h13B21,4);
TASK_PP(16'h13B22,4);
TASK_PP(16'h13B23,4);
TASK_PP(16'h13B24,4);
TASK_PP(16'h13B25,4);
TASK_PP(16'h13B26,4);
TASK_PP(16'h13B27,4);
TASK_PP(16'h13B28,4);
TASK_PP(16'h13B29,4);
TASK_PP(16'h13B2A,4);
TASK_PP(16'h13B2B,4);
TASK_PP(16'h13B2C,4);
TASK_PP(16'h13B2D,4);
TASK_PP(16'h13B2E,4);
TASK_PP(16'h13B2F,4);
TASK_PP(16'h13B30,4);
TASK_PP(16'h13B31,4);
TASK_PP(16'h13B32,4);
TASK_PP(16'h13B33,4);
TASK_PP(16'h13B34,4);
TASK_PP(16'h13B35,4);
TASK_PP(16'h13B36,4);
TASK_PP(16'h13B37,4);
TASK_PP(16'h13B38,4);
TASK_PP(16'h13B39,4);
TASK_PP(16'h13B3A,4);
TASK_PP(16'h13B3B,4);
TASK_PP(16'h13B3C,4);
TASK_PP(16'h13B3D,4);
TASK_PP(16'h13B3E,4);
TASK_PP(16'h13B3F,4);
TASK_PP(16'h13B40,4);
TASK_PP(16'h13B41,4);
TASK_PP(16'h13B42,4);
TASK_PP(16'h13B43,4);
TASK_PP(16'h13B44,4);
TASK_PP(16'h13B45,4);
TASK_PP(16'h13B46,4);
TASK_PP(16'h13B47,4);
TASK_PP(16'h13B48,4);
TASK_PP(16'h13B49,4);
TASK_PP(16'h13B4A,4);
TASK_PP(16'h13B4B,4);
TASK_PP(16'h13B4C,4);
TASK_PP(16'h13B4D,4);
TASK_PP(16'h13B4E,4);
TASK_PP(16'h13B4F,4);
TASK_PP(16'h13B50,4);
TASK_PP(16'h13B51,4);
TASK_PP(16'h13B52,4);
TASK_PP(16'h13B53,4);
TASK_PP(16'h13B54,4);
TASK_PP(16'h13B55,4);
TASK_PP(16'h13B56,4);
TASK_PP(16'h13B57,4);
TASK_PP(16'h13B58,4);
TASK_PP(16'h13B59,4);
TASK_PP(16'h13B5A,4);
TASK_PP(16'h13B5B,4);
TASK_PP(16'h13B5C,4);
TASK_PP(16'h13B5D,4);
TASK_PP(16'h13B5E,4);
TASK_PP(16'h13B5F,4);
TASK_PP(16'h13B60,4);
TASK_PP(16'h13B61,4);
TASK_PP(16'h13B62,4);
TASK_PP(16'h13B63,4);
TASK_PP(16'h13B64,4);
TASK_PP(16'h13B65,4);
TASK_PP(16'h13B66,4);
TASK_PP(16'h13B67,4);
TASK_PP(16'h13B68,4);
TASK_PP(16'h13B69,4);
TASK_PP(16'h13B6A,4);
TASK_PP(16'h13B6B,4);
TASK_PP(16'h13B6C,4);
TASK_PP(16'h13B6D,4);
TASK_PP(16'h13B6E,4);
TASK_PP(16'h13B6F,4);
TASK_PP(16'h13B70,4);
TASK_PP(16'h13B71,4);
TASK_PP(16'h13B72,4);
TASK_PP(16'h13B73,4);
TASK_PP(16'h13B74,4);
TASK_PP(16'h13B75,4);
TASK_PP(16'h13B76,4);
TASK_PP(16'h13B77,4);
TASK_PP(16'h13B78,4);
TASK_PP(16'h13B79,4);
TASK_PP(16'h13B7A,4);
TASK_PP(16'h13B7B,4);
TASK_PP(16'h13B7C,4);
TASK_PP(16'h13B7D,4);
TASK_PP(16'h13B7E,4);
TASK_PP(16'h13B7F,4);
TASK_PP(16'h13B80,4);
TASK_PP(16'h13B81,4);
TASK_PP(16'h13B82,4);
TASK_PP(16'h13B83,4);
TASK_PP(16'h13B84,4);
TASK_PP(16'h13B85,4);
TASK_PP(16'h13B86,4);
TASK_PP(16'h13B87,4);
TASK_PP(16'h13B88,4);
TASK_PP(16'h13B89,4);
TASK_PP(16'h13B8A,4);
TASK_PP(16'h13B8B,4);
TASK_PP(16'h13B8C,4);
TASK_PP(16'h13B8D,4);
TASK_PP(16'h13B8E,4);
TASK_PP(16'h13B8F,4);
TASK_PP(16'h13B90,4);
TASK_PP(16'h13B91,4);
TASK_PP(16'h13B92,4);
TASK_PP(16'h13B93,4);
TASK_PP(16'h13B94,4);
TASK_PP(16'h13B95,4);
TASK_PP(16'h13B96,4);
TASK_PP(16'h13B97,4);
TASK_PP(16'h13B98,4);
TASK_PP(16'h13B99,4);
TASK_PP(16'h13B9A,4);
TASK_PP(16'h13B9B,4);
TASK_PP(16'h13B9C,4);
TASK_PP(16'h13B9D,4);
TASK_PP(16'h13B9E,4);
TASK_PP(16'h13B9F,4);
TASK_PP(16'h13BA0,4);
TASK_PP(16'h13BA1,4);
TASK_PP(16'h13BA2,4);
TASK_PP(16'h13BA3,4);
TASK_PP(16'h13BA4,4);
TASK_PP(16'h13BA5,4);
TASK_PP(16'h13BA6,4);
TASK_PP(16'h13BA7,4);
TASK_PP(16'h13BA8,4);
TASK_PP(16'h13BA9,4);
TASK_PP(16'h13BAA,4);
TASK_PP(16'h13BAB,4);
TASK_PP(16'h13BAC,4);
TASK_PP(16'h13BAD,4);
TASK_PP(16'h13BAE,4);
TASK_PP(16'h13BAF,4);
TASK_PP(16'h13BB0,4);
TASK_PP(16'h13BB1,4);
TASK_PP(16'h13BB2,4);
TASK_PP(16'h13BB3,4);
TASK_PP(16'h13BB4,4);
TASK_PP(16'h13BB5,4);
TASK_PP(16'h13BB6,4);
TASK_PP(16'h13BB7,4);
TASK_PP(16'h13BB8,4);
TASK_PP(16'h13BB9,4);
TASK_PP(16'h13BBA,4);
TASK_PP(16'h13BBB,4);
TASK_PP(16'h13BBC,4);
TASK_PP(16'h13BBD,4);
TASK_PP(16'h13BBE,4);
TASK_PP(16'h13BBF,4);
TASK_PP(16'h13BC0,4);
TASK_PP(16'h13BC1,4);
TASK_PP(16'h13BC2,4);
TASK_PP(16'h13BC3,4);
TASK_PP(16'h13BC4,4);
TASK_PP(16'h13BC5,4);
TASK_PP(16'h13BC6,4);
TASK_PP(16'h13BC7,4);
TASK_PP(16'h13BC8,4);
TASK_PP(16'h13BC9,4);
TASK_PP(16'h13BCA,4);
TASK_PP(16'h13BCB,4);
TASK_PP(16'h13BCC,4);
TASK_PP(16'h13BCD,4);
TASK_PP(16'h13BCE,4);
TASK_PP(16'h13BCF,4);
TASK_PP(16'h13BD0,4);
TASK_PP(16'h13BD1,4);
TASK_PP(16'h13BD2,4);
TASK_PP(16'h13BD3,4);
TASK_PP(16'h13BD4,4);
TASK_PP(16'h13BD5,4);
TASK_PP(16'h13BD6,4);
TASK_PP(16'h13BD7,4);
TASK_PP(16'h13BD8,4);
TASK_PP(16'h13BD9,4);
TASK_PP(16'h13BDA,4);
TASK_PP(16'h13BDB,4);
TASK_PP(16'h13BDC,4);
TASK_PP(16'h13BDD,4);
TASK_PP(16'h13BDE,4);
TASK_PP(16'h13BDF,4);
TASK_PP(16'h13BE0,4);
TASK_PP(16'h13BE1,4);
TASK_PP(16'h13BE2,4);
TASK_PP(16'h13BE3,4);
TASK_PP(16'h13BE4,4);
TASK_PP(16'h13BE5,4);
TASK_PP(16'h13BE6,4);
TASK_PP(16'h13BE7,4);
TASK_PP(16'h13BE8,4);
TASK_PP(16'h13BE9,4);
TASK_PP(16'h13BEA,4);
TASK_PP(16'h13BEB,4);
TASK_PP(16'h13BEC,4);
TASK_PP(16'h13BED,4);
TASK_PP(16'h13BEE,4);
TASK_PP(16'h13BEF,4);
TASK_PP(16'h13BF0,4);
TASK_PP(16'h13BF1,4);
TASK_PP(16'h13BF2,4);
TASK_PP(16'h13BF3,4);
TASK_PP(16'h13BF4,4);
TASK_PP(16'h13BF5,4);
TASK_PP(16'h13BF6,4);
TASK_PP(16'h13BF7,4);
TASK_PP(16'h13BF8,4);
TASK_PP(16'h13BF9,4);
TASK_PP(16'h13BFA,4);
TASK_PP(16'h13BFB,4);
TASK_PP(16'h13BFC,4);
TASK_PP(16'h13BFD,4);
TASK_PP(16'h13BFE,4);
TASK_PP(16'h13BFF,4);
TASK_PP(16'h13C00,4);
TASK_PP(16'h13C01,4);
TASK_PP(16'h13C02,4);
TASK_PP(16'h13C03,4);
TASK_PP(16'h13C04,4);
TASK_PP(16'h13C05,4);
TASK_PP(16'h13C06,4);
TASK_PP(16'h13C07,4);
TASK_PP(16'h13C08,4);
TASK_PP(16'h13C09,4);
TASK_PP(16'h13C0A,4);
TASK_PP(16'h13C0B,4);
TASK_PP(16'h13C0C,4);
TASK_PP(16'h13C0D,4);
TASK_PP(16'h13C0E,4);
TASK_PP(16'h13C0F,4);
TASK_PP(16'h13C10,4);
TASK_PP(16'h13C11,4);
TASK_PP(16'h13C12,4);
TASK_PP(16'h13C13,4);
TASK_PP(16'h13C14,4);
TASK_PP(16'h13C15,4);
TASK_PP(16'h13C16,4);
TASK_PP(16'h13C17,4);
TASK_PP(16'h13C18,4);
TASK_PP(16'h13C19,4);
TASK_PP(16'h13C1A,4);
TASK_PP(16'h13C1B,4);
TASK_PP(16'h13C1C,4);
TASK_PP(16'h13C1D,4);
TASK_PP(16'h13C1E,4);
TASK_PP(16'h13C1F,4);
TASK_PP(16'h13C20,4);
TASK_PP(16'h13C21,4);
TASK_PP(16'h13C22,4);
TASK_PP(16'h13C23,4);
TASK_PP(16'h13C24,4);
TASK_PP(16'h13C25,4);
TASK_PP(16'h13C26,4);
TASK_PP(16'h13C27,4);
TASK_PP(16'h13C28,4);
TASK_PP(16'h13C29,4);
TASK_PP(16'h13C2A,4);
TASK_PP(16'h13C2B,4);
TASK_PP(16'h13C2C,4);
TASK_PP(16'h13C2D,4);
TASK_PP(16'h13C2E,4);
TASK_PP(16'h13C2F,4);
TASK_PP(16'h13C30,4);
TASK_PP(16'h13C31,4);
TASK_PP(16'h13C32,4);
TASK_PP(16'h13C33,4);
TASK_PP(16'h13C34,4);
TASK_PP(16'h13C35,4);
TASK_PP(16'h13C36,4);
TASK_PP(16'h13C37,4);
TASK_PP(16'h13C38,4);
TASK_PP(16'h13C39,4);
TASK_PP(16'h13C3A,4);
TASK_PP(16'h13C3B,4);
TASK_PP(16'h13C3C,4);
TASK_PP(16'h13C3D,4);
TASK_PP(16'h13C3E,4);
TASK_PP(16'h13C3F,4);
TASK_PP(16'h13C40,4);
TASK_PP(16'h13C41,4);
TASK_PP(16'h13C42,4);
TASK_PP(16'h13C43,4);
TASK_PP(16'h13C44,4);
TASK_PP(16'h13C45,4);
TASK_PP(16'h13C46,4);
TASK_PP(16'h13C47,4);
TASK_PP(16'h13C48,4);
TASK_PP(16'h13C49,4);
TASK_PP(16'h13C4A,4);
TASK_PP(16'h13C4B,4);
TASK_PP(16'h13C4C,4);
TASK_PP(16'h13C4D,4);
TASK_PP(16'h13C4E,4);
TASK_PP(16'h13C4F,4);
TASK_PP(16'h13C50,4);
TASK_PP(16'h13C51,4);
TASK_PP(16'h13C52,4);
TASK_PP(16'h13C53,4);
TASK_PP(16'h13C54,4);
TASK_PP(16'h13C55,4);
TASK_PP(16'h13C56,4);
TASK_PP(16'h13C57,4);
TASK_PP(16'h13C58,4);
TASK_PP(16'h13C59,4);
TASK_PP(16'h13C5A,4);
TASK_PP(16'h13C5B,4);
TASK_PP(16'h13C5C,4);
TASK_PP(16'h13C5D,4);
TASK_PP(16'h13C5E,4);
TASK_PP(16'h13C5F,4);
TASK_PP(16'h13C60,4);
TASK_PP(16'h13C61,4);
TASK_PP(16'h13C62,4);
TASK_PP(16'h13C63,4);
TASK_PP(16'h13C64,4);
TASK_PP(16'h13C65,4);
TASK_PP(16'h13C66,4);
TASK_PP(16'h13C67,4);
TASK_PP(16'h13C68,4);
TASK_PP(16'h13C69,4);
TASK_PP(16'h13C6A,4);
TASK_PP(16'h13C6B,4);
TASK_PP(16'h13C6C,4);
TASK_PP(16'h13C6D,4);
TASK_PP(16'h13C6E,4);
TASK_PP(16'h13C6F,4);
TASK_PP(16'h13C70,4);
TASK_PP(16'h13C71,4);
TASK_PP(16'h13C72,4);
TASK_PP(16'h13C73,4);
TASK_PP(16'h13C74,4);
TASK_PP(16'h13C75,4);
TASK_PP(16'h13C76,4);
TASK_PP(16'h13C77,4);
TASK_PP(16'h13C78,4);
TASK_PP(16'h13C79,4);
TASK_PP(16'h13C7A,4);
TASK_PP(16'h13C7B,4);
TASK_PP(16'h13C7C,4);
TASK_PP(16'h13C7D,4);
TASK_PP(16'h13C7E,4);
TASK_PP(16'h13C7F,4);
TASK_PP(16'h13C80,4);
TASK_PP(16'h13C81,4);
TASK_PP(16'h13C82,4);
TASK_PP(16'h13C83,4);
TASK_PP(16'h13C84,4);
TASK_PP(16'h13C85,4);
TASK_PP(16'h13C86,4);
TASK_PP(16'h13C87,4);
TASK_PP(16'h13C88,4);
TASK_PP(16'h13C89,4);
TASK_PP(16'h13C8A,4);
TASK_PP(16'h13C8B,4);
TASK_PP(16'h13C8C,4);
TASK_PP(16'h13C8D,4);
TASK_PP(16'h13C8E,4);
TASK_PP(16'h13C8F,4);
TASK_PP(16'h13C90,4);
TASK_PP(16'h13C91,4);
TASK_PP(16'h13C92,4);
TASK_PP(16'h13C93,4);
TASK_PP(16'h13C94,4);
TASK_PP(16'h13C95,4);
TASK_PP(16'h13C96,4);
TASK_PP(16'h13C97,4);
TASK_PP(16'h13C98,4);
TASK_PP(16'h13C99,4);
TASK_PP(16'h13C9A,4);
TASK_PP(16'h13C9B,4);
TASK_PP(16'h13C9C,4);
TASK_PP(16'h13C9D,4);
TASK_PP(16'h13C9E,4);
TASK_PP(16'h13C9F,4);
TASK_PP(16'h13CA0,4);
TASK_PP(16'h13CA1,4);
TASK_PP(16'h13CA2,4);
TASK_PP(16'h13CA3,4);
TASK_PP(16'h13CA4,4);
TASK_PP(16'h13CA5,4);
TASK_PP(16'h13CA6,4);
TASK_PP(16'h13CA7,4);
TASK_PP(16'h13CA8,4);
TASK_PP(16'h13CA9,4);
TASK_PP(16'h13CAA,4);
TASK_PP(16'h13CAB,4);
TASK_PP(16'h13CAC,4);
TASK_PP(16'h13CAD,4);
TASK_PP(16'h13CAE,4);
TASK_PP(16'h13CAF,4);
TASK_PP(16'h13CB0,4);
TASK_PP(16'h13CB1,4);
TASK_PP(16'h13CB2,4);
TASK_PP(16'h13CB3,4);
TASK_PP(16'h13CB4,4);
TASK_PP(16'h13CB5,4);
TASK_PP(16'h13CB6,4);
TASK_PP(16'h13CB7,4);
TASK_PP(16'h13CB8,4);
TASK_PP(16'h13CB9,4);
TASK_PP(16'h13CBA,4);
TASK_PP(16'h13CBB,4);
TASK_PP(16'h13CBC,4);
TASK_PP(16'h13CBD,4);
TASK_PP(16'h13CBE,4);
TASK_PP(16'h13CBF,4);
TASK_PP(16'h13CC0,4);
TASK_PP(16'h13CC1,4);
TASK_PP(16'h13CC2,4);
TASK_PP(16'h13CC3,4);
TASK_PP(16'h13CC4,4);
TASK_PP(16'h13CC5,4);
TASK_PP(16'h13CC6,4);
TASK_PP(16'h13CC7,4);
TASK_PP(16'h13CC8,4);
TASK_PP(16'h13CC9,4);
TASK_PP(16'h13CCA,4);
TASK_PP(16'h13CCB,4);
TASK_PP(16'h13CCC,4);
TASK_PP(16'h13CCD,4);
TASK_PP(16'h13CCE,4);
TASK_PP(16'h13CCF,4);
TASK_PP(16'h13CD0,4);
TASK_PP(16'h13CD1,4);
TASK_PP(16'h13CD2,4);
TASK_PP(16'h13CD3,4);
TASK_PP(16'h13CD4,4);
TASK_PP(16'h13CD5,4);
TASK_PP(16'h13CD6,4);
TASK_PP(16'h13CD7,4);
TASK_PP(16'h13CD8,4);
TASK_PP(16'h13CD9,4);
TASK_PP(16'h13CDA,4);
TASK_PP(16'h13CDB,4);
TASK_PP(16'h13CDC,4);
TASK_PP(16'h13CDD,4);
TASK_PP(16'h13CDE,4);
TASK_PP(16'h13CDF,4);
TASK_PP(16'h13CE0,4);
TASK_PP(16'h13CE1,4);
TASK_PP(16'h13CE2,4);
TASK_PP(16'h13CE3,4);
TASK_PP(16'h13CE4,4);
TASK_PP(16'h13CE5,4);
TASK_PP(16'h13CE6,4);
TASK_PP(16'h13CE7,4);
TASK_PP(16'h13CE8,4);
TASK_PP(16'h13CE9,4);
TASK_PP(16'h13CEA,4);
TASK_PP(16'h13CEB,4);
TASK_PP(16'h13CEC,4);
TASK_PP(16'h13CED,4);
TASK_PP(16'h13CEE,4);
TASK_PP(16'h13CEF,4);
TASK_PP(16'h13CF0,4);
TASK_PP(16'h13CF1,4);
TASK_PP(16'h13CF2,4);
TASK_PP(16'h13CF3,4);
TASK_PP(16'h13CF4,4);
TASK_PP(16'h13CF5,4);
TASK_PP(16'h13CF6,4);
TASK_PP(16'h13CF7,4);
TASK_PP(16'h13CF8,4);
TASK_PP(16'h13CF9,4);
TASK_PP(16'h13CFA,4);
TASK_PP(16'h13CFB,4);
TASK_PP(16'h13CFC,4);
TASK_PP(16'h13CFD,4);
TASK_PP(16'h13CFE,4);
TASK_PP(16'h13CFF,4);
TASK_PP(16'h13D00,4);
TASK_PP(16'h13D01,4);
TASK_PP(16'h13D02,4);
TASK_PP(16'h13D03,4);
TASK_PP(16'h13D04,4);
TASK_PP(16'h13D05,4);
TASK_PP(16'h13D06,4);
TASK_PP(16'h13D07,4);
TASK_PP(16'h13D08,4);
TASK_PP(16'h13D09,4);
TASK_PP(16'h13D0A,4);
TASK_PP(16'h13D0B,4);
TASK_PP(16'h13D0C,4);
TASK_PP(16'h13D0D,4);
TASK_PP(16'h13D0E,4);
TASK_PP(16'h13D0F,4);
TASK_PP(16'h13D10,4);
TASK_PP(16'h13D11,4);
TASK_PP(16'h13D12,4);
TASK_PP(16'h13D13,4);
TASK_PP(16'h13D14,4);
TASK_PP(16'h13D15,4);
TASK_PP(16'h13D16,4);
TASK_PP(16'h13D17,4);
TASK_PP(16'h13D18,4);
TASK_PP(16'h13D19,4);
TASK_PP(16'h13D1A,4);
TASK_PP(16'h13D1B,4);
TASK_PP(16'h13D1C,4);
TASK_PP(16'h13D1D,4);
TASK_PP(16'h13D1E,4);
TASK_PP(16'h13D1F,4);
TASK_PP(16'h13D20,4);
TASK_PP(16'h13D21,4);
TASK_PP(16'h13D22,4);
TASK_PP(16'h13D23,4);
TASK_PP(16'h13D24,4);
TASK_PP(16'h13D25,4);
TASK_PP(16'h13D26,4);
TASK_PP(16'h13D27,4);
TASK_PP(16'h13D28,4);
TASK_PP(16'h13D29,4);
TASK_PP(16'h13D2A,4);
TASK_PP(16'h13D2B,4);
TASK_PP(16'h13D2C,4);
TASK_PP(16'h13D2D,4);
TASK_PP(16'h13D2E,4);
TASK_PP(16'h13D2F,4);
TASK_PP(16'h13D30,4);
TASK_PP(16'h13D31,4);
TASK_PP(16'h13D32,4);
TASK_PP(16'h13D33,4);
TASK_PP(16'h13D34,4);
TASK_PP(16'h13D35,4);
TASK_PP(16'h13D36,4);
TASK_PP(16'h13D37,4);
TASK_PP(16'h13D38,4);
TASK_PP(16'h13D39,4);
TASK_PP(16'h13D3A,4);
TASK_PP(16'h13D3B,4);
TASK_PP(16'h13D3C,4);
TASK_PP(16'h13D3D,4);
TASK_PP(16'h13D3E,4);
TASK_PP(16'h13D3F,4);
TASK_PP(16'h13D40,4);
TASK_PP(16'h13D41,4);
TASK_PP(16'h13D42,4);
TASK_PP(16'h13D43,4);
TASK_PP(16'h13D44,4);
TASK_PP(16'h13D45,4);
TASK_PP(16'h13D46,4);
TASK_PP(16'h13D47,4);
TASK_PP(16'h13D48,4);
TASK_PP(16'h13D49,4);
TASK_PP(16'h13D4A,4);
TASK_PP(16'h13D4B,4);
TASK_PP(16'h13D4C,4);
TASK_PP(16'h13D4D,4);
TASK_PP(16'h13D4E,4);
TASK_PP(16'h13D4F,4);
TASK_PP(16'h13D50,4);
TASK_PP(16'h13D51,4);
TASK_PP(16'h13D52,4);
TASK_PP(16'h13D53,4);
TASK_PP(16'h13D54,4);
TASK_PP(16'h13D55,4);
TASK_PP(16'h13D56,4);
TASK_PP(16'h13D57,4);
TASK_PP(16'h13D58,4);
TASK_PP(16'h13D59,4);
TASK_PP(16'h13D5A,4);
TASK_PP(16'h13D5B,4);
TASK_PP(16'h13D5C,4);
TASK_PP(16'h13D5D,4);
TASK_PP(16'h13D5E,4);
TASK_PP(16'h13D5F,4);
TASK_PP(16'h13D60,4);
TASK_PP(16'h13D61,4);
TASK_PP(16'h13D62,4);
TASK_PP(16'h13D63,4);
TASK_PP(16'h13D64,4);
TASK_PP(16'h13D65,4);
TASK_PP(16'h13D66,4);
TASK_PP(16'h13D67,4);
TASK_PP(16'h13D68,4);
TASK_PP(16'h13D69,4);
TASK_PP(16'h13D6A,4);
TASK_PP(16'h13D6B,4);
TASK_PP(16'h13D6C,4);
TASK_PP(16'h13D6D,4);
TASK_PP(16'h13D6E,4);
TASK_PP(16'h13D6F,4);
TASK_PP(16'h13D70,4);
TASK_PP(16'h13D71,4);
TASK_PP(16'h13D72,4);
TASK_PP(16'h13D73,4);
TASK_PP(16'h13D74,4);
TASK_PP(16'h13D75,4);
TASK_PP(16'h13D76,4);
TASK_PP(16'h13D77,4);
TASK_PP(16'h13D78,4);
TASK_PP(16'h13D79,4);
TASK_PP(16'h13D7A,4);
TASK_PP(16'h13D7B,4);
TASK_PP(16'h13D7C,4);
TASK_PP(16'h13D7D,4);
TASK_PP(16'h13D7E,4);
TASK_PP(16'h13D7F,4);
TASK_PP(16'h13D80,4);
TASK_PP(16'h13D81,4);
TASK_PP(16'h13D82,4);
TASK_PP(16'h13D83,4);
TASK_PP(16'h13D84,4);
TASK_PP(16'h13D85,4);
TASK_PP(16'h13D86,4);
TASK_PP(16'h13D87,4);
TASK_PP(16'h13D88,4);
TASK_PP(16'h13D89,4);
TASK_PP(16'h13D8A,4);
TASK_PP(16'h13D8B,4);
TASK_PP(16'h13D8C,4);
TASK_PP(16'h13D8D,4);
TASK_PP(16'h13D8E,4);
TASK_PP(16'h13D8F,4);
TASK_PP(16'h13D90,4);
TASK_PP(16'h13D91,4);
TASK_PP(16'h13D92,4);
TASK_PP(16'h13D93,4);
TASK_PP(16'h13D94,4);
TASK_PP(16'h13D95,4);
TASK_PP(16'h13D96,4);
TASK_PP(16'h13D97,4);
TASK_PP(16'h13D98,4);
TASK_PP(16'h13D99,4);
TASK_PP(16'h13D9A,4);
TASK_PP(16'h13D9B,4);
TASK_PP(16'h13D9C,4);
TASK_PP(16'h13D9D,4);
TASK_PP(16'h13D9E,4);
TASK_PP(16'h13D9F,4);
TASK_PP(16'h13DA0,4);
TASK_PP(16'h13DA1,4);
TASK_PP(16'h13DA2,4);
TASK_PP(16'h13DA3,4);
TASK_PP(16'h13DA4,4);
TASK_PP(16'h13DA5,4);
TASK_PP(16'h13DA6,4);
TASK_PP(16'h13DA7,4);
TASK_PP(16'h13DA8,4);
TASK_PP(16'h13DA9,4);
TASK_PP(16'h13DAA,4);
TASK_PP(16'h13DAB,4);
TASK_PP(16'h13DAC,4);
TASK_PP(16'h13DAD,4);
TASK_PP(16'h13DAE,4);
TASK_PP(16'h13DAF,4);
TASK_PP(16'h13DB0,4);
TASK_PP(16'h13DB1,4);
TASK_PP(16'h13DB2,4);
TASK_PP(16'h13DB3,4);
TASK_PP(16'h13DB4,4);
TASK_PP(16'h13DB5,4);
TASK_PP(16'h13DB6,4);
TASK_PP(16'h13DB7,4);
TASK_PP(16'h13DB8,4);
TASK_PP(16'h13DB9,4);
TASK_PP(16'h13DBA,4);
TASK_PP(16'h13DBB,4);
TASK_PP(16'h13DBC,4);
TASK_PP(16'h13DBD,4);
TASK_PP(16'h13DBE,4);
TASK_PP(16'h13DBF,4);
TASK_PP(16'h13DC0,4);
TASK_PP(16'h13DC1,4);
TASK_PP(16'h13DC2,4);
TASK_PP(16'h13DC3,4);
TASK_PP(16'h13DC4,4);
TASK_PP(16'h13DC5,4);
TASK_PP(16'h13DC6,4);
TASK_PP(16'h13DC7,4);
TASK_PP(16'h13DC8,4);
TASK_PP(16'h13DC9,4);
TASK_PP(16'h13DCA,4);
TASK_PP(16'h13DCB,4);
TASK_PP(16'h13DCC,4);
TASK_PP(16'h13DCD,4);
TASK_PP(16'h13DCE,4);
TASK_PP(16'h13DCF,4);
TASK_PP(16'h13DD0,4);
TASK_PP(16'h13DD1,4);
TASK_PP(16'h13DD2,4);
TASK_PP(16'h13DD3,4);
TASK_PP(16'h13DD4,4);
TASK_PP(16'h13DD5,4);
TASK_PP(16'h13DD6,4);
TASK_PP(16'h13DD7,4);
TASK_PP(16'h13DD8,4);
TASK_PP(16'h13DD9,4);
TASK_PP(16'h13DDA,4);
TASK_PP(16'h13DDB,4);
TASK_PP(16'h13DDC,4);
TASK_PP(16'h13DDD,4);
TASK_PP(16'h13DDE,4);
TASK_PP(16'h13DDF,4);
TASK_PP(16'h13DE0,4);
TASK_PP(16'h13DE1,4);
TASK_PP(16'h13DE2,4);
TASK_PP(16'h13DE3,4);
TASK_PP(16'h13DE4,4);
TASK_PP(16'h13DE5,4);
TASK_PP(16'h13DE6,4);
TASK_PP(16'h13DE7,4);
TASK_PP(16'h13DE8,4);
TASK_PP(16'h13DE9,4);
TASK_PP(16'h13DEA,4);
TASK_PP(16'h13DEB,4);
TASK_PP(16'h13DEC,4);
TASK_PP(16'h13DED,4);
TASK_PP(16'h13DEE,4);
TASK_PP(16'h13DEF,4);
TASK_PP(16'h13DF0,4);
TASK_PP(16'h13DF1,4);
TASK_PP(16'h13DF2,4);
TASK_PP(16'h13DF3,4);
TASK_PP(16'h13DF4,4);
TASK_PP(16'h13DF5,4);
TASK_PP(16'h13DF6,4);
TASK_PP(16'h13DF7,4);
TASK_PP(16'h13DF8,4);
TASK_PP(16'h13DF9,4);
TASK_PP(16'h13DFA,4);
TASK_PP(16'h13DFB,4);
TASK_PP(16'h13DFC,4);
TASK_PP(16'h13DFD,4);
TASK_PP(16'h13DFE,4);
TASK_PP(16'h13DFF,4);
TASK_PP(16'h13E00,4);
TASK_PP(16'h13E01,4);
TASK_PP(16'h13E02,4);
TASK_PP(16'h13E03,4);
TASK_PP(16'h13E04,4);
TASK_PP(16'h13E05,4);
TASK_PP(16'h13E06,4);
TASK_PP(16'h13E07,4);
TASK_PP(16'h13E08,4);
TASK_PP(16'h13E09,4);
TASK_PP(16'h13E0A,4);
TASK_PP(16'h13E0B,4);
TASK_PP(16'h13E0C,4);
TASK_PP(16'h13E0D,4);
TASK_PP(16'h13E0E,4);
TASK_PP(16'h13E0F,4);
TASK_PP(16'h13E10,4);
TASK_PP(16'h13E11,4);
TASK_PP(16'h13E12,4);
TASK_PP(16'h13E13,4);
TASK_PP(16'h13E14,4);
TASK_PP(16'h13E15,4);
TASK_PP(16'h13E16,4);
TASK_PP(16'h13E17,4);
TASK_PP(16'h13E18,4);
TASK_PP(16'h13E19,4);
TASK_PP(16'h13E1A,4);
TASK_PP(16'h13E1B,4);
TASK_PP(16'h13E1C,4);
TASK_PP(16'h13E1D,4);
TASK_PP(16'h13E1E,4);
TASK_PP(16'h13E1F,4);
TASK_PP(16'h13E20,4);
TASK_PP(16'h13E21,4);
TASK_PP(16'h13E22,4);
TASK_PP(16'h13E23,4);
TASK_PP(16'h13E24,4);
TASK_PP(16'h13E25,4);
TASK_PP(16'h13E26,4);
TASK_PP(16'h13E27,4);
TASK_PP(16'h13E28,4);
TASK_PP(16'h13E29,4);
TASK_PP(16'h13E2A,4);
TASK_PP(16'h13E2B,4);
TASK_PP(16'h13E2C,4);
TASK_PP(16'h13E2D,4);
TASK_PP(16'h13E2E,4);
TASK_PP(16'h13E2F,4);
TASK_PP(16'h13E30,4);
TASK_PP(16'h13E31,4);
TASK_PP(16'h13E32,4);
TASK_PP(16'h13E33,4);
TASK_PP(16'h13E34,4);
TASK_PP(16'h13E35,4);
TASK_PP(16'h13E36,4);
TASK_PP(16'h13E37,4);
TASK_PP(16'h13E38,4);
TASK_PP(16'h13E39,4);
TASK_PP(16'h13E3A,4);
TASK_PP(16'h13E3B,4);
TASK_PP(16'h13E3C,4);
TASK_PP(16'h13E3D,4);
TASK_PP(16'h13E3E,4);
TASK_PP(16'h13E3F,4);
TASK_PP(16'h13E40,4);
TASK_PP(16'h13E41,4);
TASK_PP(16'h13E42,4);
TASK_PP(16'h13E43,4);
TASK_PP(16'h13E44,4);
TASK_PP(16'h13E45,4);
TASK_PP(16'h13E46,4);
TASK_PP(16'h13E47,4);
TASK_PP(16'h13E48,4);
TASK_PP(16'h13E49,4);
TASK_PP(16'h13E4A,4);
TASK_PP(16'h13E4B,4);
TASK_PP(16'h13E4C,4);
TASK_PP(16'h13E4D,4);
TASK_PP(16'h13E4E,4);
TASK_PP(16'h13E4F,4);
TASK_PP(16'h13E50,4);
TASK_PP(16'h13E51,4);
TASK_PP(16'h13E52,4);
TASK_PP(16'h13E53,4);
TASK_PP(16'h13E54,4);
TASK_PP(16'h13E55,4);
TASK_PP(16'h13E56,4);
TASK_PP(16'h13E57,4);
TASK_PP(16'h13E58,4);
TASK_PP(16'h13E59,4);
TASK_PP(16'h13E5A,4);
TASK_PP(16'h13E5B,4);
TASK_PP(16'h13E5C,4);
TASK_PP(16'h13E5D,4);
TASK_PP(16'h13E5E,4);
TASK_PP(16'h13E5F,4);
TASK_PP(16'h13E60,4);
TASK_PP(16'h13E61,4);
TASK_PP(16'h13E62,4);
TASK_PP(16'h13E63,4);
TASK_PP(16'h13E64,4);
TASK_PP(16'h13E65,4);
TASK_PP(16'h13E66,4);
TASK_PP(16'h13E67,4);
TASK_PP(16'h13E68,4);
TASK_PP(16'h13E69,4);
TASK_PP(16'h13E6A,4);
TASK_PP(16'h13E6B,4);
TASK_PP(16'h13E6C,4);
TASK_PP(16'h13E6D,4);
TASK_PP(16'h13E6E,4);
TASK_PP(16'h13E6F,4);
TASK_PP(16'h13E70,4);
TASK_PP(16'h13E71,4);
TASK_PP(16'h13E72,4);
TASK_PP(16'h13E73,4);
TASK_PP(16'h13E74,4);
TASK_PP(16'h13E75,4);
TASK_PP(16'h13E76,4);
TASK_PP(16'h13E77,4);
TASK_PP(16'h13E78,4);
TASK_PP(16'h13E79,4);
TASK_PP(16'h13E7A,4);
TASK_PP(16'h13E7B,4);
TASK_PP(16'h13E7C,4);
TASK_PP(16'h13E7D,4);
TASK_PP(16'h13E7E,4);
TASK_PP(16'h13E7F,4);
TASK_PP(16'h13E80,4);
TASK_PP(16'h13E81,4);
TASK_PP(16'h13E82,4);
TASK_PP(16'h13E83,4);
TASK_PP(16'h13E84,4);
TASK_PP(16'h13E85,4);
TASK_PP(16'h13E86,4);
TASK_PP(16'h13E87,4);
TASK_PP(16'h13E88,4);
TASK_PP(16'h13E89,4);
TASK_PP(16'h13E8A,4);
TASK_PP(16'h13E8B,4);
TASK_PP(16'h13E8C,4);
TASK_PP(16'h13E8D,4);
TASK_PP(16'h13E8E,4);
TASK_PP(16'h13E8F,4);
TASK_PP(16'h13E90,4);
TASK_PP(16'h13E91,4);
TASK_PP(16'h13E92,4);
TASK_PP(16'h13E93,4);
TASK_PP(16'h13E94,4);
TASK_PP(16'h13E95,4);
TASK_PP(16'h13E96,4);
TASK_PP(16'h13E97,4);
TASK_PP(16'h13E98,4);
TASK_PP(16'h13E99,4);
TASK_PP(16'h13E9A,4);
TASK_PP(16'h13E9B,4);
TASK_PP(16'h13E9C,4);
TASK_PP(16'h13E9D,4);
TASK_PP(16'h13E9E,4);
TASK_PP(16'h13E9F,4);
TASK_PP(16'h13EA0,4);
TASK_PP(16'h13EA1,4);
TASK_PP(16'h13EA2,4);
TASK_PP(16'h13EA3,4);
TASK_PP(16'h13EA4,4);
TASK_PP(16'h13EA5,4);
TASK_PP(16'h13EA6,4);
TASK_PP(16'h13EA7,4);
TASK_PP(16'h13EA8,4);
TASK_PP(16'h13EA9,4);
TASK_PP(16'h13EAA,4);
TASK_PP(16'h13EAB,4);
TASK_PP(16'h13EAC,4);
TASK_PP(16'h13EAD,4);
TASK_PP(16'h13EAE,4);
TASK_PP(16'h13EAF,4);
TASK_PP(16'h13EB0,4);
TASK_PP(16'h13EB1,4);
TASK_PP(16'h13EB2,4);
TASK_PP(16'h13EB3,4);
TASK_PP(16'h13EB4,4);
TASK_PP(16'h13EB5,4);
TASK_PP(16'h13EB6,4);
TASK_PP(16'h13EB7,4);
TASK_PP(16'h13EB8,4);
TASK_PP(16'h13EB9,4);
TASK_PP(16'h13EBA,4);
TASK_PP(16'h13EBB,4);
TASK_PP(16'h13EBC,4);
TASK_PP(16'h13EBD,4);
TASK_PP(16'h13EBE,4);
TASK_PP(16'h13EBF,4);
TASK_PP(16'h13EC0,4);
TASK_PP(16'h13EC1,4);
TASK_PP(16'h13EC2,4);
TASK_PP(16'h13EC3,4);
TASK_PP(16'h13EC4,4);
TASK_PP(16'h13EC5,4);
TASK_PP(16'h13EC6,4);
TASK_PP(16'h13EC7,4);
TASK_PP(16'h13EC8,4);
TASK_PP(16'h13EC9,4);
TASK_PP(16'h13ECA,4);
TASK_PP(16'h13ECB,4);
TASK_PP(16'h13ECC,4);
TASK_PP(16'h13ECD,4);
TASK_PP(16'h13ECE,4);
TASK_PP(16'h13ECF,4);
TASK_PP(16'h13ED0,4);
TASK_PP(16'h13ED1,4);
TASK_PP(16'h13ED2,4);
TASK_PP(16'h13ED3,4);
TASK_PP(16'h13ED4,4);
TASK_PP(16'h13ED5,4);
TASK_PP(16'h13ED6,4);
TASK_PP(16'h13ED7,4);
TASK_PP(16'h13ED8,4);
TASK_PP(16'h13ED9,4);
TASK_PP(16'h13EDA,4);
TASK_PP(16'h13EDB,4);
TASK_PP(16'h13EDC,4);
TASK_PP(16'h13EDD,4);
TASK_PP(16'h13EDE,4);
TASK_PP(16'h13EDF,4);
TASK_PP(16'h13EE0,4);
TASK_PP(16'h13EE1,4);
TASK_PP(16'h13EE2,4);
TASK_PP(16'h13EE3,4);
TASK_PP(16'h13EE4,4);
TASK_PP(16'h13EE5,4);
TASK_PP(16'h13EE6,4);
TASK_PP(16'h13EE7,4);
TASK_PP(16'h13EE8,4);
TASK_PP(16'h13EE9,4);
TASK_PP(16'h13EEA,4);
TASK_PP(16'h13EEB,4);
TASK_PP(16'h13EEC,4);
TASK_PP(16'h13EED,4);
TASK_PP(16'h13EEE,4);
TASK_PP(16'h13EEF,4);
TASK_PP(16'h13EF0,4);
TASK_PP(16'h13EF1,4);
TASK_PP(16'h13EF2,4);
TASK_PP(16'h13EF3,4);
TASK_PP(16'h13EF4,4);
TASK_PP(16'h13EF5,4);
TASK_PP(16'h13EF6,4);
TASK_PP(16'h13EF7,4);
TASK_PP(16'h13EF8,4);
TASK_PP(16'h13EF9,4);
TASK_PP(16'h13EFA,4);
TASK_PP(16'h13EFB,4);
TASK_PP(16'h13EFC,4);
TASK_PP(16'h13EFD,4);
TASK_PP(16'h13EFE,4);
TASK_PP(16'h13EFF,4);
TASK_PP(16'h13F00,4);
TASK_PP(16'h13F01,4);
TASK_PP(16'h13F02,4);
TASK_PP(16'h13F03,4);
TASK_PP(16'h13F04,4);
TASK_PP(16'h13F05,4);
TASK_PP(16'h13F06,4);
TASK_PP(16'h13F07,4);
TASK_PP(16'h13F08,4);
TASK_PP(16'h13F09,4);
TASK_PP(16'h13F0A,4);
TASK_PP(16'h13F0B,4);
TASK_PP(16'h13F0C,4);
TASK_PP(16'h13F0D,4);
TASK_PP(16'h13F0E,4);
TASK_PP(16'h13F0F,4);
TASK_PP(16'h13F10,4);
TASK_PP(16'h13F11,4);
TASK_PP(16'h13F12,4);
TASK_PP(16'h13F13,4);
TASK_PP(16'h13F14,4);
TASK_PP(16'h13F15,4);
TASK_PP(16'h13F16,4);
TASK_PP(16'h13F17,4);
TASK_PP(16'h13F18,4);
TASK_PP(16'h13F19,4);
TASK_PP(16'h13F1A,4);
TASK_PP(16'h13F1B,4);
TASK_PP(16'h13F1C,4);
TASK_PP(16'h13F1D,4);
TASK_PP(16'h13F1E,4);
TASK_PP(16'h13F1F,4);
TASK_PP(16'h13F20,4);
TASK_PP(16'h13F21,4);
TASK_PP(16'h13F22,4);
TASK_PP(16'h13F23,4);
TASK_PP(16'h13F24,4);
TASK_PP(16'h13F25,4);
TASK_PP(16'h13F26,4);
TASK_PP(16'h13F27,4);
TASK_PP(16'h13F28,4);
TASK_PP(16'h13F29,4);
TASK_PP(16'h13F2A,4);
TASK_PP(16'h13F2B,4);
TASK_PP(16'h13F2C,4);
TASK_PP(16'h13F2D,4);
TASK_PP(16'h13F2E,4);
TASK_PP(16'h13F2F,4);
TASK_PP(16'h13F30,4);
TASK_PP(16'h13F31,4);
TASK_PP(16'h13F32,4);
TASK_PP(16'h13F33,4);
TASK_PP(16'h13F34,4);
TASK_PP(16'h13F35,4);
TASK_PP(16'h13F36,4);
TASK_PP(16'h13F37,4);
TASK_PP(16'h13F38,4);
TASK_PP(16'h13F39,4);
TASK_PP(16'h13F3A,4);
TASK_PP(16'h13F3B,4);
TASK_PP(16'h13F3C,4);
TASK_PP(16'h13F3D,4);
TASK_PP(16'h13F3E,4);
TASK_PP(16'h13F3F,4);
TASK_PP(16'h13F40,4);
TASK_PP(16'h13F41,4);
TASK_PP(16'h13F42,4);
TASK_PP(16'h13F43,4);
TASK_PP(16'h13F44,4);
TASK_PP(16'h13F45,4);
TASK_PP(16'h13F46,4);
TASK_PP(16'h13F47,4);
TASK_PP(16'h13F48,4);
TASK_PP(16'h13F49,4);
TASK_PP(16'h13F4A,4);
TASK_PP(16'h13F4B,4);
TASK_PP(16'h13F4C,4);
TASK_PP(16'h13F4D,4);
TASK_PP(16'h13F4E,4);
TASK_PP(16'h13F4F,4);
TASK_PP(16'h13F50,4);
TASK_PP(16'h13F51,4);
TASK_PP(16'h13F52,4);
TASK_PP(16'h13F53,4);
TASK_PP(16'h13F54,4);
TASK_PP(16'h13F55,4);
TASK_PP(16'h13F56,4);
TASK_PP(16'h13F57,4);
TASK_PP(16'h13F58,4);
TASK_PP(16'h13F59,4);
TASK_PP(16'h13F5A,4);
TASK_PP(16'h13F5B,4);
TASK_PP(16'h13F5C,4);
TASK_PP(16'h13F5D,4);
TASK_PP(16'h13F5E,4);
TASK_PP(16'h13F5F,4);
TASK_PP(16'h13F60,4);
TASK_PP(16'h13F61,4);
TASK_PP(16'h13F62,4);
TASK_PP(16'h13F63,4);
TASK_PP(16'h13F64,4);
TASK_PP(16'h13F65,4);
TASK_PP(16'h13F66,4);
TASK_PP(16'h13F67,4);
TASK_PP(16'h13F68,4);
TASK_PP(16'h13F69,4);
TASK_PP(16'h13F6A,4);
TASK_PP(16'h13F6B,4);
TASK_PP(16'h13F6C,4);
TASK_PP(16'h13F6D,4);
TASK_PP(16'h13F6E,4);
TASK_PP(16'h13F6F,4);
TASK_PP(16'h13F70,4);
TASK_PP(16'h13F71,4);
TASK_PP(16'h13F72,4);
TASK_PP(16'h13F73,4);
TASK_PP(16'h13F74,4);
TASK_PP(16'h13F75,4);
TASK_PP(16'h13F76,4);
TASK_PP(16'h13F77,4);
TASK_PP(16'h13F78,4);
TASK_PP(16'h13F79,4);
TASK_PP(16'h13F7A,4);
TASK_PP(16'h13F7B,4);
TASK_PP(16'h13F7C,4);
TASK_PP(16'h13F7D,4);
TASK_PP(16'h13F7E,4);
TASK_PP(16'h13F7F,4);
TASK_PP(16'h13F80,4);
TASK_PP(16'h13F81,4);
TASK_PP(16'h13F82,4);
TASK_PP(16'h13F83,4);
TASK_PP(16'h13F84,4);
TASK_PP(16'h13F85,4);
TASK_PP(16'h13F86,4);
TASK_PP(16'h13F87,4);
TASK_PP(16'h13F88,4);
TASK_PP(16'h13F89,4);
TASK_PP(16'h13F8A,4);
TASK_PP(16'h13F8B,4);
TASK_PP(16'h13F8C,4);
TASK_PP(16'h13F8D,4);
TASK_PP(16'h13F8E,4);
TASK_PP(16'h13F8F,4);
TASK_PP(16'h13F90,4);
TASK_PP(16'h13F91,4);
TASK_PP(16'h13F92,4);
TASK_PP(16'h13F93,4);
TASK_PP(16'h13F94,4);
TASK_PP(16'h13F95,4);
TASK_PP(16'h13F96,4);
TASK_PP(16'h13F97,4);
TASK_PP(16'h13F98,4);
TASK_PP(16'h13F99,4);
TASK_PP(16'h13F9A,4);
TASK_PP(16'h13F9B,4);
TASK_PP(16'h13F9C,4);
TASK_PP(16'h13F9D,4);
TASK_PP(16'h13F9E,4);
TASK_PP(16'h13F9F,4);
TASK_PP(16'h13FA0,4);
TASK_PP(16'h13FA1,4);
TASK_PP(16'h13FA2,4);
TASK_PP(16'h13FA3,4);
TASK_PP(16'h13FA4,4);
TASK_PP(16'h13FA5,4);
TASK_PP(16'h13FA6,4);
TASK_PP(16'h13FA7,4);
TASK_PP(16'h13FA8,4);
TASK_PP(16'h13FA9,4);
TASK_PP(16'h13FAA,4);
TASK_PP(16'h13FAB,4);
TASK_PP(16'h13FAC,4);
TASK_PP(16'h13FAD,4);
TASK_PP(16'h13FAE,4);
TASK_PP(16'h13FAF,4);
TASK_PP(16'h13FB0,4);
TASK_PP(16'h13FB1,4);
TASK_PP(16'h13FB2,4);
TASK_PP(16'h13FB3,4);
TASK_PP(16'h13FB4,4);
TASK_PP(16'h13FB5,4);
TASK_PP(16'h13FB6,4);
TASK_PP(16'h13FB7,4);
TASK_PP(16'h13FB8,4);
TASK_PP(16'h13FB9,4);
TASK_PP(16'h13FBA,4);
TASK_PP(16'h13FBB,4);
TASK_PP(16'h13FBC,4);
TASK_PP(16'h13FBD,4);
TASK_PP(16'h13FBE,4);
TASK_PP(16'h13FBF,4);
TASK_PP(16'h13FC0,4);
TASK_PP(16'h13FC1,4);
TASK_PP(16'h13FC2,4);
TASK_PP(16'h13FC3,4);
TASK_PP(16'h13FC4,4);
TASK_PP(16'h13FC5,4);
TASK_PP(16'h13FC6,4);
TASK_PP(16'h13FC7,4);
TASK_PP(16'h13FC8,4);
TASK_PP(16'h13FC9,4);
TASK_PP(16'h13FCA,4);
TASK_PP(16'h13FCB,4);
TASK_PP(16'h13FCC,4);
TASK_PP(16'h13FCD,4);
TASK_PP(16'h13FCE,4);
TASK_PP(16'h13FCF,4);
TASK_PP(16'h13FD0,4);
TASK_PP(16'h13FD1,4);
TASK_PP(16'h13FD2,4);
TASK_PP(16'h13FD3,4);
TASK_PP(16'h13FD4,4);
TASK_PP(16'h13FD5,4);
TASK_PP(16'h13FD6,4);
TASK_PP(16'h13FD7,4);
TASK_PP(16'h13FD8,4);
TASK_PP(16'h13FD9,4);
TASK_PP(16'h13FDA,4);
TASK_PP(16'h13FDB,4);
TASK_PP(16'h13FDC,4);
TASK_PP(16'h13FDD,4);
TASK_PP(16'h13FDE,4);
TASK_PP(16'h13FDF,4);
TASK_PP(16'h13FE0,4);
TASK_PP(16'h13FE1,4);
TASK_PP(16'h13FE2,4);
TASK_PP(16'h13FE3,4);
TASK_PP(16'h13FE4,4);
TASK_PP(16'h13FE5,4);
TASK_PP(16'h13FE6,4);
TASK_PP(16'h13FE7,4);
TASK_PP(16'h13FE8,4);
TASK_PP(16'h13FE9,4);
TASK_PP(16'h13FEA,4);
TASK_PP(16'h13FEB,4);
TASK_PP(16'h13FEC,4);
TASK_PP(16'h13FED,4);
TASK_PP(16'h13FEE,4);
TASK_PP(16'h13FEF,4);
TASK_PP(16'h13FF0,4);
TASK_PP(16'h13FF1,4);
TASK_PP(16'h13FF2,4);
TASK_PP(16'h13FF3,4);
TASK_PP(16'h13FF4,4);
TASK_PP(16'h13FF5,4);
TASK_PP(16'h13FF6,4);
TASK_PP(16'h13FF7,4);
TASK_PP(16'h13FF8,4);
TASK_PP(16'h13FF9,4);
TASK_PP(16'h13FFA,4);
TASK_PP(16'h13FFB,4);
TASK_PP(16'h13FFC,4);
TASK_PP(16'h13FFD,4);
TASK_PP(16'h13FFE,4);
TASK_PP(16'h13FFF,4);
TASK_PP(16'h14000,4);
TASK_PP(16'h14001,4);
TASK_PP(16'h14002,4);
TASK_PP(16'h14003,4);
TASK_PP(16'h14004,4);
TASK_PP(16'h14005,4);
TASK_PP(16'h14006,4);
TASK_PP(16'h14007,4);
TASK_PP(16'h14008,4);
TASK_PP(16'h14009,4);
TASK_PP(16'h1400A,4);
TASK_PP(16'h1400B,4);
TASK_PP(16'h1400C,4);
TASK_PP(16'h1400D,4);
TASK_PP(16'h1400E,4);
TASK_PP(16'h1400F,4);
TASK_PP(16'h14010,4);
TASK_PP(16'h14011,4);
TASK_PP(16'h14012,4);
TASK_PP(16'h14013,4);
TASK_PP(16'h14014,4);
TASK_PP(16'h14015,4);
TASK_PP(16'h14016,4);
TASK_PP(16'h14017,4);
TASK_PP(16'h14018,4);
TASK_PP(16'h14019,4);
TASK_PP(16'h1401A,4);
TASK_PP(16'h1401B,4);
TASK_PP(16'h1401C,4);
TASK_PP(16'h1401D,4);
TASK_PP(16'h1401E,4);
TASK_PP(16'h1401F,4);
TASK_PP(16'h14020,4);
TASK_PP(16'h14021,4);
TASK_PP(16'h14022,4);
TASK_PP(16'h14023,4);
TASK_PP(16'h14024,4);
TASK_PP(16'h14025,4);
TASK_PP(16'h14026,4);
TASK_PP(16'h14027,4);
TASK_PP(16'h14028,4);
TASK_PP(16'h14029,4);
TASK_PP(16'h1402A,4);
TASK_PP(16'h1402B,4);
TASK_PP(16'h1402C,4);
TASK_PP(16'h1402D,4);
TASK_PP(16'h1402E,4);
TASK_PP(16'h1402F,4);
TASK_PP(16'h14030,4);
TASK_PP(16'h14031,4);
TASK_PP(16'h14032,4);
TASK_PP(16'h14033,4);
TASK_PP(16'h14034,4);
TASK_PP(16'h14035,4);
TASK_PP(16'h14036,4);
TASK_PP(16'h14037,4);
TASK_PP(16'h14038,4);
TASK_PP(16'h14039,4);
TASK_PP(16'h1403A,4);
TASK_PP(16'h1403B,4);
TASK_PP(16'h1403C,4);
TASK_PP(16'h1403D,4);
TASK_PP(16'h1403E,4);
TASK_PP(16'h1403F,4);
TASK_PP(16'h14040,4);
TASK_PP(16'h14041,4);
TASK_PP(16'h14042,4);
TASK_PP(16'h14043,4);
TASK_PP(16'h14044,4);
TASK_PP(16'h14045,4);
TASK_PP(16'h14046,4);
TASK_PP(16'h14047,4);
TASK_PP(16'h14048,4);
TASK_PP(16'h14049,4);
TASK_PP(16'h1404A,4);
TASK_PP(16'h1404B,4);
TASK_PP(16'h1404C,4);
TASK_PP(16'h1404D,4);
TASK_PP(16'h1404E,4);
TASK_PP(16'h1404F,4);
TASK_PP(16'h14050,4);
TASK_PP(16'h14051,4);
TASK_PP(16'h14052,4);
TASK_PP(16'h14053,4);
TASK_PP(16'h14054,4);
TASK_PP(16'h14055,4);
TASK_PP(16'h14056,4);
TASK_PP(16'h14057,4);
TASK_PP(16'h14058,4);
TASK_PP(16'h14059,4);
TASK_PP(16'h1405A,4);
TASK_PP(16'h1405B,4);
TASK_PP(16'h1405C,4);
TASK_PP(16'h1405D,4);
TASK_PP(16'h1405E,4);
TASK_PP(16'h1405F,4);
TASK_PP(16'h14060,4);
TASK_PP(16'h14061,4);
TASK_PP(16'h14062,4);
TASK_PP(16'h14063,4);
TASK_PP(16'h14064,4);
TASK_PP(16'h14065,4);
TASK_PP(16'h14066,4);
TASK_PP(16'h14067,4);
TASK_PP(16'h14068,4);
TASK_PP(16'h14069,4);
TASK_PP(16'h1406A,4);
TASK_PP(16'h1406B,4);
TASK_PP(16'h1406C,4);
TASK_PP(16'h1406D,4);
TASK_PP(16'h1406E,4);
TASK_PP(16'h1406F,4);
TASK_PP(16'h14070,4);
TASK_PP(16'h14071,4);
TASK_PP(16'h14072,4);
TASK_PP(16'h14073,4);
TASK_PP(16'h14074,4);
TASK_PP(16'h14075,4);
TASK_PP(16'h14076,4);
TASK_PP(16'h14077,4);
TASK_PP(16'h14078,4);
TASK_PP(16'h14079,4);
TASK_PP(16'h1407A,4);
TASK_PP(16'h1407B,4);
TASK_PP(16'h1407C,4);
TASK_PP(16'h1407D,4);
TASK_PP(16'h1407E,4);
TASK_PP(16'h1407F,4);
TASK_PP(16'h14080,4);
TASK_PP(16'h14081,4);
TASK_PP(16'h14082,4);
TASK_PP(16'h14083,4);
TASK_PP(16'h14084,4);
TASK_PP(16'h14085,4);
TASK_PP(16'h14086,4);
TASK_PP(16'h14087,4);
TASK_PP(16'h14088,4);
TASK_PP(16'h14089,4);
TASK_PP(16'h1408A,4);
TASK_PP(16'h1408B,4);
TASK_PP(16'h1408C,4);
TASK_PP(16'h1408D,4);
TASK_PP(16'h1408E,4);
TASK_PP(16'h1408F,4);
TASK_PP(16'h14090,4);
TASK_PP(16'h14091,4);
TASK_PP(16'h14092,4);
TASK_PP(16'h14093,4);
TASK_PP(16'h14094,4);
TASK_PP(16'h14095,4);
TASK_PP(16'h14096,4);
TASK_PP(16'h14097,4);
TASK_PP(16'h14098,4);
TASK_PP(16'h14099,4);
TASK_PP(16'h1409A,4);
TASK_PP(16'h1409B,4);
TASK_PP(16'h1409C,4);
TASK_PP(16'h1409D,4);
TASK_PP(16'h1409E,4);
TASK_PP(16'h1409F,4);
TASK_PP(16'h140A0,4);
TASK_PP(16'h140A1,4);
TASK_PP(16'h140A2,4);
TASK_PP(16'h140A3,4);
TASK_PP(16'h140A4,4);
TASK_PP(16'h140A5,4);
TASK_PP(16'h140A6,4);
TASK_PP(16'h140A7,4);
TASK_PP(16'h140A8,4);
TASK_PP(16'h140A9,4);
TASK_PP(16'h140AA,4);
TASK_PP(16'h140AB,4);
TASK_PP(16'h140AC,4);
TASK_PP(16'h140AD,4);
TASK_PP(16'h140AE,4);
TASK_PP(16'h140AF,4);
TASK_PP(16'h140B0,4);
TASK_PP(16'h140B1,4);
TASK_PP(16'h140B2,4);
TASK_PP(16'h140B3,4);
TASK_PP(16'h140B4,4);
TASK_PP(16'h140B5,4);
TASK_PP(16'h140B6,4);
TASK_PP(16'h140B7,4);
TASK_PP(16'h140B8,4);
TASK_PP(16'h140B9,4);
TASK_PP(16'h140BA,4);
TASK_PP(16'h140BB,4);
TASK_PP(16'h140BC,4);
TASK_PP(16'h140BD,4);
TASK_PP(16'h140BE,4);
TASK_PP(16'h140BF,4);
TASK_PP(16'h140C0,4);
TASK_PP(16'h140C1,4);
TASK_PP(16'h140C2,4);
TASK_PP(16'h140C3,4);
TASK_PP(16'h140C4,4);
TASK_PP(16'h140C5,4);
TASK_PP(16'h140C6,4);
TASK_PP(16'h140C7,4);
TASK_PP(16'h140C8,4);
TASK_PP(16'h140C9,4);
TASK_PP(16'h140CA,4);
TASK_PP(16'h140CB,4);
TASK_PP(16'h140CC,4);
TASK_PP(16'h140CD,4);
TASK_PP(16'h140CE,4);
TASK_PP(16'h140CF,4);
TASK_PP(16'h140D0,4);
TASK_PP(16'h140D1,4);
TASK_PP(16'h140D2,4);
TASK_PP(16'h140D3,4);
TASK_PP(16'h140D4,4);
TASK_PP(16'h140D5,4);
TASK_PP(16'h140D6,4);
TASK_PP(16'h140D7,4);
TASK_PP(16'h140D8,4);
TASK_PP(16'h140D9,4);
TASK_PP(16'h140DA,4);
TASK_PP(16'h140DB,4);
TASK_PP(16'h140DC,4);
TASK_PP(16'h140DD,4);
TASK_PP(16'h140DE,4);
TASK_PP(16'h140DF,4);
TASK_PP(16'h140E0,4);
TASK_PP(16'h140E1,4);
TASK_PP(16'h140E2,4);
TASK_PP(16'h140E3,4);
TASK_PP(16'h140E4,4);
TASK_PP(16'h140E5,4);
TASK_PP(16'h140E6,4);
TASK_PP(16'h140E7,4);
TASK_PP(16'h140E8,4);
TASK_PP(16'h140E9,4);
TASK_PP(16'h140EA,4);
TASK_PP(16'h140EB,4);
TASK_PP(16'h140EC,4);
TASK_PP(16'h140ED,4);
TASK_PP(16'h140EE,4);
TASK_PP(16'h140EF,4);
TASK_PP(16'h140F0,4);
TASK_PP(16'h140F1,4);
TASK_PP(16'h140F2,4);
TASK_PP(16'h140F3,4);
TASK_PP(16'h140F4,4);
TASK_PP(16'h140F5,4);
TASK_PP(16'h140F6,4);
TASK_PP(16'h140F7,4);
TASK_PP(16'h140F8,4);
TASK_PP(16'h140F9,4);
TASK_PP(16'h140FA,4);
TASK_PP(16'h140FB,4);
TASK_PP(16'h140FC,4);
TASK_PP(16'h140FD,4);
TASK_PP(16'h140FE,4);
TASK_PP(16'h140FF,4);
TASK_PP(16'h14100,4);
TASK_PP(16'h14101,4);
TASK_PP(16'h14102,4);
TASK_PP(16'h14103,4);
TASK_PP(16'h14104,4);
TASK_PP(16'h14105,4);
TASK_PP(16'h14106,4);
TASK_PP(16'h14107,4);
TASK_PP(16'h14108,4);
TASK_PP(16'h14109,4);
TASK_PP(16'h1410A,4);
TASK_PP(16'h1410B,4);
TASK_PP(16'h1410C,4);
TASK_PP(16'h1410D,4);
TASK_PP(16'h1410E,4);
TASK_PP(16'h1410F,4);
TASK_PP(16'h14110,4);
TASK_PP(16'h14111,4);
TASK_PP(16'h14112,4);
TASK_PP(16'h14113,4);
TASK_PP(16'h14114,4);
TASK_PP(16'h14115,4);
TASK_PP(16'h14116,4);
TASK_PP(16'h14117,4);
TASK_PP(16'h14118,4);
TASK_PP(16'h14119,4);
TASK_PP(16'h1411A,4);
TASK_PP(16'h1411B,4);
TASK_PP(16'h1411C,4);
TASK_PP(16'h1411D,4);
TASK_PP(16'h1411E,4);
TASK_PP(16'h1411F,4);
TASK_PP(16'h14120,4);
TASK_PP(16'h14121,4);
TASK_PP(16'h14122,4);
TASK_PP(16'h14123,4);
TASK_PP(16'h14124,4);
TASK_PP(16'h14125,4);
TASK_PP(16'h14126,4);
TASK_PP(16'h14127,4);
TASK_PP(16'h14128,4);
TASK_PP(16'h14129,4);
TASK_PP(16'h1412A,4);
TASK_PP(16'h1412B,4);
TASK_PP(16'h1412C,4);
TASK_PP(16'h1412D,4);
TASK_PP(16'h1412E,4);
TASK_PP(16'h1412F,4);
TASK_PP(16'h14130,4);
TASK_PP(16'h14131,4);
TASK_PP(16'h14132,4);
TASK_PP(16'h14133,4);
TASK_PP(16'h14134,4);
TASK_PP(16'h14135,4);
TASK_PP(16'h14136,4);
TASK_PP(16'h14137,4);
TASK_PP(16'h14138,4);
TASK_PP(16'h14139,4);
TASK_PP(16'h1413A,4);
TASK_PP(16'h1413B,4);
TASK_PP(16'h1413C,4);
TASK_PP(16'h1413D,4);
TASK_PP(16'h1413E,4);
TASK_PP(16'h1413F,4);
TASK_PP(16'h14140,4);
TASK_PP(16'h14141,4);
TASK_PP(16'h14142,4);
TASK_PP(16'h14143,4);
TASK_PP(16'h14144,4);
TASK_PP(16'h14145,4);
TASK_PP(16'h14146,4);
TASK_PP(16'h14147,4);
TASK_PP(16'h14148,4);
TASK_PP(16'h14149,4);
TASK_PP(16'h1414A,4);
TASK_PP(16'h1414B,4);
TASK_PP(16'h1414C,4);
TASK_PP(16'h1414D,4);
TASK_PP(16'h1414E,4);
TASK_PP(16'h1414F,4);
TASK_PP(16'h14150,4);
TASK_PP(16'h14151,4);
TASK_PP(16'h14152,4);
TASK_PP(16'h14153,4);
TASK_PP(16'h14154,4);
TASK_PP(16'h14155,4);
TASK_PP(16'h14156,4);
TASK_PP(16'h14157,4);
TASK_PP(16'h14158,4);
TASK_PP(16'h14159,4);
TASK_PP(16'h1415A,4);
TASK_PP(16'h1415B,4);
TASK_PP(16'h1415C,4);
TASK_PP(16'h1415D,4);
TASK_PP(16'h1415E,4);
TASK_PP(16'h1415F,4);
TASK_PP(16'h14160,4);
TASK_PP(16'h14161,4);
TASK_PP(16'h14162,4);
TASK_PP(16'h14163,4);
TASK_PP(16'h14164,4);
TASK_PP(16'h14165,4);
TASK_PP(16'h14166,4);
TASK_PP(16'h14167,4);
TASK_PP(16'h14168,4);
TASK_PP(16'h14169,4);
TASK_PP(16'h1416A,4);
TASK_PP(16'h1416B,4);
TASK_PP(16'h1416C,4);
TASK_PP(16'h1416D,4);
TASK_PP(16'h1416E,4);
TASK_PP(16'h1416F,4);
TASK_PP(16'h14170,4);
TASK_PP(16'h14171,4);
TASK_PP(16'h14172,4);
TASK_PP(16'h14173,4);
TASK_PP(16'h14174,4);
TASK_PP(16'h14175,4);
TASK_PP(16'h14176,4);
TASK_PP(16'h14177,4);
TASK_PP(16'h14178,4);
TASK_PP(16'h14179,4);
TASK_PP(16'h1417A,4);
TASK_PP(16'h1417B,4);
TASK_PP(16'h1417C,4);
TASK_PP(16'h1417D,4);
TASK_PP(16'h1417E,4);
TASK_PP(16'h1417F,4);
TASK_PP(16'h14180,4);
TASK_PP(16'h14181,4);
TASK_PP(16'h14182,4);
TASK_PP(16'h14183,4);
TASK_PP(16'h14184,4);
TASK_PP(16'h14185,4);
TASK_PP(16'h14186,4);
TASK_PP(16'h14187,4);
TASK_PP(16'h14188,4);
TASK_PP(16'h14189,4);
TASK_PP(16'h1418A,4);
TASK_PP(16'h1418B,4);
TASK_PP(16'h1418C,4);
TASK_PP(16'h1418D,4);
TASK_PP(16'h1418E,4);
TASK_PP(16'h1418F,4);
TASK_PP(16'h14190,4);
TASK_PP(16'h14191,4);
TASK_PP(16'h14192,4);
TASK_PP(16'h14193,4);
TASK_PP(16'h14194,4);
TASK_PP(16'h14195,4);
TASK_PP(16'h14196,4);
TASK_PP(16'h14197,4);
TASK_PP(16'h14198,4);
TASK_PP(16'h14199,4);
TASK_PP(16'h1419A,4);
TASK_PP(16'h1419B,4);
TASK_PP(16'h1419C,4);
TASK_PP(16'h1419D,4);
TASK_PP(16'h1419E,4);
TASK_PP(16'h1419F,4);
TASK_PP(16'h141A0,4);
TASK_PP(16'h141A1,4);
TASK_PP(16'h141A2,4);
TASK_PP(16'h141A3,4);
TASK_PP(16'h141A4,4);
TASK_PP(16'h141A5,4);
TASK_PP(16'h141A6,4);
TASK_PP(16'h141A7,4);
TASK_PP(16'h141A8,4);
TASK_PP(16'h141A9,4);
TASK_PP(16'h141AA,4);
TASK_PP(16'h141AB,4);
TASK_PP(16'h141AC,4);
TASK_PP(16'h141AD,4);
TASK_PP(16'h141AE,4);
TASK_PP(16'h141AF,4);
TASK_PP(16'h141B0,4);
TASK_PP(16'h141B1,4);
TASK_PP(16'h141B2,4);
TASK_PP(16'h141B3,4);
TASK_PP(16'h141B4,4);
TASK_PP(16'h141B5,4);
TASK_PP(16'h141B6,4);
TASK_PP(16'h141B7,4);
TASK_PP(16'h141B8,4);
TASK_PP(16'h141B9,4);
TASK_PP(16'h141BA,4);
TASK_PP(16'h141BB,4);
TASK_PP(16'h141BC,4);
TASK_PP(16'h141BD,4);
TASK_PP(16'h141BE,4);
TASK_PP(16'h141BF,4);
TASK_PP(16'h141C0,4);
TASK_PP(16'h141C1,4);
TASK_PP(16'h141C2,4);
TASK_PP(16'h141C3,4);
TASK_PP(16'h141C4,4);
TASK_PP(16'h141C5,4);
TASK_PP(16'h141C6,4);
TASK_PP(16'h141C7,4);
TASK_PP(16'h141C8,4);
TASK_PP(16'h141C9,4);
TASK_PP(16'h141CA,4);
TASK_PP(16'h141CB,4);
TASK_PP(16'h141CC,4);
TASK_PP(16'h141CD,4);
TASK_PP(16'h141CE,4);
TASK_PP(16'h141CF,4);
TASK_PP(16'h141D0,4);
TASK_PP(16'h141D1,4);
TASK_PP(16'h141D2,4);
TASK_PP(16'h141D3,4);
TASK_PP(16'h141D4,4);
TASK_PP(16'h141D5,4);
TASK_PP(16'h141D6,4);
TASK_PP(16'h141D7,4);
TASK_PP(16'h141D8,4);
TASK_PP(16'h141D9,4);
TASK_PP(16'h141DA,4);
TASK_PP(16'h141DB,4);
TASK_PP(16'h141DC,4);
TASK_PP(16'h141DD,4);
TASK_PP(16'h141DE,4);
TASK_PP(16'h141DF,4);
TASK_PP(16'h141E0,4);
TASK_PP(16'h141E1,4);
TASK_PP(16'h141E2,4);
TASK_PP(16'h141E3,4);
TASK_PP(16'h141E4,4);
TASK_PP(16'h141E5,4);
TASK_PP(16'h141E6,4);
TASK_PP(16'h141E7,4);
TASK_PP(16'h141E8,4);
TASK_PP(16'h141E9,4);
TASK_PP(16'h141EA,4);
TASK_PP(16'h141EB,4);
TASK_PP(16'h141EC,4);
TASK_PP(16'h141ED,4);
TASK_PP(16'h141EE,4);
TASK_PP(16'h141EF,4);
TASK_PP(16'h141F0,4);
TASK_PP(16'h141F1,4);
TASK_PP(16'h141F2,4);
TASK_PP(16'h141F3,4);
TASK_PP(16'h141F4,4);
TASK_PP(16'h141F5,4);
TASK_PP(16'h141F6,4);
TASK_PP(16'h141F7,4);
TASK_PP(16'h141F8,4);
TASK_PP(16'h141F9,4);
TASK_PP(16'h141FA,4);
TASK_PP(16'h141FB,4);
TASK_PP(16'h141FC,4);
TASK_PP(16'h141FD,4);
TASK_PP(16'h141FE,4);
TASK_PP(16'h141FF,4);
TASK_PP(16'h14200,4);
TASK_PP(16'h14201,4);
TASK_PP(16'h14202,4);
TASK_PP(16'h14203,4);
TASK_PP(16'h14204,4);
TASK_PP(16'h14205,4);
TASK_PP(16'h14206,4);
TASK_PP(16'h14207,4);
TASK_PP(16'h14208,4);
TASK_PP(16'h14209,4);
TASK_PP(16'h1420A,4);
TASK_PP(16'h1420B,4);
TASK_PP(16'h1420C,4);
TASK_PP(16'h1420D,4);
TASK_PP(16'h1420E,4);
TASK_PP(16'h1420F,4);
TASK_PP(16'h14210,4);
TASK_PP(16'h14211,4);
TASK_PP(16'h14212,4);
TASK_PP(16'h14213,4);
TASK_PP(16'h14214,4);
TASK_PP(16'h14215,4);
TASK_PP(16'h14216,4);
TASK_PP(16'h14217,4);
TASK_PP(16'h14218,4);
TASK_PP(16'h14219,4);
TASK_PP(16'h1421A,4);
TASK_PP(16'h1421B,4);
TASK_PP(16'h1421C,4);
TASK_PP(16'h1421D,4);
TASK_PP(16'h1421E,4);
TASK_PP(16'h1421F,4);
TASK_PP(16'h14220,4);
TASK_PP(16'h14221,4);
TASK_PP(16'h14222,4);
TASK_PP(16'h14223,4);
TASK_PP(16'h14224,4);
TASK_PP(16'h14225,4);
TASK_PP(16'h14226,4);
TASK_PP(16'h14227,4);
TASK_PP(16'h14228,4);
TASK_PP(16'h14229,4);
TASK_PP(16'h1422A,4);
TASK_PP(16'h1422B,4);
TASK_PP(16'h1422C,4);
TASK_PP(16'h1422D,4);
TASK_PP(16'h1422E,4);
TASK_PP(16'h1422F,4);
TASK_PP(16'h14230,4);
TASK_PP(16'h14231,4);
TASK_PP(16'h14232,4);
TASK_PP(16'h14233,4);
TASK_PP(16'h14234,4);
TASK_PP(16'h14235,4);
TASK_PP(16'h14236,4);
TASK_PP(16'h14237,4);
TASK_PP(16'h14238,4);
TASK_PP(16'h14239,4);
TASK_PP(16'h1423A,4);
TASK_PP(16'h1423B,4);
TASK_PP(16'h1423C,4);
TASK_PP(16'h1423D,4);
TASK_PP(16'h1423E,4);
TASK_PP(16'h1423F,4);
TASK_PP(16'h14240,4);
TASK_PP(16'h14241,4);
TASK_PP(16'h14242,4);
TASK_PP(16'h14243,4);
TASK_PP(16'h14244,4);
TASK_PP(16'h14245,4);
TASK_PP(16'h14246,4);
TASK_PP(16'h14247,4);
TASK_PP(16'h14248,4);
TASK_PP(16'h14249,4);
TASK_PP(16'h1424A,4);
TASK_PP(16'h1424B,4);
TASK_PP(16'h1424C,4);
TASK_PP(16'h1424D,4);
TASK_PP(16'h1424E,4);
TASK_PP(16'h1424F,4);
TASK_PP(16'h14250,4);
TASK_PP(16'h14251,4);
TASK_PP(16'h14252,4);
TASK_PP(16'h14253,4);
TASK_PP(16'h14254,4);
TASK_PP(16'h14255,4);
TASK_PP(16'h14256,4);
TASK_PP(16'h14257,4);
TASK_PP(16'h14258,4);
TASK_PP(16'h14259,4);
TASK_PP(16'h1425A,4);
TASK_PP(16'h1425B,4);
TASK_PP(16'h1425C,4);
TASK_PP(16'h1425D,4);
TASK_PP(16'h1425E,4);
TASK_PP(16'h1425F,4);
TASK_PP(16'h14260,4);
TASK_PP(16'h14261,4);
TASK_PP(16'h14262,4);
TASK_PP(16'h14263,4);
TASK_PP(16'h14264,4);
TASK_PP(16'h14265,4);
TASK_PP(16'h14266,4);
TASK_PP(16'h14267,4);
TASK_PP(16'h14268,4);
TASK_PP(16'h14269,4);
TASK_PP(16'h1426A,4);
TASK_PP(16'h1426B,4);
TASK_PP(16'h1426C,4);
TASK_PP(16'h1426D,4);
TASK_PP(16'h1426E,4);
TASK_PP(16'h1426F,4);
TASK_PP(16'h14270,4);
TASK_PP(16'h14271,4);
TASK_PP(16'h14272,4);
TASK_PP(16'h14273,4);
TASK_PP(16'h14274,4);
TASK_PP(16'h14275,4);
TASK_PP(16'h14276,4);
TASK_PP(16'h14277,4);
TASK_PP(16'h14278,4);
TASK_PP(16'h14279,4);
TASK_PP(16'h1427A,4);
TASK_PP(16'h1427B,4);
TASK_PP(16'h1427C,4);
TASK_PP(16'h1427D,4);
TASK_PP(16'h1427E,4);
TASK_PP(16'h1427F,4);
TASK_PP(16'h14280,4);
TASK_PP(16'h14281,4);
TASK_PP(16'h14282,4);
TASK_PP(16'h14283,4);
TASK_PP(16'h14284,4);
TASK_PP(16'h14285,4);
TASK_PP(16'h14286,4);
TASK_PP(16'h14287,4);
TASK_PP(16'h14288,4);
TASK_PP(16'h14289,4);
TASK_PP(16'h1428A,4);
TASK_PP(16'h1428B,4);
TASK_PP(16'h1428C,4);
TASK_PP(16'h1428D,4);
TASK_PP(16'h1428E,4);
TASK_PP(16'h1428F,4);
TASK_PP(16'h14290,4);
TASK_PP(16'h14291,4);
TASK_PP(16'h14292,4);
TASK_PP(16'h14293,4);
TASK_PP(16'h14294,4);
TASK_PP(16'h14295,4);
TASK_PP(16'h14296,4);
TASK_PP(16'h14297,4);
TASK_PP(16'h14298,4);
TASK_PP(16'h14299,4);
TASK_PP(16'h1429A,4);
TASK_PP(16'h1429B,4);
TASK_PP(16'h1429C,4);
TASK_PP(16'h1429D,4);
TASK_PP(16'h1429E,4);
TASK_PP(16'h1429F,4);
TASK_PP(16'h142A0,4);
TASK_PP(16'h142A1,4);
TASK_PP(16'h142A2,4);
TASK_PP(16'h142A3,4);
TASK_PP(16'h142A4,4);
TASK_PP(16'h142A5,4);
TASK_PP(16'h142A6,4);
TASK_PP(16'h142A7,4);
TASK_PP(16'h142A8,4);
TASK_PP(16'h142A9,4);
TASK_PP(16'h142AA,4);
TASK_PP(16'h142AB,4);
TASK_PP(16'h142AC,4);
TASK_PP(16'h142AD,4);
TASK_PP(16'h142AE,4);
TASK_PP(16'h142AF,4);
TASK_PP(16'h142B0,4);
TASK_PP(16'h142B1,4);
TASK_PP(16'h142B2,4);
TASK_PP(16'h142B3,4);
TASK_PP(16'h142B4,4);
TASK_PP(16'h142B5,4);
TASK_PP(16'h142B6,4);
TASK_PP(16'h142B7,4);
TASK_PP(16'h142B8,4);
TASK_PP(16'h142B9,4);
TASK_PP(16'h142BA,4);
TASK_PP(16'h142BB,4);
TASK_PP(16'h142BC,4);
TASK_PP(16'h142BD,4);
TASK_PP(16'h142BE,4);
TASK_PP(16'h142BF,4);
TASK_PP(16'h142C0,4);
TASK_PP(16'h142C1,4);
TASK_PP(16'h142C2,4);
TASK_PP(16'h142C3,4);
TASK_PP(16'h142C4,4);
TASK_PP(16'h142C5,4);
TASK_PP(16'h142C6,4);
TASK_PP(16'h142C7,4);
TASK_PP(16'h142C8,4);
TASK_PP(16'h142C9,4);
TASK_PP(16'h142CA,4);
TASK_PP(16'h142CB,4);
TASK_PP(16'h142CC,4);
TASK_PP(16'h142CD,4);
TASK_PP(16'h142CE,4);
TASK_PP(16'h142CF,4);
TASK_PP(16'h142D0,4);
TASK_PP(16'h142D1,4);
TASK_PP(16'h142D2,4);
TASK_PP(16'h142D3,4);
TASK_PP(16'h142D4,4);
TASK_PP(16'h142D5,4);
TASK_PP(16'h142D6,4);
TASK_PP(16'h142D7,4);
TASK_PP(16'h142D8,4);
TASK_PP(16'h142D9,4);
TASK_PP(16'h142DA,4);
TASK_PP(16'h142DB,4);
TASK_PP(16'h142DC,4);
TASK_PP(16'h142DD,4);
TASK_PP(16'h142DE,4);
TASK_PP(16'h142DF,4);
TASK_PP(16'h142E0,4);
TASK_PP(16'h142E1,4);
TASK_PP(16'h142E2,4);
TASK_PP(16'h142E3,4);
TASK_PP(16'h142E4,4);
TASK_PP(16'h142E5,4);
TASK_PP(16'h142E6,4);
TASK_PP(16'h142E7,4);
TASK_PP(16'h142E8,4);
TASK_PP(16'h142E9,4);
TASK_PP(16'h142EA,4);
TASK_PP(16'h142EB,4);
TASK_PP(16'h142EC,4);
TASK_PP(16'h142ED,4);
TASK_PP(16'h142EE,4);
TASK_PP(16'h142EF,4);
TASK_PP(16'h142F0,4);
TASK_PP(16'h142F1,4);
TASK_PP(16'h142F2,4);
TASK_PP(16'h142F3,4);
TASK_PP(16'h142F4,4);
TASK_PP(16'h142F5,4);
TASK_PP(16'h142F6,4);
TASK_PP(16'h142F7,4);
TASK_PP(16'h142F8,4);
TASK_PP(16'h142F9,4);
TASK_PP(16'h142FA,4);
TASK_PP(16'h142FB,4);
TASK_PP(16'h142FC,4);
TASK_PP(16'h142FD,4);
TASK_PP(16'h142FE,4);
TASK_PP(16'h142FF,4);
TASK_PP(16'h14300,4);
TASK_PP(16'h14301,4);
TASK_PP(16'h14302,4);
TASK_PP(16'h14303,4);
TASK_PP(16'h14304,4);
TASK_PP(16'h14305,4);
TASK_PP(16'h14306,4);
TASK_PP(16'h14307,4);
TASK_PP(16'h14308,4);
TASK_PP(16'h14309,4);
TASK_PP(16'h1430A,4);
TASK_PP(16'h1430B,4);
TASK_PP(16'h1430C,4);
TASK_PP(16'h1430D,4);
TASK_PP(16'h1430E,4);
TASK_PP(16'h1430F,4);
TASK_PP(16'h14310,4);
TASK_PP(16'h14311,4);
TASK_PP(16'h14312,4);
TASK_PP(16'h14313,4);
TASK_PP(16'h14314,4);
TASK_PP(16'h14315,4);
TASK_PP(16'h14316,4);
TASK_PP(16'h14317,4);
TASK_PP(16'h14318,4);
TASK_PP(16'h14319,4);
TASK_PP(16'h1431A,4);
TASK_PP(16'h1431B,4);
TASK_PP(16'h1431C,4);
TASK_PP(16'h1431D,4);
TASK_PP(16'h1431E,4);
TASK_PP(16'h1431F,4);
TASK_PP(16'h14320,4);
TASK_PP(16'h14321,4);
TASK_PP(16'h14322,4);
TASK_PP(16'h14323,4);
TASK_PP(16'h14324,4);
TASK_PP(16'h14325,4);
TASK_PP(16'h14326,4);
TASK_PP(16'h14327,4);
TASK_PP(16'h14328,4);
TASK_PP(16'h14329,4);
TASK_PP(16'h1432A,4);
TASK_PP(16'h1432B,4);
TASK_PP(16'h1432C,4);
TASK_PP(16'h1432D,4);
TASK_PP(16'h1432E,4);
TASK_PP(16'h1432F,4);
TASK_PP(16'h14330,4);
TASK_PP(16'h14331,4);
TASK_PP(16'h14332,4);
TASK_PP(16'h14333,4);
TASK_PP(16'h14334,4);
TASK_PP(16'h14335,4);
TASK_PP(16'h14336,4);
TASK_PP(16'h14337,4);
TASK_PP(16'h14338,4);
TASK_PP(16'h14339,4);
TASK_PP(16'h1433A,4);
TASK_PP(16'h1433B,4);
TASK_PP(16'h1433C,4);
TASK_PP(16'h1433D,4);
TASK_PP(16'h1433E,4);
TASK_PP(16'h1433F,4);
TASK_PP(16'h14340,4);
TASK_PP(16'h14341,4);
TASK_PP(16'h14342,4);
TASK_PP(16'h14343,4);
TASK_PP(16'h14344,4);
TASK_PP(16'h14345,4);
TASK_PP(16'h14346,4);
TASK_PP(16'h14347,4);
TASK_PP(16'h14348,4);
TASK_PP(16'h14349,4);
TASK_PP(16'h1434A,4);
TASK_PP(16'h1434B,4);
TASK_PP(16'h1434C,4);
TASK_PP(16'h1434D,4);
TASK_PP(16'h1434E,4);
TASK_PP(16'h1434F,4);
TASK_PP(16'h14350,4);
TASK_PP(16'h14351,4);
TASK_PP(16'h14352,4);
TASK_PP(16'h14353,4);
TASK_PP(16'h14354,4);
TASK_PP(16'h14355,4);
TASK_PP(16'h14356,4);
TASK_PP(16'h14357,4);
TASK_PP(16'h14358,4);
TASK_PP(16'h14359,4);
TASK_PP(16'h1435A,4);
TASK_PP(16'h1435B,4);
TASK_PP(16'h1435C,4);
TASK_PP(16'h1435D,4);
TASK_PP(16'h1435E,4);
TASK_PP(16'h1435F,4);
TASK_PP(16'h14360,4);
TASK_PP(16'h14361,4);
TASK_PP(16'h14362,4);
TASK_PP(16'h14363,4);
TASK_PP(16'h14364,4);
TASK_PP(16'h14365,4);
TASK_PP(16'h14366,4);
TASK_PP(16'h14367,4);
TASK_PP(16'h14368,4);
TASK_PP(16'h14369,4);
TASK_PP(16'h1436A,4);
TASK_PP(16'h1436B,4);
TASK_PP(16'h1436C,4);
TASK_PP(16'h1436D,4);
TASK_PP(16'h1436E,4);
TASK_PP(16'h1436F,4);
TASK_PP(16'h14370,4);
TASK_PP(16'h14371,4);
TASK_PP(16'h14372,4);
TASK_PP(16'h14373,4);
TASK_PP(16'h14374,4);
TASK_PP(16'h14375,4);
TASK_PP(16'h14376,4);
TASK_PP(16'h14377,4);
TASK_PP(16'h14378,4);
TASK_PP(16'h14379,4);
TASK_PP(16'h1437A,4);
TASK_PP(16'h1437B,4);
TASK_PP(16'h1437C,4);
TASK_PP(16'h1437D,4);
TASK_PP(16'h1437E,4);
TASK_PP(16'h1437F,4);
TASK_PP(16'h14380,4);
TASK_PP(16'h14381,4);
TASK_PP(16'h14382,4);
TASK_PP(16'h14383,4);
TASK_PP(16'h14384,4);
TASK_PP(16'h14385,4);
TASK_PP(16'h14386,4);
TASK_PP(16'h14387,4);
TASK_PP(16'h14388,4);
TASK_PP(16'h14389,4);
TASK_PP(16'h1438A,4);
TASK_PP(16'h1438B,4);
TASK_PP(16'h1438C,4);
TASK_PP(16'h1438D,4);
TASK_PP(16'h1438E,4);
TASK_PP(16'h1438F,4);
TASK_PP(16'h14390,4);
TASK_PP(16'h14391,4);
TASK_PP(16'h14392,4);
TASK_PP(16'h14393,4);
TASK_PP(16'h14394,4);
TASK_PP(16'h14395,4);
TASK_PP(16'h14396,4);
TASK_PP(16'h14397,4);
TASK_PP(16'h14398,4);
TASK_PP(16'h14399,4);
TASK_PP(16'h1439A,4);
TASK_PP(16'h1439B,4);
TASK_PP(16'h1439C,4);
TASK_PP(16'h1439D,4);
TASK_PP(16'h1439E,4);
TASK_PP(16'h1439F,4);
TASK_PP(16'h143A0,4);
TASK_PP(16'h143A1,4);
TASK_PP(16'h143A2,4);
TASK_PP(16'h143A3,4);
TASK_PP(16'h143A4,4);
TASK_PP(16'h143A5,4);
TASK_PP(16'h143A6,4);
TASK_PP(16'h143A7,4);
TASK_PP(16'h143A8,4);
TASK_PP(16'h143A9,4);
TASK_PP(16'h143AA,4);
TASK_PP(16'h143AB,4);
TASK_PP(16'h143AC,4);
TASK_PP(16'h143AD,4);
TASK_PP(16'h143AE,4);
TASK_PP(16'h143AF,4);
TASK_PP(16'h143B0,4);
TASK_PP(16'h143B1,4);
TASK_PP(16'h143B2,4);
TASK_PP(16'h143B3,4);
TASK_PP(16'h143B4,4);
TASK_PP(16'h143B5,4);
TASK_PP(16'h143B6,4);
TASK_PP(16'h143B7,4);
TASK_PP(16'h143B8,4);
TASK_PP(16'h143B9,4);
TASK_PP(16'h143BA,4);
TASK_PP(16'h143BB,4);
TASK_PP(16'h143BC,4);
TASK_PP(16'h143BD,4);
TASK_PP(16'h143BE,4);
TASK_PP(16'h143BF,4);
TASK_PP(16'h143C0,4);
TASK_PP(16'h143C1,4);
TASK_PP(16'h143C2,4);
TASK_PP(16'h143C3,4);
TASK_PP(16'h143C4,4);
TASK_PP(16'h143C5,4);
TASK_PP(16'h143C6,4);
TASK_PP(16'h143C7,4);
TASK_PP(16'h143C8,4);
TASK_PP(16'h143C9,4);
TASK_PP(16'h143CA,4);
TASK_PP(16'h143CB,4);
TASK_PP(16'h143CC,4);
TASK_PP(16'h143CD,4);
TASK_PP(16'h143CE,4);
TASK_PP(16'h143CF,4);
TASK_PP(16'h143D0,4);
TASK_PP(16'h143D1,4);
TASK_PP(16'h143D2,4);
TASK_PP(16'h143D3,4);
TASK_PP(16'h143D4,4);
TASK_PP(16'h143D5,4);
TASK_PP(16'h143D6,4);
TASK_PP(16'h143D7,4);
TASK_PP(16'h143D8,4);
TASK_PP(16'h143D9,4);
TASK_PP(16'h143DA,4);
TASK_PP(16'h143DB,4);
TASK_PP(16'h143DC,4);
TASK_PP(16'h143DD,4);
TASK_PP(16'h143DE,4);
TASK_PP(16'h143DF,4);
TASK_PP(16'h143E0,4);
TASK_PP(16'h143E1,4);
TASK_PP(16'h143E2,4);
TASK_PP(16'h143E3,4);
TASK_PP(16'h143E4,4);
TASK_PP(16'h143E5,4);
TASK_PP(16'h143E6,4);
TASK_PP(16'h143E7,4);
TASK_PP(16'h143E8,4);
TASK_PP(16'h143E9,4);
TASK_PP(16'h143EA,4);
TASK_PP(16'h143EB,4);
TASK_PP(16'h143EC,4);
TASK_PP(16'h143ED,4);
TASK_PP(16'h143EE,4);
TASK_PP(16'h143EF,4);
TASK_PP(16'h143F0,4);
TASK_PP(16'h143F1,4);
TASK_PP(16'h143F2,4);
TASK_PP(16'h143F3,4);
TASK_PP(16'h143F4,4);
TASK_PP(16'h143F5,4);
TASK_PP(16'h143F6,4);
TASK_PP(16'h143F7,4);
TASK_PP(16'h143F8,4);
TASK_PP(16'h143F9,4);
TASK_PP(16'h143FA,4);
TASK_PP(16'h143FB,4);
TASK_PP(16'h143FC,4);
TASK_PP(16'h143FD,4);
TASK_PP(16'h143FE,4);
TASK_PP(16'h143FF,4);
TASK_PP(16'h14400,4);
TASK_PP(16'h14401,4);
TASK_PP(16'h14402,4);
TASK_PP(16'h14403,4);
TASK_PP(16'h14404,4);
TASK_PP(16'h14405,4);
TASK_PP(16'h14406,4);
TASK_PP(16'h14407,4);
TASK_PP(16'h14408,4);
TASK_PP(16'h14409,4);
TASK_PP(16'h1440A,4);
TASK_PP(16'h1440B,4);
TASK_PP(16'h1440C,4);
TASK_PP(16'h1440D,4);
TASK_PP(16'h1440E,4);
TASK_PP(16'h1440F,4);
TASK_PP(16'h14410,4);
TASK_PP(16'h14411,4);
TASK_PP(16'h14412,4);
TASK_PP(16'h14413,4);
TASK_PP(16'h14414,4);
TASK_PP(16'h14415,4);
TASK_PP(16'h14416,4);
TASK_PP(16'h14417,4);
TASK_PP(16'h14418,4);
TASK_PP(16'h14419,4);
TASK_PP(16'h1441A,4);
TASK_PP(16'h1441B,4);
TASK_PP(16'h1441C,4);
TASK_PP(16'h1441D,4);
TASK_PP(16'h1441E,4);
TASK_PP(16'h1441F,4);
TASK_PP(16'h14420,4);
TASK_PP(16'h14421,4);
TASK_PP(16'h14422,4);
TASK_PP(16'h14423,4);
TASK_PP(16'h14424,4);
TASK_PP(16'h14425,4);
TASK_PP(16'h14426,4);
TASK_PP(16'h14427,4);
TASK_PP(16'h14428,4);
TASK_PP(16'h14429,4);
TASK_PP(16'h1442A,4);
TASK_PP(16'h1442B,4);
TASK_PP(16'h1442C,4);
TASK_PP(16'h1442D,4);
TASK_PP(16'h1442E,4);
TASK_PP(16'h1442F,4);
TASK_PP(16'h14430,4);
TASK_PP(16'h14431,4);
TASK_PP(16'h14432,4);
TASK_PP(16'h14433,4);
TASK_PP(16'h14434,4);
TASK_PP(16'h14435,4);
TASK_PP(16'h14436,4);
TASK_PP(16'h14437,4);
TASK_PP(16'h14438,4);
TASK_PP(16'h14439,4);
TASK_PP(16'h1443A,4);
TASK_PP(16'h1443B,4);
TASK_PP(16'h1443C,4);
TASK_PP(16'h1443D,4);
TASK_PP(16'h1443E,4);
TASK_PP(16'h1443F,4);
TASK_PP(16'h14440,4);
TASK_PP(16'h14441,4);
TASK_PP(16'h14442,4);
TASK_PP(16'h14443,4);
TASK_PP(16'h14444,4);
TASK_PP(16'h14445,4);
TASK_PP(16'h14446,4);
TASK_PP(16'h14447,4);
TASK_PP(16'h14448,4);
TASK_PP(16'h14449,4);
TASK_PP(16'h1444A,4);
TASK_PP(16'h1444B,4);
TASK_PP(16'h1444C,4);
TASK_PP(16'h1444D,4);
TASK_PP(16'h1444E,4);
TASK_PP(16'h1444F,4);
TASK_PP(16'h14450,4);
TASK_PP(16'h14451,4);
TASK_PP(16'h14452,4);
TASK_PP(16'h14453,4);
TASK_PP(16'h14454,4);
TASK_PP(16'h14455,4);
TASK_PP(16'h14456,4);
TASK_PP(16'h14457,4);
TASK_PP(16'h14458,4);
TASK_PP(16'h14459,4);
TASK_PP(16'h1445A,4);
TASK_PP(16'h1445B,4);
TASK_PP(16'h1445C,4);
TASK_PP(16'h1445D,4);
TASK_PP(16'h1445E,4);
TASK_PP(16'h1445F,4);
TASK_PP(16'h14460,4);
TASK_PP(16'h14461,4);
TASK_PP(16'h14462,4);
TASK_PP(16'h14463,4);
TASK_PP(16'h14464,4);
TASK_PP(16'h14465,4);
TASK_PP(16'h14466,4);
TASK_PP(16'h14467,4);
TASK_PP(16'h14468,4);
TASK_PP(16'h14469,4);
TASK_PP(16'h1446A,4);
TASK_PP(16'h1446B,4);
TASK_PP(16'h1446C,4);
TASK_PP(16'h1446D,4);
TASK_PP(16'h1446E,4);
TASK_PP(16'h1446F,4);
TASK_PP(16'h14470,4);
TASK_PP(16'h14471,4);
TASK_PP(16'h14472,4);
TASK_PP(16'h14473,4);
TASK_PP(16'h14474,4);
TASK_PP(16'h14475,4);
TASK_PP(16'h14476,4);
TASK_PP(16'h14477,4);
TASK_PP(16'h14478,4);
TASK_PP(16'h14479,4);
TASK_PP(16'h1447A,4);
TASK_PP(16'h1447B,4);
TASK_PP(16'h1447C,4);
TASK_PP(16'h1447D,4);
TASK_PP(16'h1447E,4);
TASK_PP(16'h1447F,4);
TASK_PP(16'h14480,4);
TASK_PP(16'h14481,4);
TASK_PP(16'h14482,4);
TASK_PP(16'h14483,4);
TASK_PP(16'h14484,4);
TASK_PP(16'h14485,4);
TASK_PP(16'h14486,4);
TASK_PP(16'h14487,4);
TASK_PP(16'h14488,4);
TASK_PP(16'h14489,4);
TASK_PP(16'h1448A,4);
TASK_PP(16'h1448B,4);
TASK_PP(16'h1448C,4);
TASK_PP(16'h1448D,4);
TASK_PP(16'h1448E,4);
TASK_PP(16'h1448F,4);
TASK_PP(16'h14490,4);
TASK_PP(16'h14491,4);
TASK_PP(16'h14492,4);
TASK_PP(16'h14493,4);
TASK_PP(16'h14494,4);
TASK_PP(16'h14495,4);
TASK_PP(16'h14496,4);
TASK_PP(16'h14497,4);
TASK_PP(16'h14498,4);
TASK_PP(16'h14499,4);
TASK_PP(16'h1449A,4);
TASK_PP(16'h1449B,4);
TASK_PP(16'h1449C,4);
TASK_PP(16'h1449D,4);
TASK_PP(16'h1449E,4);
TASK_PP(16'h1449F,4);
TASK_PP(16'h144A0,4);
TASK_PP(16'h144A1,4);
TASK_PP(16'h144A2,4);
TASK_PP(16'h144A3,4);
TASK_PP(16'h144A4,4);
TASK_PP(16'h144A5,4);
TASK_PP(16'h144A6,4);
TASK_PP(16'h144A7,4);
TASK_PP(16'h144A8,4);
TASK_PP(16'h144A9,4);
TASK_PP(16'h144AA,4);
TASK_PP(16'h144AB,4);
TASK_PP(16'h144AC,4);
TASK_PP(16'h144AD,4);
TASK_PP(16'h144AE,4);
TASK_PP(16'h144AF,4);
TASK_PP(16'h144B0,4);
TASK_PP(16'h144B1,4);
TASK_PP(16'h144B2,4);
TASK_PP(16'h144B3,4);
TASK_PP(16'h144B4,4);
TASK_PP(16'h144B5,4);
TASK_PP(16'h144B6,4);
TASK_PP(16'h144B7,4);
TASK_PP(16'h144B8,4);
TASK_PP(16'h144B9,4);
TASK_PP(16'h144BA,4);
TASK_PP(16'h144BB,4);
TASK_PP(16'h144BC,4);
TASK_PP(16'h144BD,4);
TASK_PP(16'h144BE,4);
TASK_PP(16'h144BF,4);
TASK_PP(16'h144C0,4);
TASK_PP(16'h144C1,4);
TASK_PP(16'h144C2,4);
TASK_PP(16'h144C3,4);
TASK_PP(16'h144C4,4);
TASK_PP(16'h144C5,4);
TASK_PP(16'h144C6,4);
TASK_PP(16'h144C7,4);
TASK_PP(16'h144C8,4);
TASK_PP(16'h144C9,4);
TASK_PP(16'h144CA,4);
TASK_PP(16'h144CB,4);
TASK_PP(16'h144CC,4);
TASK_PP(16'h144CD,4);
TASK_PP(16'h144CE,4);
TASK_PP(16'h144CF,4);
TASK_PP(16'h144D0,4);
TASK_PP(16'h144D1,4);
TASK_PP(16'h144D2,4);
TASK_PP(16'h144D3,4);
TASK_PP(16'h144D4,4);
TASK_PP(16'h144D5,4);
TASK_PP(16'h144D6,4);
TASK_PP(16'h144D7,4);
TASK_PP(16'h144D8,4);
TASK_PP(16'h144D9,4);
TASK_PP(16'h144DA,4);
TASK_PP(16'h144DB,4);
TASK_PP(16'h144DC,4);
TASK_PP(16'h144DD,4);
TASK_PP(16'h144DE,4);
TASK_PP(16'h144DF,4);
TASK_PP(16'h144E0,4);
TASK_PP(16'h144E1,4);
TASK_PP(16'h144E2,4);
TASK_PP(16'h144E3,4);
TASK_PP(16'h144E4,4);
TASK_PP(16'h144E5,4);
TASK_PP(16'h144E6,4);
TASK_PP(16'h144E7,4);
TASK_PP(16'h144E8,4);
TASK_PP(16'h144E9,4);
TASK_PP(16'h144EA,4);
TASK_PP(16'h144EB,4);
TASK_PP(16'h144EC,4);
TASK_PP(16'h144ED,4);
TASK_PP(16'h144EE,4);
TASK_PP(16'h144EF,4);
TASK_PP(16'h144F0,4);
TASK_PP(16'h144F1,4);
TASK_PP(16'h144F2,4);
TASK_PP(16'h144F3,4);
TASK_PP(16'h144F4,4);
TASK_PP(16'h144F5,4);
TASK_PP(16'h144F6,4);
TASK_PP(16'h144F7,4);
TASK_PP(16'h144F8,4);
TASK_PP(16'h144F9,4);
TASK_PP(16'h144FA,4);
TASK_PP(16'h144FB,4);
TASK_PP(16'h144FC,4);
TASK_PP(16'h144FD,4);
TASK_PP(16'h144FE,4);
TASK_PP(16'h144FF,4);
TASK_PP(16'h14500,4);
TASK_PP(16'h14501,4);
TASK_PP(16'h14502,4);
TASK_PP(16'h14503,4);
TASK_PP(16'h14504,4);
TASK_PP(16'h14505,4);
TASK_PP(16'h14506,4);
TASK_PP(16'h14507,4);
TASK_PP(16'h14508,4);
TASK_PP(16'h14509,4);
TASK_PP(16'h1450A,4);
TASK_PP(16'h1450B,4);
TASK_PP(16'h1450C,4);
TASK_PP(16'h1450D,4);
TASK_PP(16'h1450E,4);
TASK_PP(16'h1450F,4);
TASK_PP(16'h14510,4);
TASK_PP(16'h14511,4);
TASK_PP(16'h14512,4);
TASK_PP(16'h14513,4);
TASK_PP(16'h14514,4);
TASK_PP(16'h14515,4);
TASK_PP(16'h14516,4);
TASK_PP(16'h14517,4);
TASK_PP(16'h14518,4);
TASK_PP(16'h14519,4);
TASK_PP(16'h1451A,4);
TASK_PP(16'h1451B,4);
TASK_PP(16'h1451C,4);
TASK_PP(16'h1451D,4);
TASK_PP(16'h1451E,4);
TASK_PP(16'h1451F,4);
TASK_PP(16'h14520,4);
TASK_PP(16'h14521,4);
TASK_PP(16'h14522,4);
TASK_PP(16'h14523,4);
TASK_PP(16'h14524,4);
TASK_PP(16'h14525,4);
TASK_PP(16'h14526,4);
TASK_PP(16'h14527,4);
TASK_PP(16'h14528,4);
TASK_PP(16'h14529,4);
TASK_PP(16'h1452A,4);
TASK_PP(16'h1452B,4);
TASK_PP(16'h1452C,4);
TASK_PP(16'h1452D,4);
TASK_PP(16'h1452E,4);
TASK_PP(16'h1452F,4);
TASK_PP(16'h14530,4);
TASK_PP(16'h14531,4);
TASK_PP(16'h14532,4);
TASK_PP(16'h14533,4);
TASK_PP(16'h14534,4);
TASK_PP(16'h14535,4);
TASK_PP(16'h14536,4);
TASK_PP(16'h14537,4);
TASK_PP(16'h14538,4);
TASK_PP(16'h14539,4);
TASK_PP(16'h1453A,4);
TASK_PP(16'h1453B,4);
TASK_PP(16'h1453C,4);
TASK_PP(16'h1453D,4);
TASK_PP(16'h1453E,4);
TASK_PP(16'h1453F,4);
TASK_PP(16'h14540,4);
TASK_PP(16'h14541,4);
TASK_PP(16'h14542,4);
TASK_PP(16'h14543,4);
TASK_PP(16'h14544,4);
TASK_PP(16'h14545,4);
TASK_PP(16'h14546,4);
TASK_PP(16'h14547,4);
TASK_PP(16'h14548,4);
TASK_PP(16'h14549,4);
TASK_PP(16'h1454A,4);
TASK_PP(16'h1454B,4);
TASK_PP(16'h1454C,4);
TASK_PP(16'h1454D,4);
TASK_PP(16'h1454E,4);
TASK_PP(16'h1454F,4);
TASK_PP(16'h14550,4);
TASK_PP(16'h14551,4);
TASK_PP(16'h14552,4);
TASK_PP(16'h14553,4);
TASK_PP(16'h14554,4);
TASK_PP(16'h14555,4);
TASK_PP(16'h14556,4);
TASK_PP(16'h14557,4);
TASK_PP(16'h14558,4);
TASK_PP(16'h14559,4);
TASK_PP(16'h1455A,4);
TASK_PP(16'h1455B,4);
TASK_PP(16'h1455C,4);
TASK_PP(16'h1455D,4);
TASK_PP(16'h1455E,4);
TASK_PP(16'h1455F,4);
TASK_PP(16'h14560,4);
TASK_PP(16'h14561,4);
TASK_PP(16'h14562,4);
TASK_PP(16'h14563,4);
TASK_PP(16'h14564,4);
TASK_PP(16'h14565,4);
TASK_PP(16'h14566,4);
TASK_PP(16'h14567,4);
TASK_PP(16'h14568,4);
TASK_PP(16'h14569,4);
TASK_PP(16'h1456A,4);
TASK_PP(16'h1456B,4);
TASK_PP(16'h1456C,4);
TASK_PP(16'h1456D,4);
TASK_PP(16'h1456E,4);
TASK_PP(16'h1456F,4);
TASK_PP(16'h14570,4);
TASK_PP(16'h14571,4);
TASK_PP(16'h14572,4);
TASK_PP(16'h14573,4);
TASK_PP(16'h14574,4);
TASK_PP(16'h14575,4);
TASK_PP(16'h14576,4);
TASK_PP(16'h14577,4);
TASK_PP(16'h14578,4);
TASK_PP(16'h14579,4);
TASK_PP(16'h1457A,4);
TASK_PP(16'h1457B,4);
TASK_PP(16'h1457C,4);
TASK_PP(16'h1457D,4);
TASK_PP(16'h1457E,4);
TASK_PP(16'h1457F,4);
TASK_PP(16'h14580,4);
TASK_PP(16'h14581,4);
TASK_PP(16'h14582,4);
TASK_PP(16'h14583,4);
TASK_PP(16'h14584,4);
TASK_PP(16'h14585,4);
TASK_PP(16'h14586,4);
TASK_PP(16'h14587,4);
TASK_PP(16'h14588,4);
TASK_PP(16'h14589,4);
TASK_PP(16'h1458A,4);
TASK_PP(16'h1458B,4);
TASK_PP(16'h1458C,4);
TASK_PP(16'h1458D,4);
TASK_PP(16'h1458E,4);
TASK_PP(16'h1458F,4);
TASK_PP(16'h14590,4);
TASK_PP(16'h14591,4);
TASK_PP(16'h14592,4);
TASK_PP(16'h14593,4);
TASK_PP(16'h14594,4);
TASK_PP(16'h14595,4);
TASK_PP(16'h14596,4);
TASK_PP(16'h14597,4);
TASK_PP(16'h14598,4);
TASK_PP(16'h14599,4);
TASK_PP(16'h1459A,4);
TASK_PP(16'h1459B,4);
TASK_PP(16'h1459C,4);
TASK_PP(16'h1459D,4);
TASK_PP(16'h1459E,4);
TASK_PP(16'h1459F,4);
TASK_PP(16'h145A0,4);
TASK_PP(16'h145A1,4);
TASK_PP(16'h145A2,4);
TASK_PP(16'h145A3,4);
TASK_PP(16'h145A4,4);
TASK_PP(16'h145A5,4);
TASK_PP(16'h145A6,4);
TASK_PP(16'h145A7,4);
TASK_PP(16'h145A8,4);
TASK_PP(16'h145A9,4);
TASK_PP(16'h145AA,4);
TASK_PP(16'h145AB,4);
TASK_PP(16'h145AC,4);
TASK_PP(16'h145AD,4);
TASK_PP(16'h145AE,4);
TASK_PP(16'h145AF,4);
TASK_PP(16'h145B0,4);
TASK_PP(16'h145B1,4);
TASK_PP(16'h145B2,4);
TASK_PP(16'h145B3,4);
TASK_PP(16'h145B4,4);
TASK_PP(16'h145B5,4);
TASK_PP(16'h145B6,4);
TASK_PP(16'h145B7,4);
TASK_PP(16'h145B8,4);
TASK_PP(16'h145B9,4);
TASK_PP(16'h145BA,4);
TASK_PP(16'h145BB,4);
TASK_PP(16'h145BC,4);
TASK_PP(16'h145BD,4);
TASK_PP(16'h145BE,4);
TASK_PP(16'h145BF,4);
TASK_PP(16'h145C0,4);
TASK_PP(16'h145C1,4);
TASK_PP(16'h145C2,4);
TASK_PP(16'h145C3,4);
TASK_PP(16'h145C4,4);
TASK_PP(16'h145C5,4);
TASK_PP(16'h145C6,4);
TASK_PP(16'h145C7,4);
TASK_PP(16'h145C8,4);
TASK_PP(16'h145C9,4);
TASK_PP(16'h145CA,4);
TASK_PP(16'h145CB,4);
TASK_PP(16'h145CC,4);
TASK_PP(16'h145CD,4);
TASK_PP(16'h145CE,4);
TASK_PP(16'h145CF,4);
TASK_PP(16'h145D0,4);
TASK_PP(16'h145D1,4);
TASK_PP(16'h145D2,4);
TASK_PP(16'h145D3,4);
TASK_PP(16'h145D4,4);
TASK_PP(16'h145D5,4);
TASK_PP(16'h145D6,4);
TASK_PP(16'h145D7,4);
TASK_PP(16'h145D8,4);
TASK_PP(16'h145D9,4);
TASK_PP(16'h145DA,4);
TASK_PP(16'h145DB,4);
TASK_PP(16'h145DC,4);
TASK_PP(16'h145DD,4);
TASK_PP(16'h145DE,4);
TASK_PP(16'h145DF,4);
TASK_PP(16'h145E0,4);
TASK_PP(16'h145E1,4);
TASK_PP(16'h145E2,4);
TASK_PP(16'h145E3,4);
TASK_PP(16'h145E4,4);
TASK_PP(16'h145E5,4);
TASK_PP(16'h145E6,4);
TASK_PP(16'h145E7,4);
TASK_PP(16'h145E8,4);
TASK_PP(16'h145E9,4);
TASK_PP(16'h145EA,4);
TASK_PP(16'h145EB,4);
TASK_PP(16'h145EC,4);
TASK_PP(16'h145ED,4);
TASK_PP(16'h145EE,4);
TASK_PP(16'h145EF,4);
TASK_PP(16'h145F0,4);
TASK_PP(16'h145F1,4);
TASK_PP(16'h145F2,4);
TASK_PP(16'h145F3,4);
TASK_PP(16'h145F4,4);
TASK_PP(16'h145F5,4);
TASK_PP(16'h145F6,4);
TASK_PP(16'h145F7,4);
TASK_PP(16'h145F8,4);
TASK_PP(16'h145F9,4);
TASK_PP(16'h145FA,4);
TASK_PP(16'h145FB,4);
TASK_PP(16'h145FC,4);
TASK_PP(16'h145FD,4);
TASK_PP(16'h145FE,4);
TASK_PP(16'h145FF,4);
TASK_PP(16'h14600,4);
TASK_PP(16'h14601,4);
TASK_PP(16'h14602,4);
TASK_PP(16'h14603,4);
TASK_PP(16'h14604,4);
TASK_PP(16'h14605,4);
TASK_PP(16'h14606,4);
TASK_PP(16'h14607,4);
TASK_PP(16'h14608,4);
TASK_PP(16'h14609,4);
TASK_PP(16'h1460A,4);
TASK_PP(16'h1460B,4);
TASK_PP(16'h1460C,4);
TASK_PP(16'h1460D,4);
TASK_PP(16'h1460E,4);
TASK_PP(16'h1460F,4);
TASK_PP(16'h14610,4);
TASK_PP(16'h14611,4);
TASK_PP(16'h14612,4);
TASK_PP(16'h14613,4);
TASK_PP(16'h14614,4);
TASK_PP(16'h14615,4);
TASK_PP(16'h14616,4);
TASK_PP(16'h14617,4);
TASK_PP(16'h14618,4);
TASK_PP(16'h14619,4);
TASK_PP(16'h1461A,4);
TASK_PP(16'h1461B,4);
TASK_PP(16'h1461C,4);
TASK_PP(16'h1461D,4);
TASK_PP(16'h1461E,4);
TASK_PP(16'h1461F,4);
TASK_PP(16'h14620,4);
TASK_PP(16'h14621,4);
TASK_PP(16'h14622,4);
TASK_PP(16'h14623,4);
TASK_PP(16'h14624,4);
TASK_PP(16'h14625,4);
TASK_PP(16'h14626,4);
TASK_PP(16'h14627,4);
TASK_PP(16'h14628,4);
TASK_PP(16'h14629,4);
TASK_PP(16'h1462A,4);
TASK_PP(16'h1462B,4);
TASK_PP(16'h1462C,4);
TASK_PP(16'h1462D,4);
TASK_PP(16'h1462E,4);
TASK_PP(16'h1462F,4);
TASK_PP(16'h14630,4);
TASK_PP(16'h14631,4);
TASK_PP(16'h14632,4);
TASK_PP(16'h14633,4);
TASK_PP(16'h14634,4);
TASK_PP(16'h14635,4);
TASK_PP(16'h14636,4);
TASK_PP(16'h14637,4);
TASK_PP(16'h14638,4);
TASK_PP(16'h14639,4);
TASK_PP(16'h1463A,4);
TASK_PP(16'h1463B,4);
TASK_PP(16'h1463C,4);
TASK_PP(16'h1463D,4);
TASK_PP(16'h1463E,4);
TASK_PP(16'h1463F,4);
TASK_PP(16'h14640,4);
TASK_PP(16'h14641,4);
TASK_PP(16'h14642,4);
TASK_PP(16'h14643,4);
TASK_PP(16'h14644,4);
TASK_PP(16'h14645,4);
TASK_PP(16'h14646,4);
TASK_PP(16'h14647,4);
TASK_PP(16'h14648,4);
TASK_PP(16'h14649,4);
TASK_PP(16'h1464A,4);
TASK_PP(16'h1464B,4);
TASK_PP(16'h1464C,4);
TASK_PP(16'h1464D,4);
TASK_PP(16'h1464E,4);
TASK_PP(16'h1464F,4);
TASK_PP(16'h14650,4);
TASK_PP(16'h14651,4);
TASK_PP(16'h14652,4);
TASK_PP(16'h14653,4);
TASK_PP(16'h14654,4);
TASK_PP(16'h14655,4);
TASK_PP(16'h14656,4);
TASK_PP(16'h14657,4);
TASK_PP(16'h14658,4);
TASK_PP(16'h14659,4);
TASK_PP(16'h1465A,4);
TASK_PP(16'h1465B,4);
TASK_PP(16'h1465C,4);
TASK_PP(16'h1465D,4);
TASK_PP(16'h1465E,4);
TASK_PP(16'h1465F,4);
TASK_PP(16'h14660,4);
TASK_PP(16'h14661,4);
TASK_PP(16'h14662,4);
TASK_PP(16'h14663,4);
TASK_PP(16'h14664,4);
TASK_PP(16'h14665,4);
TASK_PP(16'h14666,4);
TASK_PP(16'h14667,4);
TASK_PP(16'h14668,4);
TASK_PP(16'h14669,4);
TASK_PP(16'h1466A,4);
TASK_PP(16'h1466B,4);
TASK_PP(16'h1466C,4);
TASK_PP(16'h1466D,4);
TASK_PP(16'h1466E,4);
TASK_PP(16'h1466F,4);
TASK_PP(16'h14670,4);
TASK_PP(16'h14671,4);
TASK_PP(16'h14672,4);
TASK_PP(16'h14673,4);
TASK_PP(16'h14674,4);
TASK_PP(16'h14675,4);
TASK_PP(16'h14676,4);
TASK_PP(16'h14677,4);
TASK_PP(16'h14678,4);
TASK_PP(16'h14679,4);
TASK_PP(16'h1467A,4);
TASK_PP(16'h1467B,4);
TASK_PP(16'h1467C,4);
TASK_PP(16'h1467D,4);
TASK_PP(16'h1467E,4);
TASK_PP(16'h1467F,4);
TASK_PP(16'h14680,4);
TASK_PP(16'h14681,4);
TASK_PP(16'h14682,4);
TASK_PP(16'h14683,4);
TASK_PP(16'h14684,4);
TASK_PP(16'h14685,4);
TASK_PP(16'h14686,4);
TASK_PP(16'h14687,4);
TASK_PP(16'h14688,4);
TASK_PP(16'h14689,4);
TASK_PP(16'h1468A,4);
TASK_PP(16'h1468B,4);
TASK_PP(16'h1468C,4);
TASK_PP(16'h1468D,4);
TASK_PP(16'h1468E,4);
TASK_PP(16'h1468F,4);
TASK_PP(16'h14690,4);
TASK_PP(16'h14691,4);
TASK_PP(16'h14692,4);
TASK_PP(16'h14693,4);
TASK_PP(16'h14694,4);
TASK_PP(16'h14695,4);
TASK_PP(16'h14696,4);
TASK_PP(16'h14697,4);
TASK_PP(16'h14698,4);
TASK_PP(16'h14699,4);
TASK_PP(16'h1469A,4);
TASK_PP(16'h1469B,4);
TASK_PP(16'h1469C,4);
TASK_PP(16'h1469D,4);
TASK_PP(16'h1469E,4);
TASK_PP(16'h1469F,4);
TASK_PP(16'h146A0,4);
TASK_PP(16'h146A1,4);
TASK_PP(16'h146A2,4);
TASK_PP(16'h146A3,4);
TASK_PP(16'h146A4,4);
TASK_PP(16'h146A5,4);
TASK_PP(16'h146A6,4);
TASK_PP(16'h146A7,4);
TASK_PP(16'h146A8,4);
TASK_PP(16'h146A9,4);
TASK_PP(16'h146AA,4);
TASK_PP(16'h146AB,4);
TASK_PP(16'h146AC,4);
TASK_PP(16'h146AD,4);
TASK_PP(16'h146AE,4);
TASK_PP(16'h146AF,4);
TASK_PP(16'h146B0,4);
TASK_PP(16'h146B1,4);
TASK_PP(16'h146B2,4);
TASK_PP(16'h146B3,4);
TASK_PP(16'h146B4,4);
TASK_PP(16'h146B5,4);
TASK_PP(16'h146B6,4);
TASK_PP(16'h146B7,4);
TASK_PP(16'h146B8,4);
TASK_PP(16'h146B9,4);
TASK_PP(16'h146BA,4);
TASK_PP(16'h146BB,4);
TASK_PP(16'h146BC,4);
TASK_PP(16'h146BD,4);
TASK_PP(16'h146BE,4);
TASK_PP(16'h146BF,4);
TASK_PP(16'h146C0,4);
TASK_PP(16'h146C1,4);
TASK_PP(16'h146C2,4);
TASK_PP(16'h146C3,4);
TASK_PP(16'h146C4,4);
TASK_PP(16'h146C5,4);
TASK_PP(16'h146C6,4);
TASK_PP(16'h146C7,4);
TASK_PP(16'h146C8,4);
TASK_PP(16'h146C9,4);
TASK_PP(16'h146CA,4);
TASK_PP(16'h146CB,4);
TASK_PP(16'h146CC,4);
TASK_PP(16'h146CD,4);
TASK_PP(16'h146CE,4);
TASK_PP(16'h146CF,4);
TASK_PP(16'h146D0,4);
TASK_PP(16'h146D1,4);
TASK_PP(16'h146D2,4);
TASK_PP(16'h146D3,4);
TASK_PP(16'h146D4,4);
TASK_PP(16'h146D5,4);
TASK_PP(16'h146D6,4);
TASK_PP(16'h146D7,4);
TASK_PP(16'h146D8,4);
TASK_PP(16'h146D9,4);
TASK_PP(16'h146DA,4);
TASK_PP(16'h146DB,4);
TASK_PP(16'h146DC,4);
TASK_PP(16'h146DD,4);
TASK_PP(16'h146DE,4);
TASK_PP(16'h146DF,4);
TASK_PP(16'h146E0,4);
TASK_PP(16'h146E1,4);
TASK_PP(16'h146E2,4);
TASK_PP(16'h146E3,4);
TASK_PP(16'h146E4,4);
TASK_PP(16'h146E5,4);
TASK_PP(16'h146E6,4);
TASK_PP(16'h146E7,4);
TASK_PP(16'h146E8,4);
TASK_PP(16'h146E9,4);
TASK_PP(16'h146EA,4);
TASK_PP(16'h146EB,4);
TASK_PP(16'h146EC,4);
TASK_PP(16'h146ED,4);
TASK_PP(16'h146EE,4);
TASK_PP(16'h146EF,4);
TASK_PP(16'h146F0,4);
TASK_PP(16'h146F1,4);
TASK_PP(16'h146F2,4);
TASK_PP(16'h146F3,4);
TASK_PP(16'h146F4,4);
TASK_PP(16'h146F5,4);
TASK_PP(16'h146F6,4);
TASK_PP(16'h146F7,4);
TASK_PP(16'h146F8,4);
TASK_PP(16'h146F9,4);
TASK_PP(16'h146FA,4);
TASK_PP(16'h146FB,4);
TASK_PP(16'h146FC,4);
TASK_PP(16'h146FD,4);
TASK_PP(16'h146FE,4);
TASK_PP(16'h146FF,4);
TASK_PP(16'h14700,4);
TASK_PP(16'h14701,4);
TASK_PP(16'h14702,4);
TASK_PP(16'h14703,4);
TASK_PP(16'h14704,4);
TASK_PP(16'h14705,4);
TASK_PP(16'h14706,4);
TASK_PP(16'h14707,4);
TASK_PP(16'h14708,4);
TASK_PP(16'h14709,4);
TASK_PP(16'h1470A,4);
TASK_PP(16'h1470B,4);
TASK_PP(16'h1470C,4);
TASK_PP(16'h1470D,4);
TASK_PP(16'h1470E,4);
TASK_PP(16'h1470F,4);
TASK_PP(16'h14710,4);
TASK_PP(16'h14711,4);
TASK_PP(16'h14712,4);
TASK_PP(16'h14713,4);
TASK_PP(16'h14714,4);
TASK_PP(16'h14715,4);
TASK_PP(16'h14716,4);
TASK_PP(16'h14717,4);
TASK_PP(16'h14718,4);
TASK_PP(16'h14719,4);
TASK_PP(16'h1471A,4);
TASK_PP(16'h1471B,4);
TASK_PP(16'h1471C,4);
TASK_PP(16'h1471D,4);
TASK_PP(16'h1471E,4);
TASK_PP(16'h1471F,4);
TASK_PP(16'h14720,4);
TASK_PP(16'h14721,4);
TASK_PP(16'h14722,4);
TASK_PP(16'h14723,4);
TASK_PP(16'h14724,4);
TASK_PP(16'h14725,4);
TASK_PP(16'h14726,4);
TASK_PP(16'h14727,4);
TASK_PP(16'h14728,4);
TASK_PP(16'h14729,4);
TASK_PP(16'h1472A,4);
TASK_PP(16'h1472B,4);
TASK_PP(16'h1472C,4);
TASK_PP(16'h1472D,4);
TASK_PP(16'h1472E,4);
TASK_PP(16'h1472F,4);
TASK_PP(16'h14730,4);
TASK_PP(16'h14731,4);
TASK_PP(16'h14732,4);
TASK_PP(16'h14733,4);
TASK_PP(16'h14734,4);
TASK_PP(16'h14735,4);
TASK_PP(16'h14736,4);
TASK_PP(16'h14737,4);
TASK_PP(16'h14738,4);
TASK_PP(16'h14739,4);
TASK_PP(16'h1473A,4);
TASK_PP(16'h1473B,4);
TASK_PP(16'h1473C,4);
TASK_PP(16'h1473D,4);
TASK_PP(16'h1473E,4);
TASK_PP(16'h1473F,4);
TASK_PP(16'h14740,4);
TASK_PP(16'h14741,4);
TASK_PP(16'h14742,4);
TASK_PP(16'h14743,4);
TASK_PP(16'h14744,4);
TASK_PP(16'h14745,4);
TASK_PP(16'h14746,4);
TASK_PP(16'h14747,4);
TASK_PP(16'h14748,4);
TASK_PP(16'h14749,4);
TASK_PP(16'h1474A,4);
TASK_PP(16'h1474B,4);
TASK_PP(16'h1474C,4);
TASK_PP(16'h1474D,4);
TASK_PP(16'h1474E,4);
TASK_PP(16'h1474F,4);
TASK_PP(16'h14750,4);
TASK_PP(16'h14751,4);
TASK_PP(16'h14752,4);
TASK_PP(16'h14753,4);
TASK_PP(16'h14754,4);
TASK_PP(16'h14755,4);
TASK_PP(16'h14756,4);
TASK_PP(16'h14757,4);
TASK_PP(16'h14758,4);
TASK_PP(16'h14759,4);
TASK_PP(16'h1475A,4);
TASK_PP(16'h1475B,4);
TASK_PP(16'h1475C,4);
TASK_PP(16'h1475D,4);
TASK_PP(16'h1475E,4);
TASK_PP(16'h1475F,4);
TASK_PP(16'h14760,4);
TASK_PP(16'h14761,4);
TASK_PP(16'h14762,4);
TASK_PP(16'h14763,4);
TASK_PP(16'h14764,4);
TASK_PP(16'h14765,4);
TASK_PP(16'h14766,4);
TASK_PP(16'h14767,4);
TASK_PP(16'h14768,4);
TASK_PP(16'h14769,4);
TASK_PP(16'h1476A,4);
TASK_PP(16'h1476B,4);
TASK_PP(16'h1476C,4);
TASK_PP(16'h1476D,4);
TASK_PP(16'h1476E,4);
TASK_PP(16'h1476F,4);
TASK_PP(16'h14770,4);
TASK_PP(16'h14771,4);
TASK_PP(16'h14772,4);
TASK_PP(16'h14773,4);
TASK_PP(16'h14774,4);
TASK_PP(16'h14775,4);
TASK_PP(16'h14776,4);
TASK_PP(16'h14777,4);
TASK_PP(16'h14778,4);
TASK_PP(16'h14779,4);
TASK_PP(16'h1477A,4);
TASK_PP(16'h1477B,4);
TASK_PP(16'h1477C,4);
TASK_PP(16'h1477D,4);
TASK_PP(16'h1477E,4);
TASK_PP(16'h1477F,4);
TASK_PP(16'h14780,4);
TASK_PP(16'h14781,4);
TASK_PP(16'h14782,4);
TASK_PP(16'h14783,4);
TASK_PP(16'h14784,4);
TASK_PP(16'h14785,4);
TASK_PP(16'h14786,4);
TASK_PP(16'h14787,4);
TASK_PP(16'h14788,4);
TASK_PP(16'h14789,4);
TASK_PP(16'h1478A,4);
TASK_PP(16'h1478B,4);
TASK_PP(16'h1478C,4);
TASK_PP(16'h1478D,4);
TASK_PP(16'h1478E,4);
TASK_PP(16'h1478F,4);
TASK_PP(16'h14790,4);
TASK_PP(16'h14791,4);
TASK_PP(16'h14792,4);
TASK_PP(16'h14793,4);
TASK_PP(16'h14794,4);
TASK_PP(16'h14795,4);
TASK_PP(16'h14796,4);
TASK_PP(16'h14797,4);
TASK_PP(16'h14798,4);
TASK_PP(16'h14799,4);
TASK_PP(16'h1479A,4);
TASK_PP(16'h1479B,4);
TASK_PP(16'h1479C,4);
TASK_PP(16'h1479D,4);
TASK_PP(16'h1479E,4);
TASK_PP(16'h1479F,4);
TASK_PP(16'h147A0,4);
TASK_PP(16'h147A1,4);
TASK_PP(16'h147A2,4);
TASK_PP(16'h147A3,4);
TASK_PP(16'h147A4,4);
TASK_PP(16'h147A5,4);
TASK_PP(16'h147A6,4);
TASK_PP(16'h147A7,4);
TASK_PP(16'h147A8,4);
TASK_PP(16'h147A9,4);
TASK_PP(16'h147AA,4);
TASK_PP(16'h147AB,4);
TASK_PP(16'h147AC,4);
TASK_PP(16'h147AD,4);
TASK_PP(16'h147AE,4);
TASK_PP(16'h147AF,4);
TASK_PP(16'h147B0,4);
TASK_PP(16'h147B1,4);
TASK_PP(16'h147B2,4);
TASK_PP(16'h147B3,4);
TASK_PP(16'h147B4,4);
TASK_PP(16'h147B5,4);
TASK_PP(16'h147B6,4);
TASK_PP(16'h147B7,4);
TASK_PP(16'h147B8,4);
TASK_PP(16'h147B9,4);
TASK_PP(16'h147BA,4);
TASK_PP(16'h147BB,4);
TASK_PP(16'h147BC,4);
TASK_PP(16'h147BD,4);
TASK_PP(16'h147BE,4);
TASK_PP(16'h147BF,4);
TASK_PP(16'h147C0,4);
TASK_PP(16'h147C1,4);
TASK_PP(16'h147C2,4);
TASK_PP(16'h147C3,4);
TASK_PP(16'h147C4,4);
TASK_PP(16'h147C5,4);
TASK_PP(16'h147C6,4);
TASK_PP(16'h147C7,4);
TASK_PP(16'h147C8,4);
TASK_PP(16'h147C9,4);
TASK_PP(16'h147CA,4);
TASK_PP(16'h147CB,4);
TASK_PP(16'h147CC,4);
TASK_PP(16'h147CD,4);
TASK_PP(16'h147CE,4);
TASK_PP(16'h147CF,4);
TASK_PP(16'h147D0,4);
TASK_PP(16'h147D1,4);
TASK_PP(16'h147D2,4);
TASK_PP(16'h147D3,4);
TASK_PP(16'h147D4,4);
TASK_PP(16'h147D5,4);
TASK_PP(16'h147D6,4);
TASK_PP(16'h147D7,4);
TASK_PP(16'h147D8,4);
TASK_PP(16'h147D9,4);
TASK_PP(16'h147DA,4);
TASK_PP(16'h147DB,4);
TASK_PP(16'h147DC,4);
TASK_PP(16'h147DD,4);
TASK_PP(16'h147DE,4);
TASK_PP(16'h147DF,4);
TASK_PP(16'h147E0,4);
TASK_PP(16'h147E1,4);
TASK_PP(16'h147E2,4);
TASK_PP(16'h147E3,4);
TASK_PP(16'h147E4,4);
TASK_PP(16'h147E5,4);
TASK_PP(16'h147E6,4);
TASK_PP(16'h147E7,4);
TASK_PP(16'h147E8,4);
TASK_PP(16'h147E9,4);
TASK_PP(16'h147EA,4);
TASK_PP(16'h147EB,4);
TASK_PP(16'h147EC,4);
TASK_PP(16'h147ED,4);
TASK_PP(16'h147EE,4);
TASK_PP(16'h147EF,4);
TASK_PP(16'h147F0,4);
TASK_PP(16'h147F1,4);
TASK_PP(16'h147F2,4);
TASK_PP(16'h147F3,4);
TASK_PP(16'h147F4,4);
TASK_PP(16'h147F5,4);
TASK_PP(16'h147F6,4);
TASK_PP(16'h147F7,4);
TASK_PP(16'h147F8,4);
TASK_PP(16'h147F9,4);
TASK_PP(16'h147FA,4);
TASK_PP(16'h147FB,4);
TASK_PP(16'h147FC,4);
TASK_PP(16'h147FD,4);
TASK_PP(16'h147FE,4);
TASK_PP(16'h147FF,4);
TASK_PP(16'h14800,4);
TASK_PP(16'h14801,4);
TASK_PP(16'h14802,4);
TASK_PP(16'h14803,4);
TASK_PP(16'h14804,4);
TASK_PP(16'h14805,4);
TASK_PP(16'h14806,4);
TASK_PP(16'h14807,4);
TASK_PP(16'h14808,4);
TASK_PP(16'h14809,4);
TASK_PP(16'h1480A,4);
TASK_PP(16'h1480B,4);
TASK_PP(16'h1480C,4);
TASK_PP(16'h1480D,4);
TASK_PP(16'h1480E,4);
TASK_PP(16'h1480F,4);
TASK_PP(16'h14810,4);
TASK_PP(16'h14811,4);
TASK_PP(16'h14812,4);
TASK_PP(16'h14813,4);
TASK_PP(16'h14814,4);
TASK_PP(16'h14815,4);
TASK_PP(16'h14816,4);
TASK_PP(16'h14817,4);
TASK_PP(16'h14818,4);
TASK_PP(16'h14819,4);
TASK_PP(16'h1481A,4);
TASK_PP(16'h1481B,4);
TASK_PP(16'h1481C,4);
TASK_PP(16'h1481D,4);
TASK_PP(16'h1481E,4);
TASK_PP(16'h1481F,4);
TASK_PP(16'h14820,4);
TASK_PP(16'h14821,4);
TASK_PP(16'h14822,4);
TASK_PP(16'h14823,4);
TASK_PP(16'h14824,4);
TASK_PP(16'h14825,4);
TASK_PP(16'h14826,4);
TASK_PP(16'h14827,4);
TASK_PP(16'h14828,4);
TASK_PP(16'h14829,4);
TASK_PP(16'h1482A,4);
TASK_PP(16'h1482B,4);
TASK_PP(16'h1482C,4);
TASK_PP(16'h1482D,4);
TASK_PP(16'h1482E,4);
TASK_PP(16'h1482F,4);
TASK_PP(16'h14830,4);
TASK_PP(16'h14831,4);
TASK_PP(16'h14832,4);
TASK_PP(16'h14833,4);
TASK_PP(16'h14834,4);
TASK_PP(16'h14835,4);
TASK_PP(16'h14836,4);
TASK_PP(16'h14837,4);
TASK_PP(16'h14838,4);
TASK_PP(16'h14839,4);
TASK_PP(16'h1483A,4);
TASK_PP(16'h1483B,4);
TASK_PP(16'h1483C,4);
TASK_PP(16'h1483D,4);
TASK_PP(16'h1483E,4);
TASK_PP(16'h1483F,4);
TASK_PP(16'h14840,4);
TASK_PP(16'h14841,4);
TASK_PP(16'h14842,4);
TASK_PP(16'h14843,4);
TASK_PP(16'h14844,4);
TASK_PP(16'h14845,4);
TASK_PP(16'h14846,4);
TASK_PP(16'h14847,4);
TASK_PP(16'h14848,4);
TASK_PP(16'h14849,4);
TASK_PP(16'h1484A,4);
TASK_PP(16'h1484B,4);
TASK_PP(16'h1484C,4);
TASK_PP(16'h1484D,4);
TASK_PP(16'h1484E,4);
TASK_PP(16'h1484F,4);
TASK_PP(16'h14850,4);
TASK_PP(16'h14851,4);
TASK_PP(16'h14852,4);
TASK_PP(16'h14853,4);
TASK_PP(16'h14854,4);
TASK_PP(16'h14855,4);
TASK_PP(16'h14856,4);
TASK_PP(16'h14857,4);
TASK_PP(16'h14858,4);
TASK_PP(16'h14859,4);
TASK_PP(16'h1485A,4);
TASK_PP(16'h1485B,4);
TASK_PP(16'h1485C,4);
TASK_PP(16'h1485D,4);
TASK_PP(16'h1485E,4);
TASK_PP(16'h1485F,4);
TASK_PP(16'h14860,4);
TASK_PP(16'h14861,4);
TASK_PP(16'h14862,4);
TASK_PP(16'h14863,4);
TASK_PP(16'h14864,4);
TASK_PP(16'h14865,4);
TASK_PP(16'h14866,4);
TASK_PP(16'h14867,4);
TASK_PP(16'h14868,4);
TASK_PP(16'h14869,4);
TASK_PP(16'h1486A,4);
TASK_PP(16'h1486B,4);
TASK_PP(16'h1486C,4);
TASK_PP(16'h1486D,4);
TASK_PP(16'h1486E,4);
TASK_PP(16'h1486F,4);
TASK_PP(16'h14870,4);
TASK_PP(16'h14871,4);
TASK_PP(16'h14872,4);
TASK_PP(16'h14873,4);
TASK_PP(16'h14874,4);
TASK_PP(16'h14875,4);
TASK_PP(16'h14876,4);
TASK_PP(16'h14877,4);
TASK_PP(16'h14878,4);
TASK_PP(16'h14879,4);
TASK_PP(16'h1487A,4);
TASK_PP(16'h1487B,4);
TASK_PP(16'h1487C,4);
TASK_PP(16'h1487D,4);
TASK_PP(16'h1487E,4);
TASK_PP(16'h1487F,4);
TASK_PP(16'h14880,4);
TASK_PP(16'h14881,4);
TASK_PP(16'h14882,4);
TASK_PP(16'h14883,4);
TASK_PP(16'h14884,4);
TASK_PP(16'h14885,4);
TASK_PP(16'h14886,4);
TASK_PP(16'h14887,4);
TASK_PP(16'h14888,4);
TASK_PP(16'h14889,4);
TASK_PP(16'h1488A,4);
TASK_PP(16'h1488B,4);
TASK_PP(16'h1488C,4);
TASK_PP(16'h1488D,4);
TASK_PP(16'h1488E,4);
TASK_PP(16'h1488F,4);
TASK_PP(16'h14890,4);
TASK_PP(16'h14891,4);
TASK_PP(16'h14892,4);
TASK_PP(16'h14893,4);
TASK_PP(16'h14894,4);
TASK_PP(16'h14895,4);
TASK_PP(16'h14896,4);
TASK_PP(16'h14897,4);
TASK_PP(16'h14898,4);
TASK_PP(16'h14899,4);
TASK_PP(16'h1489A,4);
TASK_PP(16'h1489B,4);
TASK_PP(16'h1489C,4);
TASK_PP(16'h1489D,4);
TASK_PP(16'h1489E,4);
TASK_PP(16'h1489F,4);
TASK_PP(16'h148A0,4);
TASK_PP(16'h148A1,4);
TASK_PP(16'h148A2,4);
TASK_PP(16'h148A3,4);
TASK_PP(16'h148A4,4);
TASK_PP(16'h148A5,4);
TASK_PP(16'h148A6,4);
TASK_PP(16'h148A7,4);
TASK_PP(16'h148A8,4);
TASK_PP(16'h148A9,4);
TASK_PP(16'h148AA,4);
TASK_PP(16'h148AB,4);
TASK_PP(16'h148AC,4);
TASK_PP(16'h148AD,4);
TASK_PP(16'h148AE,4);
TASK_PP(16'h148AF,4);
TASK_PP(16'h148B0,4);
TASK_PP(16'h148B1,4);
TASK_PP(16'h148B2,4);
TASK_PP(16'h148B3,4);
TASK_PP(16'h148B4,4);
TASK_PP(16'h148B5,4);
TASK_PP(16'h148B6,4);
TASK_PP(16'h148B7,4);
TASK_PP(16'h148B8,4);
TASK_PP(16'h148B9,4);
TASK_PP(16'h148BA,4);
TASK_PP(16'h148BB,4);
TASK_PP(16'h148BC,4);
TASK_PP(16'h148BD,4);
TASK_PP(16'h148BE,4);
TASK_PP(16'h148BF,4);
TASK_PP(16'h148C0,4);
TASK_PP(16'h148C1,4);
TASK_PP(16'h148C2,4);
TASK_PP(16'h148C3,4);
TASK_PP(16'h148C4,4);
TASK_PP(16'h148C5,4);
TASK_PP(16'h148C6,4);
TASK_PP(16'h148C7,4);
TASK_PP(16'h148C8,4);
TASK_PP(16'h148C9,4);
TASK_PP(16'h148CA,4);
TASK_PP(16'h148CB,4);
TASK_PP(16'h148CC,4);
TASK_PP(16'h148CD,4);
TASK_PP(16'h148CE,4);
TASK_PP(16'h148CF,4);
TASK_PP(16'h148D0,4);
TASK_PP(16'h148D1,4);
TASK_PP(16'h148D2,4);
TASK_PP(16'h148D3,4);
TASK_PP(16'h148D4,4);
TASK_PP(16'h148D5,4);
TASK_PP(16'h148D6,4);
TASK_PP(16'h148D7,4);
TASK_PP(16'h148D8,4);
TASK_PP(16'h148D9,4);
TASK_PP(16'h148DA,4);
TASK_PP(16'h148DB,4);
TASK_PP(16'h148DC,4);
TASK_PP(16'h148DD,4);
TASK_PP(16'h148DE,4);
TASK_PP(16'h148DF,4);
TASK_PP(16'h148E0,4);
TASK_PP(16'h148E1,4);
TASK_PP(16'h148E2,4);
TASK_PP(16'h148E3,4);
TASK_PP(16'h148E4,4);
TASK_PP(16'h148E5,4);
TASK_PP(16'h148E6,4);
TASK_PP(16'h148E7,4);
TASK_PP(16'h148E8,4);
TASK_PP(16'h148E9,4);
TASK_PP(16'h148EA,4);
TASK_PP(16'h148EB,4);
TASK_PP(16'h148EC,4);
TASK_PP(16'h148ED,4);
TASK_PP(16'h148EE,4);
TASK_PP(16'h148EF,4);
TASK_PP(16'h148F0,4);
TASK_PP(16'h148F1,4);
TASK_PP(16'h148F2,4);
TASK_PP(16'h148F3,4);
TASK_PP(16'h148F4,4);
TASK_PP(16'h148F5,4);
TASK_PP(16'h148F6,4);
TASK_PP(16'h148F7,4);
TASK_PP(16'h148F8,4);
TASK_PP(16'h148F9,4);
TASK_PP(16'h148FA,4);
TASK_PP(16'h148FB,4);
TASK_PP(16'h148FC,4);
TASK_PP(16'h148FD,4);
TASK_PP(16'h148FE,4);
TASK_PP(16'h148FF,4);
TASK_PP(16'h14900,4);
TASK_PP(16'h14901,4);
TASK_PP(16'h14902,4);
TASK_PP(16'h14903,4);
TASK_PP(16'h14904,4);
TASK_PP(16'h14905,4);
TASK_PP(16'h14906,4);
TASK_PP(16'h14907,4);
TASK_PP(16'h14908,4);
TASK_PP(16'h14909,4);
TASK_PP(16'h1490A,4);
TASK_PP(16'h1490B,4);
TASK_PP(16'h1490C,4);
TASK_PP(16'h1490D,4);
TASK_PP(16'h1490E,4);
TASK_PP(16'h1490F,4);
TASK_PP(16'h14910,4);
TASK_PP(16'h14911,4);
TASK_PP(16'h14912,4);
TASK_PP(16'h14913,4);
TASK_PP(16'h14914,4);
TASK_PP(16'h14915,4);
TASK_PP(16'h14916,4);
TASK_PP(16'h14917,4);
TASK_PP(16'h14918,4);
TASK_PP(16'h14919,4);
TASK_PP(16'h1491A,4);
TASK_PP(16'h1491B,4);
TASK_PP(16'h1491C,4);
TASK_PP(16'h1491D,4);
TASK_PP(16'h1491E,4);
TASK_PP(16'h1491F,4);
TASK_PP(16'h14920,4);
TASK_PP(16'h14921,4);
TASK_PP(16'h14922,4);
TASK_PP(16'h14923,4);
TASK_PP(16'h14924,4);
TASK_PP(16'h14925,4);
TASK_PP(16'h14926,4);
TASK_PP(16'h14927,4);
TASK_PP(16'h14928,4);
TASK_PP(16'h14929,4);
TASK_PP(16'h1492A,4);
TASK_PP(16'h1492B,4);
TASK_PP(16'h1492C,4);
TASK_PP(16'h1492D,4);
TASK_PP(16'h1492E,4);
TASK_PP(16'h1492F,4);
TASK_PP(16'h14930,4);
TASK_PP(16'h14931,4);
TASK_PP(16'h14932,4);
TASK_PP(16'h14933,4);
TASK_PP(16'h14934,4);
TASK_PP(16'h14935,4);
TASK_PP(16'h14936,4);
TASK_PP(16'h14937,4);
TASK_PP(16'h14938,4);
TASK_PP(16'h14939,4);
TASK_PP(16'h1493A,4);
TASK_PP(16'h1493B,4);
TASK_PP(16'h1493C,4);
TASK_PP(16'h1493D,4);
TASK_PP(16'h1493E,4);
TASK_PP(16'h1493F,4);
TASK_PP(16'h14940,4);
TASK_PP(16'h14941,4);
TASK_PP(16'h14942,4);
TASK_PP(16'h14943,4);
TASK_PP(16'h14944,4);
TASK_PP(16'h14945,4);
TASK_PP(16'h14946,4);
TASK_PP(16'h14947,4);
TASK_PP(16'h14948,4);
TASK_PP(16'h14949,4);
TASK_PP(16'h1494A,4);
TASK_PP(16'h1494B,4);
TASK_PP(16'h1494C,4);
TASK_PP(16'h1494D,4);
TASK_PP(16'h1494E,4);
TASK_PP(16'h1494F,4);
TASK_PP(16'h14950,4);
TASK_PP(16'h14951,4);
TASK_PP(16'h14952,4);
TASK_PP(16'h14953,4);
TASK_PP(16'h14954,4);
TASK_PP(16'h14955,4);
TASK_PP(16'h14956,4);
TASK_PP(16'h14957,4);
TASK_PP(16'h14958,4);
TASK_PP(16'h14959,4);
TASK_PP(16'h1495A,4);
TASK_PP(16'h1495B,4);
TASK_PP(16'h1495C,4);
TASK_PP(16'h1495D,4);
TASK_PP(16'h1495E,4);
TASK_PP(16'h1495F,4);
TASK_PP(16'h14960,4);
TASK_PP(16'h14961,4);
TASK_PP(16'h14962,4);
TASK_PP(16'h14963,4);
TASK_PP(16'h14964,4);
TASK_PP(16'h14965,4);
TASK_PP(16'h14966,4);
TASK_PP(16'h14967,4);
TASK_PP(16'h14968,4);
TASK_PP(16'h14969,4);
TASK_PP(16'h1496A,4);
TASK_PP(16'h1496B,4);
TASK_PP(16'h1496C,4);
TASK_PP(16'h1496D,4);
TASK_PP(16'h1496E,4);
TASK_PP(16'h1496F,4);
TASK_PP(16'h14970,4);
TASK_PP(16'h14971,4);
TASK_PP(16'h14972,4);
TASK_PP(16'h14973,4);
TASK_PP(16'h14974,4);
TASK_PP(16'h14975,4);
TASK_PP(16'h14976,4);
TASK_PP(16'h14977,4);
TASK_PP(16'h14978,4);
TASK_PP(16'h14979,4);
TASK_PP(16'h1497A,4);
TASK_PP(16'h1497B,4);
TASK_PP(16'h1497C,4);
TASK_PP(16'h1497D,4);
TASK_PP(16'h1497E,4);
TASK_PP(16'h1497F,4);
TASK_PP(16'h14980,4);
TASK_PP(16'h14981,4);
TASK_PP(16'h14982,4);
TASK_PP(16'h14983,4);
TASK_PP(16'h14984,4);
TASK_PP(16'h14985,4);
TASK_PP(16'h14986,4);
TASK_PP(16'h14987,4);
TASK_PP(16'h14988,4);
TASK_PP(16'h14989,4);
TASK_PP(16'h1498A,4);
TASK_PP(16'h1498B,4);
TASK_PP(16'h1498C,4);
TASK_PP(16'h1498D,4);
TASK_PP(16'h1498E,4);
TASK_PP(16'h1498F,4);
TASK_PP(16'h14990,4);
TASK_PP(16'h14991,4);
TASK_PP(16'h14992,4);
TASK_PP(16'h14993,4);
TASK_PP(16'h14994,4);
TASK_PP(16'h14995,4);
TASK_PP(16'h14996,4);
TASK_PP(16'h14997,4);
TASK_PP(16'h14998,4);
TASK_PP(16'h14999,4);
TASK_PP(16'h1499A,4);
TASK_PP(16'h1499B,4);
TASK_PP(16'h1499C,4);
TASK_PP(16'h1499D,4);
TASK_PP(16'h1499E,4);
TASK_PP(16'h1499F,4);
TASK_PP(16'h149A0,4);
TASK_PP(16'h149A1,4);
TASK_PP(16'h149A2,4);
TASK_PP(16'h149A3,4);
TASK_PP(16'h149A4,4);
TASK_PP(16'h149A5,4);
TASK_PP(16'h149A6,4);
TASK_PP(16'h149A7,4);
TASK_PP(16'h149A8,4);
TASK_PP(16'h149A9,4);
TASK_PP(16'h149AA,4);
TASK_PP(16'h149AB,4);
TASK_PP(16'h149AC,4);
TASK_PP(16'h149AD,4);
TASK_PP(16'h149AE,4);
TASK_PP(16'h149AF,4);
TASK_PP(16'h149B0,4);
TASK_PP(16'h149B1,4);
TASK_PP(16'h149B2,4);
TASK_PP(16'h149B3,4);
TASK_PP(16'h149B4,4);
TASK_PP(16'h149B5,4);
TASK_PP(16'h149B6,4);
TASK_PP(16'h149B7,4);
TASK_PP(16'h149B8,4);
TASK_PP(16'h149B9,4);
TASK_PP(16'h149BA,4);
TASK_PP(16'h149BB,4);
TASK_PP(16'h149BC,4);
TASK_PP(16'h149BD,4);
TASK_PP(16'h149BE,4);
TASK_PP(16'h149BF,4);
TASK_PP(16'h149C0,4);
TASK_PP(16'h149C1,4);
TASK_PP(16'h149C2,4);
TASK_PP(16'h149C3,4);
TASK_PP(16'h149C4,4);
TASK_PP(16'h149C5,4);
TASK_PP(16'h149C6,4);
TASK_PP(16'h149C7,4);
TASK_PP(16'h149C8,4);
TASK_PP(16'h149C9,4);
TASK_PP(16'h149CA,4);
TASK_PP(16'h149CB,4);
TASK_PP(16'h149CC,4);
TASK_PP(16'h149CD,4);
TASK_PP(16'h149CE,4);
TASK_PP(16'h149CF,4);
TASK_PP(16'h149D0,4);
TASK_PP(16'h149D1,4);
TASK_PP(16'h149D2,4);
TASK_PP(16'h149D3,4);
TASK_PP(16'h149D4,4);
TASK_PP(16'h149D5,4);
TASK_PP(16'h149D6,4);
TASK_PP(16'h149D7,4);
TASK_PP(16'h149D8,4);
TASK_PP(16'h149D9,4);
TASK_PP(16'h149DA,4);
TASK_PP(16'h149DB,4);
TASK_PP(16'h149DC,4);
TASK_PP(16'h149DD,4);
TASK_PP(16'h149DE,4);
TASK_PP(16'h149DF,4);
TASK_PP(16'h149E0,4);
TASK_PP(16'h149E1,4);
TASK_PP(16'h149E2,4);
TASK_PP(16'h149E3,4);
TASK_PP(16'h149E4,4);
TASK_PP(16'h149E5,4);
TASK_PP(16'h149E6,4);
TASK_PP(16'h149E7,4);
TASK_PP(16'h149E8,4);
TASK_PP(16'h149E9,4);
TASK_PP(16'h149EA,4);
TASK_PP(16'h149EB,4);
TASK_PP(16'h149EC,4);
TASK_PP(16'h149ED,4);
TASK_PP(16'h149EE,4);
TASK_PP(16'h149EF,4);
TASK_PP(16'h149F0,4);
TASK_PP(16'h149F1,4);
TASK_PP(16'h149F2,4);
TASK_PP(16'h149F3,4);
TASK_PP(16'h149F4,4);
TASK_PP(16'h149F5,4);
TASK_PP(16'h149F6,4);
TASK_PP(16'h149F7,4);
TASK_PP(16'h149F8,4);
TASK_PP(16'h149F9,4);
TASK_PP(16'h149FA,4);
TASK_PP(16'h149FB,4);
TASK_PP(16'h149FC,4);
TASK_PP(16'h149FD,4);
TASK_PP(16'h149FE,4);
TASK_PP(16'h149FF,4);
TASK_PP(16'h14A00,4);
TASK_PP(16'h14A01,4);
TASK_PP(16'h14A02,4);
TASK_PP(16'h14A03,4);
TASK_PP(16'h14A04,4);
TASK_PP(16'h14A05,4);
TASK_PP(16'h14A06,4);
TASK_PP(16'h14A07,4);
TASK_PP(16'h14A08,4);
TASK_PP(16'h14A09,4);
TASK_PP(16'h14A0A,4);
TASK_PP(16'h14A0B,4);
TASK_PP(16'h14A0C,4);
TASK_PP(16'h14A0D,4);
TASK_PP(16'h14A0E,4);
TASK_PP(16'h14A0F,4);
TASK_PP(16'h14A10,4);
TASK_PP(16'h14A11,4);
TASK_PP(16'h14A12,4);
TASK_PP(16'h14A13,4);
TASK_PP(16'h14A14,4);
TASK_PP(16'h14A15,4);
TASK_PP(16'h14A16,4);
TASK_PP(16'h14A17,4);
TASK_PP(16'h14A18,4);
TASK_PP(16'h14A19,4);
TASK_PP(16'h14A1A,4);
TASK_PP(16'h14A1B,4);
TASK_PP(16'h14A1C,4);
TASK_PP(16'h14A1D,4);
TASK_PP(16'h14A1E,4);
TASK_PP(16'h14A1F,4);
TASK_PP(16'h14A20,4);
TASK_PP(16'h14A21,4);
TASK_PP(16'h14A22,4);
TASK_PP(16'h14A23,4);
TASK_PP(16'h14A24,4);
TASK_PP(16'h14A25,4);
TASK_PP(16'h14A26,4);
TASK_PP(16'h14A27,4);
TASK_PP(16'h14A28,4);
TASK_PP(16'h14A29,4);
TASK_PP(16'h14A2A,4);
TASK_PP(16'h14A2B,4);
TASK_PP(16'h14A2C,4);
TASK_PP(16'h14A2D,4);
TASK_PP(16'h14A2E,4);
TASK_PP(16'h14A2F,4);
TASK_PP(16'h14A30,4);
TASK_PP(16'h14A31,4);
TASK_PP(16'h14A32,4);
TASK_PP(16'h14A33,4);
TASK_PP(16'h14A34,4);
TASK_PP(16'h14A35,4);
TASK_PP(16'h14A36,4);
TASK_PP(16'h14A37,4);
TASK_PP(16'h14A38,4);
TASK_PP(16'h14A39,4);
TASK_PP(16'h14A3A,4);
TASK_PP(16'h14A3B,4);
TASK_PP(16'h14A3C,4);
TASK_PP(16'h14A3D,4);
TASK_PP(16'h14A3E,4);
TASK_PP(16'h14A3F,4);
TASK_PP(16'h14A40,4);
TASK_PP(16'h14A41,4);
TASK_PP(16'h14A42,4);
TASK_PP(16'h14A43,4);
TASK_PP(16'h14A44,4);
TASK_PP(16'h14A45,4);
TASK_PP(16'h14A46,4);
TASK_PP(16'h14A47,4);
TASK_PP(16'h14A48,4);
TASK_PP(16'h14A49,4);
TASK_PP(16'h14A4A,4);
TASK_PP(16'h14A4B,4);
TASK_PP(16'h14A4C,4);
TASK_PP(16'h14A4D,4);
TASK_PP(16'h14A4E,4);
TASK_PP(16'h14A4F,4);
TASK_PP(16'h14A50,4);
TASK_PP(16'h14A51,4);
TASK_PP(16'h14A52,4);
TASK_PP(16'h14A53,4);
TASK_PP(16'h14A54,4);
TASK_PP(16'h14A55,4);
TASK_PP(16'h14A56,4);
TASK_PP(16'h14A57,4);
TASK_PP(16'h14A58,4);
TASK_PP(16'h14A59,4);
TASK_PP(16'h14A5A,4);
TASK_PP(16'h14A5B,4);
TASK_PP(16'h14A5C,4);
TASK_PP(16'h14A5D,4);
TASK_PP(16'h14A5E,4);
TASK_PP(16'h14A5F,4);
TASK_PP(16'h14A60,4);
TASK_PP(16'h14A61,4);
TASK_PP(16'h14A62,4);
TASK_PP(16'h14A63,4);
TASK_PP(16'h14A64,4);
TASK_PP(16'h14A65,4);
TASK_PP(16'h14A66,4);
TASK_PP(16'h14A67,4);
TASK_PP(16'h14A68,4);
TASK_PP(16'h14A69,4);
TASK_PP(16'h14A6A,4);
TASK_PP(16'h14A6B,4);
TASK_PP(16'h14A6C,4);
TASK_PP(16'h14A6D,4);
TASK_PP(16'h14A6E,4);
TASK_PP(16'h14A6F,4);
TASK_PP(16'h14A70,4);
TASK_PP(16'h14A71,4);
TASK_PP(16'h14A72,4);
TASK_PP(16'h14A73,4);
TASK_PP(16'h14A74,4);
TASK_PP(16'h14A75,4);
TASK_PP(16'h14A76,4);
TASK_PP(16'h14A77,4);
TASK_PP(16'h14A78,4);
TASK_PP(16'h14A79,4);
TASK_PP(16'h14A7A,4);
TASK_PP(16'h14A7B,4);
TASK_PP(16'h14A7C,4);
TASK_PP(16'h14A7D,4);
TASK_PP(16'h14A7E,4);
TASK_PP(16'h14A7F,4);
TASK_PP(16'h14A80,4);
TASK_PP(16'h14A81,4);
TASK_PP(16'h14A82,4);
TASK_PP(16'h14A83,4);
TASK_PP(16'h14A84,4);
TASK_PP(16'h14A85,4);
TASK_PP(16'h14A86,4);
TASK_PP(16'h14A87,4);
TASK_PP(16'h14A88,4);
TASK_PP(16'h14A89,4);
TASK_PP(16'h14A8A,4);
TASK_PP(16'h14A8B,4);
TASK_PP(16'h14A8C,4);
TASK_PP(16'h14A8D,4);
TASK_PP(16'h14A8E,4);
TASK_PP(16'h14A8F,4);
TASK_PP(16'h14A90,4);
TASK_PP(16'h14A91,4);
TASK_PP(16'h14A92,4);
TASK_PP(16'h14A93,4);
TASK_PP(16'h14A94,4);
TASK_PP(16'h14A95,4);
TASK_PP(16'h14A96,4);
TASK_PP(16'h14A97,4);
TASK_PP(16'h14A98,4);
TASK_PP(16'h14A99,4);
TASK_PP(16'h14A9A,4);
TASK_PP(16'h14A9B,4);
TASK_PP(16'h14A9C,4);
TASK_PP(16'h14A9D,4);
TASK_PP(16'h14A9E,4);
TASK_PP(16'h14A9F,4);
TASK_PP(16'h14AA0,4);
TASK_PP(16'h14AA1,4);
TASK_PP(16'h14AA2,4);
TASK_PP(16'h14AA3,4);
TASK_PP(16'h14AA4,4);
TASK_PP(16'h14AA5,4);
TASK_PP(16'h14AA6,4);
TASK_PP(16'h14AA7,4);
TASK_PP(16'h14AA8,4);
TASK_PP(16'h14AA9,4);
TASK_PP(16'h14AAA,4);
TASK_PP(16'h14AAB,4);
TASK_PP(16'h14AAC,4);
TASK_PP(16'h14AAD,4);
TASK_PP(16'h14AAE,4);
TASK_PP(16'h14AAF,4);
TASK_PP(16'h14AB0,4);
TASK_PP(16'h14AB1,4);
TASK_PP(16'h14AB2,4);
TASK_PP(16'h14AB3,4);
TASK_PP(16'h14AB4,4);
TASK_PP(16'h14AB5,4);
TASK_PP(16'h14AB6,4);
TASK_PP(16'h14AB7,4);
TASK_PP(16'h14AB8,4);
TASK_PP(16'h14AB9,4);
TASK_PP(16'h14ABA,4);
TASK_PP(16'h14ABB,4);
TASK_PP(16'h14ABC,4);
TASK_PP(16'h14ABD,4);
TASK_PP(16'h14ABE,4);
TASK_PP(16'h14ABF,4);
TASK_PP(16'h14AC0,4);
TASK_PP(16'h14AC1,4);
TASK_PP(16'h14AC2,4);
TASK_PP(16'h14AC3,4);
TASK_PP(16'h14AC4,4);
TASK_PP(16'h14AC5,4);
TASK_PP(16'h14AC6,4);
TASK_PP(16'h14AC7,4);
TASK_PP(16'h14AC8,4);
TASK_PP(16'h14AC9,4);
TASK_PP(16'h14ACA,4);
TASK_PP(16'h14ACB,4);
TASK_PP(16'h14ACC,4);
TASK_PP(16'h14ACD,4);
TASK_PP(16'h14ACE,4);
TASK_PP(16'h14ACF,4);
TASK_PP(16'h14AD0,4);
TASK_PP(16'h14AD1,4);
TASK_PP(16'h14AD2,4);
TASK_PP(16'h14AD3,4);
TASK_PP(16'h14AD4,4);
TASK_PP(16'h14AD5,4);
TASK_PP(16'h14AD6,4);
TASK_PP(16'h14AD7,4);
TASK_PP(16'h14AD8,4);
TASK_PP(16'h14AD9,4);
TASK_PP(16'h14ADA,4);
TASK_PP(16'h14ADB,4);
TASK_PP(16'h14ADC,4);
TASK_PP(16'h14ADD,4);
TASK_PP(16'h14ADE,4);
TASK_PP(16'h14ADF,4);
TASK_PP(16'h14AE0,4);
TASK_PP(16'h14AE1,4);
TASK_PP(16'h14AE2,4);
TASK_PP(16'h14AE3,4);
TASK_PP(16'h14AE4,4);
TASK_PP(16'h14AE5,4);
TASK_PP(16'h14AE6,4);
TASK_PP(16'h14AE7,4);
TASK_PP(16'h14AE8,4);
TASK_PP(16'h14AE9,4);
TASK_PP(16'h14AEA,4);
TASK_PP(16'h14AEB,4);
TASK_PP(16'h14AEC,4);
TASK_PP(16'h14AED,4);
TASK_PP(16'h14AEE,4);
TASK_PP(16'h14AEF,4);
TASK_PP(16'h14AF0,4);
TASK_PP(16'h14AF1,4);
TASK_PP(16'h14AF2,4);
TASK_PP(16'h14AF3,4);
TASK_PP(16'h14AF4,4);
TASK_PP(16'h14AF5,4);
TASK_PP(16'h14AF6,4);
TASK_PP(16'h14AF7,4);
TASK_PP(16'h14AF8,4);
TASK_PP(16'h14AF9,4);
TASK_PP(16'h14AFA,4);
TASK_PP(16'h14AFB,4);
TASK_PP(16'h14AFC,4);
TASK_PP(16'h14AFD,4);
TASK_PP(16'h14AFE,4);
TASK_PP(16'h14AFF,4);
TASK_PP(16'h14B00,4);
TASK_PP(16'h14B01,4);
TASK_PP(16'h14B02,4);
TASK_PP(16'h14B03,4);
TASK_PP(16'h14B04,4);
TASK_PP(16'h14B05,4);
TASK_PP(16'h14B06,4);
TASK_PP(16'h14B07,4);
TASK_PP(16'h14B08,4);
TASK_PP(16'h14B09,4);
TASK_PP(16'h14B0A,4);
TASK_PP(16'h14B0B,4);
TASK_PP(16'h14B0C,4);
TASK_PP(16'h14B0D,4);
TASK_PP(16'h14B0E,4);
TASK_PP(16'h14B0F,4);
TASK_PP(16'h14B10,4);
TASK_PP(16'h14B11,4);
TASK_PP(16'h14B12,4);
TASK_PP(16'h14B13,4);
TASK_PP(16'h14B14,4);
TASK_PP(16'h14B15,4);
TASK_PP(16'h14B16,4);
TASK_PP(16'h14B17,4);
TASK_PP(16'h14B18,4);
TASK_PP(16'h14B19,4);
TASK_PP(16'h14B1A,4);
TASK_PP(16'h14B1B,4);
TASK_PP(16'h14B1C,4);
TASK_PP(16'h14B1D,4);
TASK_PP(16'h14B1E,4);
TASK_PP(16'h14B1F,4);
TASK_PP(16'h14B20,4);
TASK_PP(16'h14B21,4);
TASK_PP(16'h14B22,4);
TASK_PP(16'h14B23,4);
TASK_PP(16'h14B24,4);
TASK_PP(16'h14B25,4);
TASK_PP(16'h14B26,4);
TASK_PP(16'h14B27,4);
TASK_PP(16'h14B28,4);
TASK_PP(16'h14B29,4);
TASK_PP(16'h14B2A,4);
TASK_PP(16'h14B2B,4);
TASK_PP(16'h14B2C,4);
TASK_PP(16'h14B2D,4);
TASK_PP(16'h14B2E,4);
TASK_PP(16'h14B2F,4);
TASK_PP(16'h14B30,4);
TASK_PP(16'h14B31,4);
TASK_PP(16'h14B32,4);
TASK_PP(16'h14B33,4);
TASK_PP(16'h14B34,4);
TASK_PP(16'h14B35,4);
TASK_PP(16'h14B36,4);
TASK_PP(16'h14B37,4);
TASK_PP(16'h14B38,4);
TASK_PP(16'h14B39,4);
TASK_PP(16'h14B3A,4);
TASK_PP(16'h14B3B,4);
TASK_PP(16'h14B3C,4);
TASK_PP(16'h14B3D,4);
TASK_PP(16'h14B3E,4);
TASK_PP(16'h14B3F,4);
TASK_PP(16'h14B40,4);
TASK_PP(16'h14B41,4);
TASK_PP(16'h14B42,4);
TASK_PP(16'h14B43,4);
TASK_PP(16'h14B44,4);
TASK_PP(16'h14B45,4);
TASK_PP(16'h14B46,4);
TASK_PP(16'h14B47,4);
TASK_PP(16'h14B48,4);
TASK_PP(16'h14B49,4);
TASK_PP(16'h14B4A,4);
TASK_PP(16'h14B4B,4);
TASK_PP(16'h14B4C,4);
TASK_PP(16'h14B4D,4);
TASK_PP(16'h14B4E,4);
TASK_PP(16'h14B4F,4);
TASK_PP(16'h14B50,4);
TASK_PP(16'h14B51,4);
TASK_PP(16'h14B52,4);
TASK_PP(16'h14B53,4);
TASK_PP(16'h14B54,4);
TASK_PP(16'h14B55,4);
TASK_PP(16'h14B56,4);
TASK_PP(16'h14B57,4);
TASK_PP(16'h14B58,4);
TASK_PP(16'h14B59,4);
TASK_PP(16'h14B5A,4);
TASK_PP(16'h14B5B,4);
TASK_PP(16'h14B5C,4);
TASK_PP(16'h14B5D,4);
TASK_PP(16'h14B5E,4);
TASK_PP(16'h14B5F,4);
TASK_PP(16'h14B60,4);
TASK_PP(16'h14B61,4);
TASK_PP(16'h14B62,4);
TASK_PP(16'h14B63,4);
TASK_PP(16'h14B64,4);
TASK_PP(16'h14B65,4);
TASK_PP(16'h14B66,4);
TASK_PP(16'h14B67,4);
TASK_PP(16'h14B68,4);
TASK_PP(16'h14B69,4);
TASK_PP(16'h14B6A,4);
TASK_PP(16'h14B6B,4);
TASK_PP(16'h14B6C,4);
TASK_PP(16'h14B6D,4);
TASK_PP(16'h14B6E,4);
TASK_PP(16'h14B6F,4);
TASK_PP(16'h14B70,4);
TASK_PP(16'h14B71,4);
TASK_PP(16'h14B72,4);
TASK_PP(16'h14B73,4);
TASK_PP(16'h14B74,4);
TASK_PP(16'h14B75,4);
TASK_PP(16'h14B76,4);
TASK_PP(16'h14B77,4);
TASK_PP(16'h14B78,4);
TASK_PP(16'h14B79,4);
TASK_PP(16'h14B7A,4);
TASK_PP(16'h14B7B,4);
TASK_PP(16'h14B7C,4);
TASK_PP(16'h14B7D,4);
TASK_PP(16'h14B7E,4);
TASK_PP(16'h14B7F,4);
TASK_PP(16'h14B80,4);
TASK_PP(16'h14B81,4);
TASK_PP(16'h14B82,4);
TASK_PP(16'h14B83,4);
TASK_PP(16'h14B84,4);
TASK_PP(16'h14B85,4);
TASK_PP(16'h14B86,4);
TASK_PP(16'h14B87,4);
TASK_PP(16'h14B88,4);
TASK_PP(16'h14B89,4);
TASK_PP(16'h14B8A,4);
TASK_PP(16'h14B8B,4);
TASK_PP(16'h14B8C,4);
TASK_PP(16'h14B8D,4);
TASK_PP(16'h14B8E,4);
TASK_PP(16'h14B8F,4);
TASK_PP(16'h14B90,4);
TASK_PP(16'h14B91,4);
TASK_PP(16'h14B92,4);
TASK_PP(16'h14B93,4);
TASK_PP(16'h14B94,4);
TASK_PP(16'h14B95,4);
TASK_PP(16'h14B96,4);
TASK_PP(16'h14B97,4);
TASK_PP(16'h14B98,4);
TASK_PP(16'h14B99,4);
TASK_PP(16'h14B9A,4);
TASK_PP(16'h14B9B,4);
TASK_PP(16'h14B9C,4);
TASK_PP(16'h14B9D,4);
TASK_PP(16'h14B9E,4);
TASK_PP(16'h14B9F,4);
TASK_PP(16'h14BA0,4);
TASK_PP(16'h14BA1,4);
TASK_PP(16'h14BA2,4);
TASK_PP(16'h14BA3,4);
TASK_PP(16'h14BA4,4);
TASK_PP(16'h14BA5,4);
TASK_PP(16'h14BA6,4);
TASK_PP(16'h14BA7,4);
TASK_PP(16'h14BA8,4);
TASK_PP(16'h14BA9,4);
TASK_PP(16'h14BAA,4);
TASK_PP(16'h14BAB,4);
TASK_PP(16'h14BAC,4);
TASK_PP(16'h14BAD,4);
TASK_PP(16'h14BAE,4);
TASK_PP(16'h14BAF,4);
TASK_PP(16'h14BB0,4);
TASK_PP(16'h14BB1,4);
TASK_PP(16'h14BB2,4);
TASK_PP(16'h14BB3,4);
TASK_PP(16'h14BB4,4);
TASK_PP(16'h14BB5,4);
TASK_PP(16'h14BB6,4);
TASK_PP(16'h14BB7,4);
TASK_PP(16'h14BB8,4);
TASK_PP(16'h14BB9,4);
TASK_PP(16'h14BBA,4);
TASK_PP(16'h14BBB,4);
TASK_PP(16'h14BBC,4);
TASK_PP(16'h14BBD,4);
TASK_PP(16'h14BBE,4);
TASK_PP(16'h14BBF,4);
TASK_PP(16'h14BC0,4);
TASK_PP(16'h14BC1,4);
TASK_PP(16'h14BC2,4);
TASK_PP(16'h14BC3,4);
TASK_PP(16'h14BC4,4);
TASK_PP(16'h14BC5,4);
TASK_PP(16'h14BC6,4);
TASK_PP(16'h14BC7,4);
TASK_PP(16'h14BC8,4);
TASK_PP(16'h14BC9,4);
TASK_PP(16'h14BCA,4);
TASK_PP(16'h14BCB,4);
TASK_PP(16'h14BCC,4);
TASK_PP(16'h14BCD,4);
TASK_PP(16'h14BCE,4);
TASK_PP(16'h14BCF,4);
TASK_PP(16'h14BD0,4);
TASK_PP(16'h14BD1,4);
TASK_PP(16'h14BD2,4);
TASK_PP(16'h14BD3,4);
TASK_PP(16'h14BD4,4);
TASK_PP(16'h14BD5,4);
TASK_PP(16'h14BD6,4);
TASK_PP(16'h14BD7,4);
TASK_PP(16'h14BD8,4);
TASK_PP(16'h14BD9,4);
TASK_PP(16'h14BDA,4);
TASK_PP(16'h14BDB,4);
TASK_PP(16'h14BDC,4);
TASK_PP(16'h14BDD,4);
TASK_PP(16'h14BDE,4);
TASK_PP(16'h14BDF,4);
TASK_PP(16'h14BE0,4);
TASK_PP(16'h14BE1,4);
TASK_PP(16'h14BE2,4);
TASK_PP(16'h14BE3,4);
TASK_PP(16'h14BE4,4);
TASK_PP(16'h14BE5,4);
TASK_PP(16'h14BE6,4);
TASK_PP(16'h14BE7,4);
TASK_PP(16'h14BE8,4);
TASK_PP(16'h14BE9,4);
TASK_PP(16'h14BEA,4);
TASK_PP(16'h14BEB,4);
TASK_PP(16'h14BEC,4);
TASK_PP(16'h14BED,4);
TASK_PP(16'h14BEE,4);
TASK_PP(16'h14BEF,4);
TASK_PP(16'h14BF0,4);
TASK_PP(16'h14BF1,4);
TASK_PP(16'h14BF2,4);
TASK_PP(16'h14BF3,4);
TASK_PP(16'h14BF4,4);
TASK_PP(16'h14BF5,4);
TASK_PP(16'h14BF6,4);
TASK_PP(16'h14BF7,4);
TASK_PP(16'h14BF8,4);
TASK_PP(16'h14BF9,4);
TASK_PP(16'h14BFA,4);
TASK_PP(16'h14BFB,4);
TASK_PP(16'h14BFC,4);
TASK_PP(16'h14BFD,4);
TASK_PP(16'h14BFE,4);
TASK_PP(16'h14BFF,4);
TASK_PP(16'h14C00,4);
TASK_PP(16'h14C01,4);
TASK_PP(16'h14C02,4);
TASK_PP(16'h14C03,4);
TASK_PP(16'h14C04,4);
TASK_PP(16'h14C05,4);
TASK_PP(16'h14C06,4);
TASK_PP(16'h14C07,4);
TASK_PP(16'h14C08,4);
TASK_PP(16'h14C09,4);
TASK_PP(16'h14C0A,4);
TASK_PP(16'h14C0B,4);
TASK_PP(16'h14C0C,4);
TASK_PP(16'h14C0D,4);
TASK_PP(16'h14C0E,4);
TASK_PP(16'h14C0F,4);
TASK_PP(16'h14C10,4);
TASK_PP(16'h14C11,4);
TASK_PP(16'h14C12,4);
TASK_PP(16'h14C13,4);
TASK_PP(16'h14C14,4);
TASK_PP(16'h14C15,4);
TASK_PP(16'h14C16,4);
TASK_PP(16'h14C17,4);
TASK_PP(16'h14C18,4);
TASK_PP(16'h14C19,4);
TASK_PP(16'h14C1A,4);
TASK_PP(16'h14C1B,4);
TASK_PP(16'h14C1C,4);
TASK_PP(16'h14C1D,4);
TASK_PP(16'h14C1E,4);
TASK_PP(16'h14C1F,4);
TASK_PP(16'h14C20,4);
TASK_PP(16'h14C21,4);
TASK_PP(16'h14C22,4);
TASK_PP(16'h14C23,4);
TASK_PP(16'h14C24,4);
TASK_PP(16'h14C25,4);
TASK_PP(16'h14C26,4);
TASK_PP(16'h14C27,4);
TASK_PP(16'h14C28,4);
TASK_PP(16'h14C29,4);
TASK_PP(16'h14C2A,4);
TASK_PP(16'h14C2B,4);
TASK_PP(16'h14C2C,4);
TASK_PP(16'h14C2D,4);
TASK_PP(16'h14C2E,4);
TASK_PP(16'h14C2F,4);
TASK_PP(16'h14C30,4);
TASK_PP(16'h14C31,4);
TASK_PP(16'h14C32,4);
TASK_PP(16'h14C33,4);
TASK_PP(16'h14C34,4);
TASK_PP(16'h14C35,4);
TASK_PP(16'h14C36,4);
TASK_PP(16'h14C37,4);
TASK_PP(16'h14C38,4);
TASK_PP(16'h14C39,4);
TASK_PP(16'h14C3A,4);
TASK_PP(16'h14C3B,4);
TASK_PP(16'h14C3C,4);
TASK_PP(16'h14C3D,4);
TASK_PP(16'h14C3E,4);
TASK_PP(16'h14C3F,4);
TASK_PP(16'h14C40,4);
TASK_PP(16'h14C41,4);
TASK_PP(16'h14C42,4);
TASK_PP(16'h14C43,4);
TASK_PP(16'h14C44,4);
TASK_PP(16'h14C45,4);
TASK_PP(16'h14C46,4);
TASK_PP(16'h14C47,4);
TASK_PP(16'h14C48,4);
TASK_PP(16'h14C49,4);
TASK_PP(16'h14C4A,4);
TASK_PP(16'h14C4B,4);
TASK_PP(16'h14C4C,4);
TASK_PP(16'h14C4D,4);
TASK_PP(16'h14C4E,4);
TASK_PP(16'h14C4F,4);
TASK_PP(16'h14C50,4);
TASK_PP(16'h14C51,4);
TASK_PP(16'h14C52,4);
TASK_PP(16'h14C53,4);
TASK_PP(16'h14C54,4);
TASK_PP(16'h14C55,4);
TASK_PP(16'h14C56,4);
TASK_PP(16'h14C57,4);
TASK_PP(16'h14C58,4);
TASK_PP(16'h14C59,4);
TASK_PP(16'h14C5A,4);
TASK_PP(16'h14C5B,4);
TASK_PP(16'h14C5C,4);
TASK_PP(16'h14C5D,4);
TASK_PP(16'h14C5E,4);
TASK_PP(16'h14C5F,4);
TASK_PP(16'h14C60,4);
TASK_PP(16'h14C61,4);
TASK_PP(16'h14C62,4);
TASK_PP(16'h14C63,4);
TASK_PP(16'h14C64,4);
TASK_PP(16'h14C65,4);
TASK_PP(16'h14C66,4);
TASK_PP(16'h14C67,4);
TASK_PP(16'h14C68,4);
TASK_PP(16'h14C69,4);
TASK_PP(16'h14C6A,4);
TASK_PP(16'h14C6B,4);
TASK_PP(16'h14C6C,4);
TASK_PP(16'h14C6D,4);
TASK_PP(16'h14C6E,4);
TASK_PP(16'h14C6F,4);
TASK_PP(16'h14C70,4);
TASK_PP(16'h14C71,4);
TASK_PP(16'h14C72,4);
TASK_PP(16'h14C73,4);
TASK_PP(16'h14C74,4);
TASK_PP(16'h14C75,4);
TASK_PP(16'h14C76,4);
TASK_PP(16'h14C77,4);
TASK_PP(16'h14C78,4);
TASK_PP(16'h14C79,4);
TASK_PP(16'h14C7A,4);
TASK_PP(16'h14C7B,4);
TASK_PP(16'h14C7C,4);
TASK_PP(16'h14C7D,4);
TASK_PP(16'h14C7E,4);
TASK_PP(16'h14C7F,4);
TASK_PP(16'h14C80,4);
TASK_PP(16'h14C81,4);
TASK_PP(16'h14C82,4);
TASK_PP(16'h14C83,4);
TASK_PP(16'h14C84,4);
TASK_PP(16'h14C85,4);
TASK_PP(16'h14C86,4);
TASK_PP(16'h14C87,4);
TASK_PP(16'h14C88,4);
TASK_PP(16'h14C89,4);
TASK_PP(16'h14C8A,4);
TASK_PP(16'h14C8B,4);
TASK_PP(16'h14C8C,4);
TASK_PP(16'h14C8D,4);
TASK_PP(16'h14C8E,4);
TASK_PP(16'h14C8F,4);
TASK_PP(16'h14C90,4);
TASK_PP(16'h14C91,4);
TASK_PP(16'h14C92,4);
TASK_PP(16'h14C93,4);
TASK_PP(16'h14C94,4);
TASK_PP(16'h14C95,4);
TASK_PP(16'h14C96,4);
TASK_PP(16'h14C97,4);
TASK_PP(16'h14C98,4);
TASK_PP(16'h14C99,4);
TASK_PP(16'h14C9A,4);
TASK_PP(16'h14C9B,4);
TASK_PP(16'h14C9C,4);
TASK_PP(16'h14C9D,4);
TASK_PP(16'h14C9E,4);
TASK_PP(16'h14C9F,4);
TASK_PP(16'h14CA0,4);
TASK_PP(16'h14CA1,4);
TASK_PP(16'h14CA2,4);
TASK_PP(16'h14CA3,4);
TASK_PP(16'h14CA4,4);
TASK_PP(16'h14CA5,4);
TASK_PP(16'h14CA6,4);
TASK_PP(16'h14CA7,4);
TASK_PP(16'h14CA8,4);
TASK_PP(16'h14CA9,4);
TASK_PP(16'h14CAA,4);
TASK_PP(16'h14CAB,4);
TASK_PP(16'h14CAC,4);
TASK_PP(16'h14CAD,4);
TASK_PP(16'h14CAE,4);
TASK_PP(16'h14CAF,4);
TASK_PP(16'h14CB0,4);
TASK_PP(16'h14CB1,4);
TASK_PP(16'h14CB2,4);
TASK_PP(16'h14CB3,4);
TASK_PP(16'h14CB4,4);
TASK_PP(16'h14CB5,4);
TASK_PP(16'h14CB6,4);
TASK_PP(16'h14CB7,4);
TASK_PP(16'h14CB8,4);
TASK_PP(16'h14CB9,4);
TASK_PP(16'h14CBA,4);
TASK_PP(16'h14CBB,4);
TASK_PP(16'h14CBC,4);
TASK_PP(16'h14CBD,4);
TASK_PP(16'h14CBE,4);
TASK_PP(16'h14CBF,4);
TASK_PP(16'h14CC0,4);
TASK_PP(16'h14CC1,4);
TASK_PP(16'h14CC2,4);
TASK_PP(16'h14CC3,4);
TASK_PP(16'h14CC4,4);
TASK_PP(16'h14CC5,4);
TASK_PP(16'h14CC6,4);
TASK_PP(16'h14CC7,4);
TASK_PP(16'h14CC8,4);
TASK_PP(16'h14CC9,4);
TASK_PP(16'h14CCA,4);
TASK_PP(16'h14CCB,4);
TASK_PP(16'h14CCC,4);
TASK_PP(16'h14CCD,4);
TASK_PP(16'h14CCE,4);
TASK_PP(16'h14CCF,4);
TASK_PP(16'h14CD0,4);
TASK_PP(16'h14CD1,4);
TASK_PP(16'h14CD2,4);
TASK_PP(16'h14CD3,4);
TASK_PP(16'h14CD4,4);
TASK_PP(16'h14CD5,4);
TASK_PP(16'h14CD6,4);
TASK_PP(16'h14CD7,4);
TASK_PP(16'h14CD8,4);
TASK_PP(16'h14CD9,4);
TASK_PP(16'h14CDA,4);
TASK_PP(16'h14CDB,4);
TASK_PP(16'h14CDC,4);
TASK_PP(16'h14CDD,4);
TASK_PP(16'h14CDE,4);
TASK_PP(16'h14CDF,4);
TASK_PP(16'h14CE0,4);
TASK_PP(16'h14CE1,4);
TASK_PP(16'h14CE2,4);
TASK_PP(16'h14CE3,4);
TASK_PP(16'h14CE4,4);
TASK_PP(16'h14CE5,4);
TASK_PP(16'h14CE6,4);
TASK_PP(16'h14CE7,4);
TASK_PP(16'h14CE8,4);
TASK_PP(16'h14CE9,4);
TASK_PP(16'h14CEA,4);
TASK_PP(16'h14CEB,4);
TASK_PP(16'h14CEC,4);
TASK_PP(16'h14CED,4);
TASK_PP(16'h14CEE,4);
TASK_PP(16'h14CEF,4);
TASK_PP(16'h14CF0,4);
TASK_PP(16'h14CF1,4);
TASK_PP(16'h14CF2,4);
TASK_PP(16'h14CF3,4);
TASK_PP(16'h14CF4,4);
TASK_PP(16'h14CF5,4);
TASK_PP(16'h14CF6,4);
TASK_PP(16'h14CF7,4);
TASK_PP(16'h14CF8,4);
TASK_PP(16'h14CF9,4);
TASK_PP(16'h14CFA,4);
TASK_PP(16'h14CFB,4);
TASK_PP(16'h14CFC,4);
TASK_PP(16'h14CFD,4);
TASK_PP(16'h14CFE,4);
TASK_PP(16'h14CFF,4);
TASK_PP(16'h14D00,4);
TASK_PP(16'h14D01,4);
TASK_PP(16'h14D02,4);
TASK_PP(16'h14D03,4);
TASK_PP(16'h14D04,4);
TASK_PP(16'h14D05,4);
TASK_PP(16'h14D06,4);
TASK_PP(16'h14D07,4);
TASK_PP(16'h14D08,4);
TASK_PP(16'h14D09,4);
TASK_PP(16'h14D0A,4);
TASK_PP(16'h14D0B,4);
TASK_PP(16'h14D0C,4);
TASK_PP(16'h14D0D,4);
TASK_PP(16'h14D0E,4);
TASK_PP(16'h14D0F,4);
TASK_PP(16'h14D10,4);
TASK_PP(16'h14D11,4);
TASK_PP(16'h14D12,4);
TASK_PP(16'h14D13,4);
TASK_PP(16'h14D14,4);
TASK_PP(16'h14D15,4);
TASK_PP(16'h14D16,4);
TASK_PP(16'h14D17,4);
TASK_PP(16'h14D18,4);
TASK_PP(16'h14D19,4);
TASK_PP(16'h14D1A,4);
TASK_PP(16'h14D1B,4);
TASK_PP(16'h14D1C,4);
TASK_PP(16'h14D1D,4);
TASK_PP(16'h14D1E,4);
TASK_PP(16'h14D1F,4);
TASK_PP(16'h14D20,4);
TASK_PP(16'h14D21,4);
TASK_PP(16'h14D22,4);
TASK_PP(16'h14D23,4);
TASK_PP(16'h14D24,4);
TASK_PP(16'h14D25,4);
TASK_PP(16'h14D26,4);
TASK_PP(16'h14D27,4);
TASK_PP(16'h14D28,4);
TASK_PP(16'h14D29,4);
TASK_PP(16'h14D2A,4);
TASK_PP(16'h14D2B,4);
TASK_PP(16'h14D2C,4);
TASK_PP(16'h14D2D,4);
TASK_PP(16'h14D2E,4);
TASK_PP(16'h14D2F,4);
TASK_PP(16'h14D30,4);
TASK_PP(16'h14D31,4);
TASK_PP(16'h14D32,4);
TASK_PP(16'h14D33,4);
TASK_PP(16'h14D34,4);
TASK_PP(16'h14D35,4);
TASK_PP(16'h14D36,4);
TASK_PP(16'h14D37,4);
TASK_PP(16'h14D38,4);
TASK_PP(16'h14D39,4);
TASK_PP(16'h14D3A,4);
TASK_PP(16'h14D3B,4);
TASK_PP(16'h14D3C,4);
TASK_PP(16'h14D3D,4);
TASK_PP(16'h14D3E,4);
TASK_PP(16'h14D3F,4);
TASK_PP(16'h14D40,4);
TASK_PP(16'h14D41,4);
TASK_PP(16'h14D42,4);
TASK_PP(16'h14D43,4);
TASK_PP(16'h14D44,4);
TASK_PP(16'h14D45,4);
TASK_PP(16'h14D46,4);
TASK_PP(16'h14D47,4);
TASK_PP(16'h14D48,4);
TASK_PP(16'h14D49,4);
TASK_PP(16'h14D4A,4);
TASK_PP(16'h14D4B,4);
TASK_PP(16'h14D4C,4);
TASK_PP(16'h14D4D,4);
TASK_PP(16'h14D4E,4);
TASK_PP(16'h14D4F,4);
TASK_PP(16'h14D50,4);
TASK_PP(16'h14D51,4);
TASK_PP(16'h14D52,4);
TASK_PP(16'h14D53,4);
TASK_PP(16'h14D54,4);
TASK_PP(16'h14D55,4);
TASK_PP(16'h14D56,4);
TASK_PP(16'h14D57,4);
TASK_PP(16'h14D58,4);
TASK_PP(16'h14D59,4);
TASK_PP(16'h14D5A,4);
TASK_PP(16'h14D5B,4);
TASK_PP(16'h14D5C,4);
TASK_PP(16'h14D5D,4);
TASK_PP(16'h14D5E,4);
TASK_PP(16'h14D5F,4);
TASK_PP(16'h14D60,4);
TASK_PP(16'h14D61,4);
TASK_PP(16'h14D62,4);
TASK_PP(16'h14D63,4);
TASK_PP(16'h14D64,4);
TASK_PP(16'h14D65,4);
TASK_PP(16'h14D66,4);
TASK_PP(16'h14D67,4);
TASK_PP(16'h14D68,4);
TASK_PP(16'h14D69,4);
TASK_PP(16'h14D6A,4);
TASK_PP(16'h14D6B,4);
TASK_PP(16'h14D6C,4);
TASK_PP(16'h14D6D,4);
TASK_PP(16'h14D6E,4);
TASK_PP(16'h14D6F,4);
TASK_PP(16'h14D70,4);
TASK_PP(16'h14D71,4);
TASK_PP(16'h14D72,4);
TASK_PP(16'h14D73,4);
TASK_PP(16'h14D74,4);
TASK_PP(16'h14D75,4);
TASK_PP(16'h14D76,4);
TASK_PP(16'h14D77,4);
TASK_PP(16'h14D78,4);
TASK_PP(16'h14D79,4);
TASK_PP(16'h14D7A,4);
TASK_PP(16'h14D7B,4);
TASK_PP(16'h14D7C,4);
TASK_PP(16'h14D7D,4);
TASK_PP(16'h14D7E,4);
TASK_PP(16'h14D7F,4);
TASK_PP(16'h14D80,4);
TASK_PP(16'h14D81,4);
TASK_PP(16'h14D82,4);
TASK_PP(16'h14D83,4);
TASK_PP(16'h14D84,4);
TASK_PP(16'h14D85,4);
TASK_PP(16'h14D86,4);
TASK_PP(16'h14D87,4);
TASK_PP(16'h14D88,4);
TASK_PP(16'h14D89,4);
TASK_PP(16'h14D8A,4);
TASK_PP(16'h14D8B,4);
TASK_PP(16'h14D8C,4);
TASK_PP(16'h14D8D,4);
TASK_PP(16'h14D8E,4);
TASK_PP(16'h14D8F,4);
TASK_PP(16'h14D90,4);
TASK_PP(16'h14D91,4);
TASK_PP(16'h14D92,4);
TASK_PP(16'h14D93,4);
TASK_PP(16'h14D94,4);
TASK_PP(16'h14D95,4);
TASK_PP(16'h14D96,4);
TASK_PP(16'h14D97,4);
TASK_PP(16'h14D98,4);
TASK_PP(16'h14D99,4);
TASK_PP(16'h14D9A,4);
TASK_PP(16'h14D9B,4);
TASK_PP(16'h14D9C,4);
TASK_PP(16'h14D9D,4);
TASK_PP(16'h14D9E,4);
TASK_PP(16'h14D9F,4);
TASK_PP(16'h14DA0,4);
TASK_PP(16'h14DA1,4);
TASK_PP(16'h14DA2,4);
TASK_PP(16'h14DA3,4);
TASK_PP(16'h14DA4,4);
TASK_PP(16'h14DA5,4);
TASK_PP(16'h14DA6,4);
TASK_PP(16'h14DA7,4);
TASK_PP(16'h14DA8,4);
TASK_PP(16'h14DA9,4);
TASK_PP(16'h14DAA,4);
TASK_PP(16'h14DAB,4);
TASK_PP(16'h14DAC,4);
TASK_PP(16'h14DAD,4);
TASK_PP(16'h14DAE,4);
TASK_PP(16'h14DAF,4);
TASK_PP(16'h14DB0,4);
TASK_PP(16'h14DB1,4);
TASK_PP(16'h14DB2,4);
TASK_PP(16'h14DB3,4);
TASK_PP(16'h14DB4,4);
TASK_PP(16'h14DB5,4);
TASK_PP(16'h14DB6,4);
TASK_PP(16'h14DB7,4);
TASK_PP(16'h14DB8,4);
TASK_PP(16'h14DB9,4);
TASK_PP(16'h14DBA,4);
TASK_PP(16'h14DBB,4);
TASK_PP(16'h14DBC,4);
TASK_PP(16'h14DBD,4);
TASK_PP(16'h14DBE,4);
TASK_PP(16'h14DBF,4);
TASK_PP(16'h14DC0,4);
TASK_PP(16'h14DC1,4);
TASK_PP(16'h14DC2,4);
TASK_PP(16'h14DC3,4);
TASK_PP(16'h14DC4,4);
TASK_PP(16'h14DC5,4);
TASK_PP(16'h14DC6,4);
TASK_PP(16'h14DC7,4);
TASK_PP(16'h14DC8,4);
TASK_PP(16'h14DC9,4);
TASK_PP(16'h14DCA,4);
TASK_PP(16'h14DCB,4);
TASK_PP(16'h14DCC,4);
TASK_PP(16'h14DCD,4);
TASK_PP(16'h14DCE,4);
TASK_PP(16'h14DCF,4);
TASK_PP(16'h14DD0,4);
TASK_PP(16'h14DD1,4);
TASK_PP(16'h14DD2,4);
TASK_PP(16'h14DD3,4);
TASK_PP(16'h14DD4,4);
TASK_PP(16'h14DD5,4);
TASK_PP(16'h14DD6,4);
TASK_PP(16'h14DD7,4);
TASK_PP(16'h14DD8,4);
TASK_PP(16'h14DD9,4);
TASK_PP(16'h14DDA,4);
TASK_PP(16'h14DDB,4);
TASK_PP(16'h14DDC,4);
TASK_PP(16'h14DDD,4);
TASK_PP(16'h14DDE,4);
TASK_PP(16'h14DDF,4);
TASK_PP(16'h14DE0,4);
TASK_PP(16'h14DE1,4);
TASK_PP(16'h14DE2,4);
TASK_PP(16'h14DE3,4);
TASK_PP(16'h14DE4,4);
TASK_PP(16'h14DE5,4);
TASK_PP(16'h14DE6,4);
TASK_PP(16'h14DE7,4);
TASK_PP(16'h14DE8,4);
TASK_PP(16'h14DE9,4);
TASK_PP(16'h14DEA,4);
TASK_PP(16'h14DEB,4);
TASK_PP(16'h14DEC,4);
TASK_PP(16'h14DED,4);
TASK_PP(16'h14DEE,4);
TASK_PP(16'h14DEF,4);
TASK_PP(16'h14DF0,4);
TASK_PP(16'h14DF1,4);
TASK_PP(16'h14DF2,4);
TASK_PP(16'h14DF3,4);
TASK_PP(16'h14DF4,4);
TASK_PP(16'h14DF5,4);
TASK_PP(16'h14DF6,4);
TASK_PP(16'h14DF7,4);
TASK_PP(16'h14DF8,4);
TASK_PP(16'h14DF9,4);
TASK_PP(16'h14DFA,4);
TASK_PP(16'h14DFB,4);
TASK_PP(16'h14DFC,4);
TASK_PP(16'h14DFD,4);
TASK_PP(16'h14DFE,4);
TASK_PP(16'h14DFF,4);
TASK_PP(16'h14E00,4);
TASK_PP(16'h14E01,4);
TASK_PP(16'h14E02,4);
TASK_PP(16'h14E03,4);
TASK_PP(16'h14E04,4);
TASK_PP(16'h14E05,4);
TASK_PP(16'h14E06,4);
TASK_PP(16'h14E07,4);
TASK_PP(16'h14E08,4);
TASK_PP(16'h14E09,4);
TASK_PP(16'h14E0A,4);
TASK_PP(16'h14E0B,4);
TASK_PP(16'h14E0C,4);
TASK_PP(16'h14E0D,4);
TASK_PP(16'h14E0E,4);
TASK_PP(16'h14E0F,4);
TASK_PP(16'h14E10,4);
TASK_PP(16'h14E11,4);
TASK_PP(16'h14E12,4);
TASK_PP(16'h14E13,4);
TASK_PP(16'h14E14,4);
TASK_PP(16'h14E15,4);
TASK_PP(16'h14E16,4);
TASK_PP(16'h14E17,4);
TASK_PP(16'h14E18,4);
TASK_PP(16'h14E19,4);
TASK_PP(16'h14E1A,4);
TASK_PP(16'h14E1B,4);
TASK_PP(16'h14E1C,4);
TASK_PP(16'h14E1D,4);
TASK_PP(16'h14E1E,4);
TASK_PP(16'h14E1F,4);
TASK_PP(16'h14E20,4);
TASK_PP(16'h14E21,4);
TASK_PP(16'h14E22,4);
TASK_PP(16'h14E23,4);
TASK_PP(16'h14E24,4);
TASK_PP(16'h14E25,4);
TASK_PP(16'h14E26,4);
TASK_PP(16'h14E27,4);
TASK_PP(16'h14E28,4);
TASK_PP(16'h14E29,4);
TASK_PP(16'h14E2A,4);
TASK_PP(16'h14E2B,4);
TASK_PP(16'h14E2C,4);
TASK_PP(16'h14E2D,4);
TASK_PP(16'h14E2E,4);
TASK_PP(16'h14E2F,4);
TASK_PP(16'h14E30,4);
TASK_PP(16'h14E31,4);
TASK_PP(16'h14E32,4);
TASK_PP(16'h14E33,4);
TASK_PP(16'h14E34,4);
TASK_PP(16'h14E35,4);
TASK_PP(16'h14E36,4);
TASK_PP(16'h14E37,4);
TASK_PP(16'h14E38,4);
TASK_PP(16'h14E39,4);
TASK_PP(16'h14E3A,4);
TASK_PP(16'h14E3B,4);
TASK_PP(16'h14E3C,4);
TASK_PP(16'h14E3D,4);
TASK_PP(16'h14E3E,4);
TASK_PP(16'h14E3F,4);
TASK_PP(16'h14E40,4);
TASK_PP(16'h14E41,4);
TASK_PP(16'h14E42,4);
TASK_PP(16'h14E43,4);
TASK_PP(16'h14E44,4);
TASK_PP(16'h14E45,4);
TASK_PP(16'h14E46,4);
TASK_PP(16'h14E47,4);
TASK_PP(16'h14E48,4);
TASK_PP(16'h14E49,4);
TASK_PP(16'h14E4A,4);
TASK_PP(16'h14E4B,4);
TASK_PP(16'h14E4C,4);
TASK_PP(16'h14E4D,4);
TASK_PP(16'h14E4E,4);
TASK_PP(16'h14E4F,4);
TASK_PP(16'h14E50,4);
TASK_PP(16'h14E51,4);
TASK_PP(16'h14E52,4);
TASK_PP(16'h14E53,4);
TASK_PP(16'h14E54,4);
TASK_PP(16'h14E55,4);
TASK_PP(16'h14E56,4);
TASK_PP(16'h14E57,4);
TASK_PP(16'h14E58,4);
TASK_PP(16'h14E59,4);
TASK_PP(16'h14E5A,4);
TASK_PP(16'h14E5B,4);
TASK_PP(16'h14E5C,4);
TASK_PP(16'h14E5D,4);
TASK_PP(16'h14E5E,4);
TASK_PP(16'h14E5F,4);
TASK_PP(16'h14E60,4);
TASK_PP(16'h14E61,4);
TASK_PP(16'h14E62,4);
TASK_PP(16'h14E63,4);
TASK_PP(16'h14E64,4);
TASK_PP(16'h14E65,4);
TASK_PP(16'h14E66,4);
TASK_PP(16'h14E67,4);
TASK_PP(16'h14E68,4);
TASK_PP(16'h14E69,4);
TASK_PP(16'h14E6A,4);
TASK_PP(16'h14E6B,4);
TASK_PP(16'h14E6C,4);
TASK_PP(16'h14E6D,4);
TASK_PP(16'h14E6E,4);
TASK_PP(16'h14E6F,4);
TASK_PP(16'h14E70,4);
TASK_PP(16'h14E71,4);
TASK_PP(16'h14E72,4);
TASK_PP(16'h14E73,4);
TASK_PP(16'h14E74,4);
TASK_PP(16'h14E75,4);
TASK_PP(16'h14E76,4);
TASK_PP(16'h14E77,4);
TASK_PP(16'h14E78,4);
TASK_PP(16'h14E79,4);
TASK_PP(16'h14E7A,4);
TASK_PP(16'h14E7B,4);
TASK_PP(16'h14E7C,4);
TASK_PP(16'h14E7D,4);
TASK_PP(16'h14E7E,4);
TASK_PP(16'h14E7F,4);
TASK_PP(16'h14E80,4);
TASK_PP(16'h14E81,4);
TASK_PP(16'h14E82,4);
TASK_PP(16'h14E83,4);
TASK_PP(16'h14E84,4);
TASK_PP(16'h14E85,4);
TASK_PP(16'h14E86,4);
TASK_PP(16'h14E87,4);
TASK_PP(16'h14E88,4);
TASK_PP(16'h14E89,4);
TASK_PP(16'h14E8A,4);
TASK_PP(16'h14E8B,4);
TASK_PP(16'h14E8C,4);
TASK_PP(16'h14E8D,4);
TASK_PP(16'h14E8E,4);
TASK_PP(16'h14E8F,4);
TASK_PP(16'h14E90,4);
TASK_PP(16'h14E91,4);
TASK_PP(16'h14E92,4);
TASK_PP(16'h14E93,4);
TASK_PP(16'h14E94,4);
TASK_PP(16'h14E95,4);
TASK_PP(16'h14E96,4);
TASK_PP(16'h14E97,4);
TASK_PP(16'h14E98,4);
TASK_PP(16'h14E99,4);
TASK_PP(16'h14E9A,4);
TASK_PP(16'h14E9B,4);
TASK_PP(16'h14E9C,4);
TASK_PP(16'h14E9D,4);
TASK_PP(16'h14E9E,4);
TASK_PP(16'h14E9F,4);
TASK_PP(16'h14EA0,4);
TASK_PP(16'h14EA1,4);
TASK_PP(16'h14EA2,4);
TASK_PP(16'h14EA3,4);
TASK_PP(16'h14EA4,4);
TASK_PP(16'h14EA5,4);
TASK_PP(16'h14EA6,4);
TASK_PP(16'h14EA7,4);
TASK_PP(16'h14EA8,4);
TASK_PP(16'h14EA9,4);
TASK_PP(16'h14EAA,4);
TASK_PP(16'h14EAB,4);
TASK_PP(16'h14EAC,4);
TASK_PP(16'h14EAD,4);
TASK_PP(16'h14EAE,4);
TASK_PP(16'h14EAF,4);
TASK_PP(16'h14EB0,4);
TASK_PP(16'h14EB1,4);
TASK_PP(16'h14EB2,4);
TASK_PP(16'h14EB3,4);
TASK_PP(16'h14EB4,4);
TASK_PP(16'h14EB5,4);
TASK_PP(16'h14EB6,4);
TASK_PP(16'h14EB7,4);
TASK_PP(16'h14EB8,4);
TASK_PP(16'h14EB9,4);
TASK_PP(16'h14EBA,4);
TASK_PP(16'h14EBB,4);
TASK_PP(16'h14EBC,4);
TASK_PP(16'h14EBD,4);
TASK_PP(16'h14EBE,4);
TASK_PP(16'h14EBF,4);
TASK_PP(16'h14EC0,4);
TASK_PP(16'h14EC1,4);
TASK_PP(16'h14EC2,4);
TASK_PP(16'h14EC3,4);
TASK_PP(16'h14EC4,4);
TASK_PP(16'h14EC5,4);
TASK_PP(16'h14EC6,4);
TASK_PP(16'h14EC7,4);
TASK_PP(16'h14EC8,4);
TASK_PP(16'h14EC9,4);
TASK_PP(16'h14ECA,4);
TASK_PP(16'h14ECB,4);
TASK_PP(16'h14ECC,4);
TASK_PP(16'h14ECD,4);
TASK_PP(16'h14ECE,4);
TASK_PP(16'h14ECF,4);
TASK_PP(16'h14ED0,4);
TASK_PP(16'h14ED1,4);
TASK_PP(16'h14ED2,4);
TASK_PP(16'h14ED3,4);
TASK_PP(16'h14ED4,4);
TASK_PP(16'h14ED5,4);
TASK_PP(16'h14ED6,4);
TASK_PP(16'h14ED7,4);
TASK_PP(16'h14ED8,4);
TASK_PP(16'h14ED9,4);
TASK_PP(16'h14EDA,4);
TASK_PP(16'h14EDB,4);
TASK_PP(16'h14EDC,4);
TASK_PP(16'h14EDD,4);
TASK_PP(16'h14EDE,4);
TASK_PP(16'h14EDF,4);
TASK_PP(16'h14EE0,4);
TASK_PP(16'h14EE1,4);
TASK_PP(16'h14EE2,4);
TASK_PP(16'h14EE3,4);
TASK_PP(16'h14EE4,4);
TASK_PP(16'h14EE5,4);
TASK_PP(16'h14EE6,4);
TASK_PP(16'h14EE7,4);
TASK_PP(16'h14EE8,4);
TASK_PP(16'h14EE9,4);
TASK_PP(16'h14EEA,4);
TASK_PP(16'h14EEB,4);
TASK_PP(16'h14EEC,4);
TASK_PP(16'h14EED,4);
TASK_PP(16'h14EEE,4);
TASK_PP(16'h14EEF,4);
TASK_PP(16'h14EF0,4);
TASK_PP(16'h14EF1,4);
TASK_PP(16'h14EF2,4);
TASK_PP(16'h14EF3,4);
TASK_PP(16'h14EF4,4);
TASK_PP(16'h14EF5,4);
TASK_PP(16'h14EF6,4);
TASK_PP(16'h14EF7,4);
TASK_PP(16'h14EF8,4);
TASK_PP(16'h14EF9,4);
TASK_PP(16'h14EFA,4);
TASK_PP(16'h14EFB,4);
TASK_PP(16'h14EFC,4);
TASK_PP(16'h14EFD,4);
TASK_PP(16'h14EFE,4);
TASK_PP(16'h14EFF,4);
TASK_PP(16'h14F00,4);
TASK_PP(16'h14F01,4);
TASK_PP(16'h14F02,4);
TASK_PP(16'h14F03,4);
TASK_PP(16'h14F04,4);
TASK_PP(16'h14F05,4);
TASK_PP(16'h14F06,4);
TASK_PP(16'h14F07,4);
TASK_PP(16'h14F08,4);
TASK_PP(16'h14F09,4);
TASK_PP(16'h14F0A,4);
TASK_PP(16'h14F0B,4);
TASK_PP(16'h14F0C,4);
TASK_PP(16'h14F0D,4);
TASK_PP(16'h14F0E,4);
TASK_PP(16'h14F0F,4);
TASK_PP(16'h14F10,4);
TASK_PP(16'h14F11,4);
TASK_PP(16'h14F12,4);
TASK_PP(16'h14F13,4);
TASK_PP(16'h14F14,4);
TASK_PP(16'h14F15,4);
TASK_PP(16'h14F16,4);
TASK_PP(16'h14F17,4);
TASK_PP(16'h14F18,4);
TASK_PP(16'h14F19,4);
TASK_PP(16'h14F1A,4);
TASK_PP(16'h14F1B,4);
TASK_PP(16'h14F1C,4);
TASK_PP(16'h14F1D,4);
TASK_PP(16'h14F1E,4);
TASK_PP(16'h14F1F,4);
TASK_PP(16'h14F20,4);
TASK_PP(16'h14F21,4);
TASK_PP(16'h14F22,4);
TASK_PP(16'h14F23,4);
TASK_PP(16'h14F24,4);
TASK_PP(16'h14F25,4);
TASK_PP(16'h14F26,4);
TASK_PP(16'h14F27,4);
TASK_PP(16'h14F28,4);
TASK_PP(16'h14F29,4);
TASK_PP(16'h14F2A,4);
TASK_PP(16'h14F2B,4);
TASK_PP(16'h14F2C,4);
TASK_PP(16'h14F2D,4);
TASK_PP(16'h14F2E,4);
TASK_PP(16'h14F2F,4);
TASK_PP(16'h14F30,4);
TASK_PP(16'h14F31,4);
TASK_PP(16'h14F32,4);
TASK_PP(16'h14F33,4);
TASK_PP(16'h14F34,4);
TASK_PP(16'h14F35,4);
TASK_PP(16'h14F36,4);
TASK_PP(16'h14F37,4);
TASK_PP(16'h14F38,4);
TASK_PP(16'h14F39,4);
TASK_PP(16'h14F3A,4);
TASK_PP(16'h14F3B,4);
TASK_PP(16'h14F3C,4);
TASK_PP(16'h14F3D,4);
TASK_PP(16'h14F3E,4);
TASK_PP(16'h14F3F,4);
TASK_PP(16'h14F40,4);
TASK_PP(16'h14F41,4);
TASK_PP(16'h14F42,4);
TASK_PP(16'h14F43,4);
TASK_PP(16'h14F44,4);
TASK_PP(16'h14F45,4);
TASK_PP(16'h14F46,4);
TASK_PP(16'h14F47,4);
TASK_PP(16'h14F48,4);
TASK_PP(16'h14F49,4);
TASK_PP(16'h14F4A,4);
TASK_PP(16'h14F4B,4);
TASK_PP(16'h14F4C,4);
TASK_PP(16'h14F4D,4);
TASK_PP(16'h14F4E,4);
TASK_PP(16'h14F4F,4);
TASK_PP(16'h14F50,4);
TASK_PP(16'h14F51,4);
TASK_PP(16'h14F52,4);
TASK_PP(16'h14F53,4);
TASK_PP(16'h14F54,4);
TASK_PP(16'h14F55,4);
TASK_PP(16'h14F56,4);
TASK_PP(16'h14F57,4);
TASK_PP(16'h14F58,4);
TASK_PP(16'h14F59,4);
TASK_PP(16'h14F5A,4);
TASK_PP(16'h14F5B,4);
TASK_PP(16'h14F5C,4);
TASK_PP(16'h14F5D,4);
TASK_PP(16'h14F5E,4);
TASK_PP(16'h14F5F,4);
TASK_PP(16'h14F60,4);
TASK_PP(16'h14F61,4);
TASK_PP(16'h14F62,4);
TASK_PP(16'h14F63,4);
TASK_PP(16'h14F64,4);
TASK_PP(16'h14F65,4);
TASK_PP(16'h14F66,4);
TASK_PP(16'h14F67,4);
TASK_PP(16'h14F68,4);
TASK_PP(16'h14F69,4);
TASK_PP(16'h14F6A,4);
TASK_PP(16'h14F6B,4);
TASK_PP(16'h14F6C,4);
TASK_PP(16'h14F6D,4);
TASK_PP(16'h14F6E,4);
TASK_PP(16'h14F6F,4);
TASK_PP(16'h14F70,4);
TASK_PP(16'h14F71,4);
TASK_PP(16'h14F72,4);
TASK_PP(16'h14F73,4);
TASK_PP(16'h14F74,4);
TASK_PP(16'h14F75,4);
TASK_PP(16'h14F76,4);
TASK_PP(16'h14F77,4);
TASK_PP(16'h14F78,4);
TASK_PP(16'h14F79,4);
TASK_PP(16'h14F7A,4);
TASK_PP(16'h14F7B,4);
TASK_PP(16'h14F7C,4);
TASK_PP(16'h14F7D,4);
TASK_PP(16'h14F7E,4);
TASK_PP(16'h14F7F,4);
TASK_PP(16'h14F80,4);
TASK_PP(16'h14F81,4);
TASK_PP(16'h14F82,4);
TASK_PP(16'h14F83,4);
TASK_PP(16'h14F84,4);
TASK_PP(16'h14F85,4);
TASK_PP(16'h14F86,4);
TASK_PP(16'h14F87,4);
TASK_PP(16'h14F88,4);
TASK_PP(16'h14F89,4);
TASK_PP(16'h14F8A,4);
TASK_PP(16'h14F8B,4);
TASK_PP(16'h14F8C,4);
TASK_PP(16'h14F8D,4);
TASK_PP(16'h14F8E,4);
TASK_PP(16'h14F8F,4);
TASK_PP(16'h14F90,4);
TASK_PP(16'h14F91,4);
TASK_PP(16'h14F92,4);
TASK_PP(16'h14F93,4);
TASK_PP(16'h14F94,4);
TASK_PP(16'h14F95,4);
TASK_PP(16'h14F96,4);
TASK_PP(16'h14F97,4);
TASK_PP(16'h14F98,4);
TASK_PP(16'h14F99,4);
TASK_PP(16'h14F9A,4);
TASK_PP(16'h14F9B,4);
TASK_PP(16'h14F9C,4);
TASK_PP(16'h14F9D,4);
TASK_PP(16'h14F9E,4);
TASK_PP(16'h14F9F,4);
TASK_PP(16'h14FA0,4);
TASK_PP(16'h14FA1,4);
TASK_PP(16'h14FA2,4);
TASK_PP(16'h14FA3,4);
TASK_PP(16'h14FA4,4);
TASK_PP(16'h14FA5,4);
TASK_PP(16'h14FA6,4);
TASK_PP(16'h14FA7,4);
TASK_PP(16'h14FA8,4);
TASK_PP(16'h14FA9,4);
TASK_PP(16'h14FAA,4);
TASK_PP(16'h14FAB,4);
TASK_PP(16'h14FAC,4);
TASK_PP(16'h14FAD,4);
TASK_PP(16'h14FAE,4);
TASK_PP(16'h14FAF,4);
TASK_PP(16'h14FB0,4);
TASK_PP(16'h14FB1,4);
TASK_PP(16'h14FB2,4);
TASK_PP(16'h14FB3,4);
TASK_PP(16'h14FB4,4);
TASK_PP(16'h14FB5,4);
TASK_PP(16'h14FB6,4);
TASK_PP(16'h14FB7,4);
TASK_PP(16'h14FB8,4);
TASK_PP(16'h14FB9,4);
TASK_PP(16'h14FBA,4);
TASK_PP(16'h14FBB,4);
TASK_PP(16'h14FBC,4);
TASK_PP(16'h14FBD,4);
TASK_PP(16'h14FBE,4);
TASK_PP(16'h14FBF,4);
TASK_PP(16'h14FC0,4);
TASK_PP(16'h14FC1,4);
TASK_PP(16'h14FC2,4);
TASK_PP(16'h14FC3,4);
TASK_PP(16'h14FC4,4);
TASK_PP(16'h14FC5,4);
TASK_PP(16'h14FC6,4);
TASK_PP(16'h14FC7,4);
TASK_PP(16'h14FC8,4);
TASK_PP(16'h14FC9,4);
TASK_PP(16'h14FCA,4);
TASK_PP(16'h14FCB,4);
TASK_PP(16'h14FCC,4);
TASK_PP(16'h14FCD,4);
TASK_PP(16'h14FCE,4);
TASK_PP(16'h14FCF,4);
TASK_PP(16'h14FD0,4);
TASK_PP(16'h14FD1,4);
TASK_PP(16'h14FD2,4);
TASK_PP(16'h14FD3,4);
TASK_PP(16'h14FD4,4);
TASK_PP(16'h14FD5,4);
TASK_PP(16'h14FD6,4);
TASK_PP(16'h14FD7,4);
TASK_PP(16'h14FD8,4);
TASK_PP(16'h14FD9,4);
TASK_PP(16'h14FDA,4);
TASK_PP(16'h14FDB,4);
TASK_PP(16'h14FDC,4);
TASK_PP(16'h14FDD,4);
TASK_PP(16'h14FDE,4);
TASK_PP(16'h14FDF,4);
TASK_PP(16'h14FE0,4);
TASK_PP(16'h14FE1,4);
TASK_PP(16'h14FE2,4);
TASK_PP(16'h14FE3,4);
TASK_PP(16'h14FE4,4);
TASK_PP(16'h14FE5,4);
TASK_PP(16'h14FE6,4);
TASK_PP(16'h14FE7,4);
TASK_PP(16'h14FE8,4);
TASK_PP(16'h14FE9,4);
TASK_PP(16'h14FEA,4);
TASK_PP(16'h14FEB,4);
TASK_PP(16'h14FEC,4);
TASK_PP(16'h14FED,4);
TASK_PP(16'h14FEE,4);
TASK_PP(16'h14FEF,4);
TASK_PP(16'h14FF0,4);
TASK_PP(16'h14FF1,4);
TASK_PP(16'h14FF2,4);
TASK_PP(16'h14FF3,4);
TASK_PP(16'h14FF4,4);
TASK_PP(16'h14FF5,4);
TASK_PP(16'h14FF6,4);
TASK_PP(16'h14FF7,4);
TASK_PP(16'h14FF8,4);
TASK_PP(16'h14FF9,4);
TASK_PP(16'h14FFA,4);
TASK_PP(16'h14FFB,4);
TASK_PP(16'h14FFC,4);
TASK_PP(16'h14FFD,4);
TASK_PP(16'h14FFE,4);
TASK_PP(16'h14FFF,4);
TASK_PP(16'h15000,4);
TASK_PP(16'h15001,4);
TASK_PP(16'h15002,4);
TASK_PP(16'h15003,4);
TASK_PP(16'h15004,4);
TASK_PP(16'h15005,4);
TASK_PP(16'h15006,4);
TASK_PP(16'h15007,4);
TASK_PP(16'h15008,4);
TASK_PP(16'h15009,4);
TASK_PP(16'h1500A,4);
TASK_PP(16'h1500B,4);
TASK_PP(16'h1500C,4);
TASK_PP(16'h1500D,4);
TASK_PP(16'h1500E,4);
TASK_PP(16'h1500F,4);
TASK_PP(16'h15010,4);
TASK_PP(16'h15011,4);
TASK_PP(16'h15012,4);
TASK_PP(16'h15013,4);
TASK_PP(16'h15014,4);
TASK_PP(16'h15015,4);
TASK_PP(16'h15016,4);
TASK_PP(16'h15017,4);
TASK_PP(16'h15018,4);
TASK_PP(16'h15019,4);
TASK_PP(16'h1501A,4);
TASK_PP(16'h1501B,4);
TASK_PP(16'h1501C,4);
TASK_PP(16'h1501D,4);
TASK_PP(16'h1501E,4);
TASK_PP(16'h1501F,4);
TASK_PP(16'h15020,4);
TASK_PP(16'h15021,4);
TASK_PP(16'h15022,4);
TASK_PP(16'h15023,4);
TASK_PP(16'h15024,4);
TASK_PP(16'h15025,4);
TASK_PP(16'h15026,4);
TASK_PP(16'h15027,4);
TASK_PP(16'h15028,4);
TASK_PP(16'h15029,4);
TASK_PP(16'h1502A,4);
TASK_PP(16'h1502B,4);
TASK_PP(16'h1502C,4);
TASK_PP(16'h1502D,4);
TASK_PP(16'h1502E,4);
TASK_PP(16'h1502F,4);
TASK_PP(16'h15030,4);
TASK_PP(16'h15031,4);
TASK_PP(16'h15032,4);
TASK_PP(16'h15033,4);
TASK_PP(16'h15034,4);
TASK_PP(16'h15035,4);
TASK_PP(16'h15036,4);
TASK_PP(16'h15037,4);
TASK_PP(16'h15038,4);
TASK_PP(16'h15039,4);
TASK_PP(16'h1503A,4);
TASK_PP(16'h1503B,4);
TASK_PP(16'h1503C,4);
TASK_PP(16'h1503D,4);
TASK_PP(16'h1503E,4);
TASK_PP(16'h1503F,4);
TASK_PP(16'h15040,4);
TASK_PP(16'h15041,4);
TASK_PP(16'h15042,4);
TASK_PP(16'h15043,4);
TASK_PP(16'h15044,4);
TASK_PP(16'h15045,4);
TASK_PP(16'h15046,4);
TASK_PP(16'h15047,4);
TASK_PP(16'h15048,4);
TASK_PP(16'h15049,4);
TASK_PP(16'h1504A,4);
TASK_PP(16'h1504B,4);
TASK_PP(16'h1504C,4);
TASK_PP(16'h1504D,4);
TASK_PP(16'h1504E,4);
TASK_PP(16'h1504F,4);
TASK_PP(16'h15050,4);
TASK_PP(16'h15051,4);
TASK_PP(16'h15052,4);
TASK_PP(16'h15053,4);
TASK_PP(16'h15054,4);
TASK_PP(16'h15055,4);
TASK_PP(16'h15056,4);
TASK_PP(16'h15057,4);
TASK_PP(16'h15058,4);
TASK_PP(16'h15059,4);
TASK_PP(16'h1505A,4);
TASK_PP(16'h1505B,4);
TASK_PP(16'h1505C,4);
TASK_PP(16'h1505D,4);
TASK_PP(16'h1505E,4);
TASK_PP(16'h1505F,4);
TASK_PP(16'h15060,4);
TASK_PP(16'h15061,4);
TASK_PP(16'h15062,4);
TASK_PP(16'h15063,4);
TASK_PP(16'h15064,4);
TASK_PP(16'h15065,4);
TASK_PP(16'h15066,4);
TASK_PP(16'h15067,4);
TASK_PP(16'h15068,4);
TASK_PP(16'h15069,4);
TASK_PP(16'h1506A,4);
TASK_PP(16'h1506B,4);
TASK_PP(16'h1506C,4);
TASK_PP(16'h1506D,4);
TASK_PP(16'h1506E,4);
TASK_PP(16'h1506F,4);
TASK_PP(16'h15070,4);
TASK_PP(16'h15071,4);
TASK_PP(16'h15072,4);
TASK_PP(16'h15073,4);
TASK_PP(16'h15074,4);
TASK_PP(16'h15075,4);
TASK_PP(16'h15076,4);
TASK_PP(16'h15077,4);
TASK_PP(16'h15078,4);
TASK_PP(16'h15079,4);
TASK_PP(16'h1507A,4);
TASK_PP(16'h1507B,4);
TASK_PP(16'h1507C,4);
TASK_PP(16'h1507D,4);
TASK_PP(16'h1507E,4);
TASK_PP(16'h1507F,4);
TASK_PP(16'h15080,4);
TASK_PP(16'h15081,4);
TASK_PP(16'h15082,4);
TASK_PP(16'h15083,4);
TASK_PP(16'h15084,4);
TASK_PP(16'h15085,4);
TASK_PP(16'h15086,4);
TASK_PP(16'h15087,4);
TASK_PP(16'h15088,4);
TASK_PP(16'h15089,4);
TASK_PP(16'h1508A,4);
TASK_PP(16'h1508B,4);
TASK_PP(16'h1508C,4);
TASK_PP(16'h1508D,4);
TASK_PP(16'h1508E,4);
TASK_PP(16'h1508F,4);
TASK_PP(16'h15090,4);
TASK_PP(16'h15091,4);
TASK_PP(16'h15092,4);
TASK_PP(16'h15093,4);
TASK_PP(16'h15094,4);
TASK_PP(16'h15095,4);
TASK_PP(16'h15096,4);
TASK_PP(16'h15097,4);
TASK_PP(16'h15098,4);
TASK_PP(16'h15099,4);
TASK_PP(16'h1509A,4);
TASK_PP(16'h1509B,4);
TASK_PP(16'h1509C,4);
TASK_PP(16'h1509D,4);
TASK_PP(16'h1509E,4);
TASK_PP(16'h1509F,4);
TASK_PP(16'h150A0,4);
TASK_PP(16'h150A1,4);
TASK_PP(16'h150A2,4);
TASK_PP(16'h150A3,4);
TASK_PP(16'h150A4,4);
TASK_PP(16'h150A5,4);
TASK_PP(16'h150A6,4);
TASK_PP(16'h150A7,4);
TASK_PP(16'h150A8,4);
TASK_PP(16'h150A9,4);
TASK_PP(16'h150AA,4);
TASK_PP(16'h150AB,4);
TASK_PP(16'h150AC,4);
TASK_PP(16'h150AD,4);
TASK_PP(16'h150AE,4);
TASK_PP(16'h150AF,4);
TASK_PP(16'h150B0,4);
TASK_PP(16'h150B1,4);
TASK_PP(16'h150B2,4);
TASK_PP(16'h150B3,4);
TASK_PP(16'h150B4,4);
TASK_PP(16'h150B5,4);
TASK_PP(16'h150B6,4);
TASK_PP(16'h150B7,4);
TASK_PP(16'h150B8,4);
TASK_PP(16'h150B9,4);
TASK_PP(16'h150BA,4);
TASK_PP(16'h150BB,4);
TASK_PP(16'h150BC,4);
TASK_PP(16'h150BD,4);
TASK_PP(16'h150BE,4);
TASK_PP(16'h150BF,4);
TASK_PP(16'h150C0,4);
TASK_PP(16'h150C1,4);
TASK_PP(16'h150C2,4);
TASK_PP(16'h150C3,4);
TASK_PP(16'h150C4,4);
TASK_PP(16'h150C5,4);
TASK_PP(16'h150C6,4);
TASK_PP(16'h150C7,4);
TASK_PP(16'h150C8,4);
TASK_PP(16'h150C9,4);
TASK_PP(16'h150CA,4);
TASK_PP(16'h150CB,4);
TASK_PP(16'h150CC,4);
TASK_PP(16'h150CD,4);
TASK_PP(16'h150CE,4);
TASK_PP(16'h150CF,4);
TASK_PP(16'h150D0,4);
TASK_PP(16'h150D1,4);
TASK_PP(16'h150D2,4);
TASK_PP(16'h150D3,4);
TASK_PP(16'h150D4,4);
TASK_PP(16'h150D5,4);
TASK_PP(16'h150D6,4);
TASK_PP(16'h150D7,4);
TASK_PP(16'h150D8,4);
TASK_PP(16'h150D9,4);
TASK_PP(16'h150DA,4);
TASK_PP(16'h150DB,4);
TASK_PP(16'h150DC,4);
TASK_PP(16'h150DD,4);
TASK_PP(16'h150DE,4);
TASK_PP(16'h150DF,4);
TASK_PP(16'h150E0,4);
TASK_PP(16'h150E1,4);
TASK_PP(16'h150E2,4);
TASK_PP(16'h150E3,4);
TASK_PP(16'h150E4,4);
TASK_PP(16'h150E5,4);
TASK_PP(16'h150E6,4);
TASK_PP(16'h150E7,4);
TASK_PP(16'h150E8,4);
TASK_PP(16'h150E9,4);
TASK_PP(16'h150EA,4);
TASK_PP(16'h150EB,4);
TASK_PP(16'h150EC,4);
TASK_PP(16'h150ED,4);
TASK_PP(16'h150EE,4);
TASK_PP(16'h150EF,4);
TASK_PP(16'h150F0,4);
TASK_PP(16'h150F1,4);
TASK_PP(16'h150F2,4);
TASK_PP(16'h150F3,4);
TASK_PP(16'h150F4,4);
TASK_PP(16'h150F5,4);
TASK_PP(16'h150F6,4);
TASK_PP(16'h150F7,4);
TASK_PP(16'h150F8,4);
TASK_PP(16'h150F9,4);
TASK_PP(16'h150FA,4);
TASK_PP(16'h150FB,4);
TASK_PP(16'h150FC,4);
TASK_PP(16'h150FD,4);
TASK_PP(16'h150FE,4);
TASK_PP(16'h150FF,4);
TASK_PP(16'h15100,4);
TASK_PP(16'h15101,4);
TASK_PP(16'h15102,4);
TASK_PP(16'h15103,4);
TASK_PP(16'h15104,4);
TASK_PP(16'h15105,4);
TASK_PP(16'h15106,4);
TASK_PP(16'h15107,4);
TASK_PP(16'h15108,4);
TASK_PP(16'h15109,4);
TASK_PP(16'h1510A,4);
TASK_PP(16'h1510B,4);
TASK_PP(16'h1510C,4);
TASK_PP(16'h1510D,4);
TASK_PP(16'h1510E,4);
TASK_PP(16'h1510F,4);
TASK_PP(16'h15110,4);
TASK_PP(16'h15111,4);
TASK_PP(16'h15112,4);
TASK_PP(16'h15113,4);
TASK_PP(16'h15114,4);
TASK_PP(16'h15115,4);
TASK_PP(16'h15116,4);
TASK_PP(16'h15117,4);
TASK_PP(16'h15118,4);
TASK_PP(16'h15119,4);
TASK_PP(16'h1511A,4);
TASK_PP(16'h1511B,4);
TASK_PP(16'h1511C,4);
TASK_PP(16'h1511D,4);
TASK_PP(16'h1511E,4);
TASK_PP(16'h1511F,4);
TASK_PP(16'h15120,4);
TASK_PP(16'h15121,4);
TASK_PP(16'h15122,4);
TASK_PP(16'h15123,4);
TASK_PP(16'h15124,4);
TASK_PP(16'h15125,4);
TASK_PP(16'h15126,4);
TASK_PP(16'h15127,4);
TASK_PP(16'h15128,4);
TASK_PP(16'h15129,4);
TASK_PP(16'h1512A,4);
TASK_PP(16'h1512B,4);
TASK_PP(16'h1512C,4);
TASK_PP(16'h1512D,4);
TASK_PP(16'h1512E,4);
TASK_PP(16'h1512F,4);
TASK_PP(16'h15130,4);
TASK_PP(16'h15131,4);
TASK_PP(16'h15132,4);
TASK_PP(16'h15133,4);
TASK_PP(16'h15134,4);
TASK_PP(16'h15135,4);
TASK_PP(16'h15136,4);
TASK_PP(16'h15137,4);
TASK_PP(16'h15138,4);
TASK_PP(16'h15139,4);
TASK_PP(16'h1513A,4);
TASK_PP(16'h1513B,4);
TASK_PP(16'h1513C,4);
TASK_PP(16'h1513D,4);
TASK_PP(16'h1513E,4);
TASK_PP(16'h1513F,4);
TASK_PP(16'h15140,4);
TASK_PP(16'h15141,4);
TASK_PP(16'h15142,4);
TASK_PP(16'h15143,4);
TASK_PP(16'h15144,4);
TASK_PP(16'h15145,4);
TASK_PP(16'h15146,4);
TASK_PP(16'h15147,4);
TASK_PP(16'h15148,4);
TASK_PP(16'h15149,4);
TASK_PP(16'h1514A,4);
TASK_PP(16'h1514B,4);
TASK_PP(16'h1514C,4);
TASK_PP(16'h1514D,4);
TASK_PP(16'h1514E,4);
TASK_PP(16'h1514F,4);
TASK_PP(16'h15150,4);
TASK_PP(16'h15151,4);
TASK_PP(16'h15152,4);
TASK_PP(16'h15153,4);
TASK_PP(16'h15154,4);
TASK_PP(16'h15155,4);
TASK_PP(16'h15156,4);
TASK_PP(16'h15157,4);
TASK_PP(16'h15158,4);
TASK_PP(16'h15159,4);
TASK_PP(16'h1515A,4);
TASK_PP(16'h1515B,4);
TASK_PP(16'h1515C,4);
TASK_PP(16'h1515D,4);
TASK_PP(16'h1515E,4);
TASK_PP(16'h1515F,4);
TASK_PP(16'h15160,4);
TASK_PP(16'h15161,4);
TASK_PP(16'h15162,4);
TASK_PP(16'h15163,4);
TASK_PP(16'h15164,4);
TASK_PP(16'h15165,4);
TASK_PP(16'h15166,4);
TASK_PP(16'h15167,4);
TASK_PP(16'h15168,4);
TASK_PP(16'h15169,4);
TASK_PP(16'h1516A,4);
TASK_PP(16'h1516B,4);
TASK_PP(16'h1516C,4);
TASK_PP(16'h1516D,4);
TASK_PP(16'h1516E,4);
TASK_PP(16'h1516F,4);
TASK_PP(16'h15170,4);
TASK_PP(16'h15171,4);
TASK_PP(16'h15172,4);
TASK_PP(16'h15173,4);
TASK_PP(16'h15174,4);
TASK_PP(16'h15175,4);
TASK_PP(16'h15176,4);
TASK_PP(16'h15177,4);
TASK_PP(16'h15178,4);
TASK_PP(16'h15179,4);
TASK_PP(16'h1517A,4);
TASK_PP(16'h1517B,4);
TASK_PP(16'h1517C,4);
TASK_PP(16'h1517D,4);
TASK_PP(16'h1517E,4);
TASK_PP(16'h1517F,4);
TASK_PP(16'h15180,4);
TASK_PP(16'h15181,4);
TASK_PP(16'h15182,4);
TASK_PP(16'h15183,4);
TASK_PP(16'h15184,4);
TASK_PP(16'h15185,4);
TASK_PP(16'h15186,4);
TASK_PP(16'h15187,4);
TASK_PP(16'h15188,4);
TASK_PP(16'h15189,4);
TASK_PP(16'h1518A,4);
TASK_PP(16'h1518B,4);
TASK_PP(16'h1518C,4);
TASK_PP(16'h1518D,4);
TASK_PP(16'h1518E,4);
TASK_PP(16'h1518F,4);
TASK_PP(16'h15190,4);
TASK_PP(16'h15191,4);
TASK_PP(16'h15192,4);
TASK_PP(16'h15193,4);
TASK_PP(16'h15194,4);
TASK_PP(16'h15195,4);
TASK_PP(16'h15196,4);
TASK_PP(16'h15197,4);
TASK_PP(16'h15198,4);
TASK_PP(16'h15199,4);
TASK_PP(16'h1519A,4);
TASK_PP(16'h1519B,4);
TASK_PP(16'h1519C,4);
TASK_PP(16'h1519D,4);
TASK_PP(16'h1519E,4);
TASK_PP(16'h1519F,4);
TASK_PP(16'h151A0,4);
TASK_PP(16'h151A1,4);
TASK_PP(16'h151A2,4);
TASK_PP(16'h151A3,4);
TASK_PP(16'h151A4,4);
TASK_PP(16'h151A5,4);
TASK_PP(16'h151A6,4);
TASK_PP(16'h151A7,4);
TASK_PP(16'h151A8,4);
TASK_PP(16'h151A9,4);
TASK_PP(16'h151AA,4);
TASK_PP(16'h151AB,4);
TASK_PP(16'h151AC,4);
TASK_PP(16'h151AD,4);
TASK_PP(16'h151AE,4);
TASK_PP(16'h151AF,4);
TASK_PP(16'h151B0,4);
TASK_PP(16'h151B1,4);
TASK_PP(16'h151B2,4);
TASK_PP(16'h151B3,4);
TASK_PP(16'h151B4,4);
TASK_PP(16'h151B5,4);
TASK_PP(16'h151B6,4);
TASK_PP(16'h151B7,4);
TASK_PP(16'h151B8,4);
TASK_PP(16'h151B9,4);
TASK_PP(16'h151BA,4);
TASK_PP(16'h151BB,4);
TASK_PP(16'h151BC,4);
TASK_PP(16'h151BD,4);
TASK_PP(16'h151BE,4);
TASK_PP(16'h151BF,4);
TASK_PP(16'h151C0,4);
TASK_PP(16'h151C1,4);
TASK_PP(16'h151C2,4);
TASK_PP(16'h151C3,4);
TASK_PP(16'h151C4,4);
TASK_PP(16'h151C5,4);
TASK_PP(16'h151C6,4);
TASK_PP(16'h151C7,4);
TASK_PP(16'h151C8,4);
TASK_PP(16'h151C9,4);
TASK_PP(16'h151CA,4);
TASK_PP(16'h151CB,4);
TASK_PP(16'h151CC,4);
TASK_PP(16'h151CD,4);
TASK_PP(16'h151CE,4);
TASK_PP(16'h151CF,4);
TASK_PP(16'h151D0,4);
TASK_PP(16'h151D1,4);
TASK_PP(16'h151D2,4);
TASK_PP(16'h151D3,4);
TASK_PP(16'h151D4,4);
TASK_PP(16'h151D5,4);
TASK_PP(16'h151D6,4);
TASK_PP(16'h151D7,4);
TASK_PP(16'h151D8,4);
TASK_PP(16'h151D9,4);
TASK_PP(16'h151DA,4);
TASK_PP(16'h151DB,4);
TASK_PP(16'h151DC,4);
TASK_PP(16'h151DD,4);
TASK_PP(16'h151DE,4);
TASK_PP(16'h151DF,4);
TASK_PP(16'h151E0,4);
TASK_PP(16'h151E1,4);
TASK_PP(16'h151E2,4);
TASK_PP(16'h151E3,4);
TASK_PP(16'h151E4,4);
TASK_PP(16'h151E5,4);
TASK_PP(16'h151E6,4);
TASK_PP(16'h151E7,4);
TASK_PP(16'h151E8,4);
TASK_PP(16'h151E9,4);
TASK_PP(16'h151EA,4);
TASK_PP(16'h151EB,4);
TASK_PP(16'h151EC,4);
TASK_PP(16'h151ED,4);
TASK_PP(16'h151EE,4);
TASK_PP(16'h151EF,4);
TASK_PP(16'h151F0,4);
TASK_PP(16'h151F1,4);
TASK_PP(16'h151F2,4);
TASK_PP(16'h151F3,4);
TASK_PP(16'h151F4,4);
TASK_PP(16'h151F5,4);
TASK_PP(16'h151F6,4);
TASK_PP(16'h151F7,4);
TASK_PP(16'h151F8,4);
TASK_PP(16'h151F9,4);
TASK_PP(16'h151FA,4);
TASK_PP(16'h151FB,4);
TASK_PP(16'h151FC,4);
TASK_PP(16'h151FD,4);
TASK_PP(16'h151FE,4);
TASK_PP(16'h151FF,4);
TASK_PP(16'h15200,4);
TASK_PP(16'h15201,4);
TASK_PP(16'h15202,4);
TASK_PP(16'h15203,4);
TASK_PP(16'h15204,4);
TASK_PP(16'h15205,4);
TASK_PP(16'h15206,4);
TASK_PP(16'h15207,4);
TASK_PP(16'h15208,4);
TASK_PP(16'h15209,4);
TASK_PP(16'h1520A,4);
TASK_PP(16'h1520B,4);
TASK_PP(16'h1520C,4);
TASK_PP(16'h1520D,4);
TASK_PP(16'h1520E,4);
TASK_PP(16'h1520F,4);
TASK_PP(16'h15210,4);
TASK_PP(16'h15211,4);
TASK_PP(16'h15212,4);
TASK_PP(16'h15213,4);
TASK_PP(16'h15214,4);
TASK_PP(16'h15215,4);
TASK_PP(16'h15216,4);
TASK_PP(16'h15217,4);
TASK_PP(16'h15218,4);
TASK_PP(16'h15219,4);
TASK_PP(16'h1521A,4);
TASK_PP(16'h1521B,4);
TASK_PP(16'h1521C,4);
TASK_PP(16'h1521D,4);
TASK_PP(16'h1521E,4);
TASK_PP(16'h1521F,4);
TASK_PP(16'h15220,4);
TASK_PP(16'h15221,4);
TASK_PP(16'h15222,4);
TASK_PP(16'h15223,4);
TASK_PP(16'h15224,4);
TASK_PP(16'h15225,4);
TASK_PP(16'h15226,4);
TASK_PP(16'h15227,4);
TASK_PP(16'h15228,4);
TASK_PP(16'h15229,4);
TASK_PP(16'h1522A,4);
TASK_PP(16'h1522B,4);
TASK_PP(16'h1522C,4);
TASK_PP(16'h1522D,4);
TASK_PP(16'h1522E,4);
TASK_PP(16'h1522F,4);
TASK_PP(16'h15230,4);
TASK_PP(16'h15231,4);
TASK_PP(16'h15232,4);
TASK_PP(16'h15233,4);
TASK_PP(16'h15234,4);
TASK_PP(16'h15235,4);
TASK_PP(16'h15236,4);
TASK_PP(16'h15237,4);
TASK_PP(16'h15238,4);
TASK_PP(16'h15239,4);
TASK_PP(16'h1523A,4);
TASK_PP(16'h1523B,4);
TASK_PP(16'h1523C,4);
TASK_PP(16'h1523D,4);
TASK_PP(16'h1523E,4);
TASK_PP(16'h1523F,4);
TASK_PP(16'h15240,4);
TASK_PP(16'h15241,4);
TASK_PP(16'h15242,4);
TASK_PP(16'h15243,4);
TASK_PP(16'h15244,4);
TASK_PP(16'h15245,4);
TASK_PP(16'h15246,4);
TASK_PP(16'h15247,4);
TASK_PP(16'h15248,4);
TASK_PP(16'h15249,4);
TASK_PP(16'h1524A,4);
TASK_PP(16'h1524B,4);
TASK_PP(16'h1524C,4);
TASK_PP(16'h1524D,4);
TASK_PP(16'h1524E,4);
TASK_PP(16'h1524F,4);
TASK_PP(16'h15250,4);
TASK_PP(16'h15251,4);
TASK_PP(16'h15252,4);
TASK_PP(16'h15253,4);
TASK_PP(16'h15254,4);
TASK_PP(16'h15255,4);
TASK_PP(16'h15256,4);
TASK_PP(16'h15257,4);
TASK_PP(16'h15258,4);
TASK_PP(16'h15259,4);
TASK_PP(16'h1525A,4);
TASK_PP(16'h1525B,4);
TASK_PP(16'h1525C,4);
TASK_PP(16'h1525D,4);
TASK_PP(16'h1525E,4);
TASK_PP(16'h1525F,4);
TASK_PP(16'h15260,4);
TASK_PP(16'h15261,4);
TASK_PP(16'h15262,4);
TASK_PP(16'h15263,4);
TASK_PP(16'h15264,4);
TASK_PP(16'h15265,4);
TASK_PP(16'h15266,4);
TASK_PP(16'h15267,4);
TASK_PP(16'h15268,4);
TASK_PP(16'h15269,4);
TASK_PP(16'h1526A,4);
TASK_PP(16'h1526B,4);
TASK_PP(16'h1526C,4);
TASK_PP(16'h1526D,4);
TASK_PP(16'h1526E,4);
TASK_PP(16'h1526F,4);
TASK_PP(16'h15270,4);
TASK_PP(16'h15271,4);
TASK_PP(16'h15272,4);
TASK_PP(16'h15273,4);
TASK_PP(16'h15274,4);
TASK_PP(16'h15275,4);
TASK_PP(16'h15276,4);
TASK_PP(16'h15277,4);
TASK_PP(16'h15278,4);
TASK_PP(16'h15279,4);
TASK_PP(16'h1527A,4);
TASK_PP(16'h1527B,4);
TASK_PP(16'h1527C,4);
TASK_PP(16'h1527D,4);
TASK_PP(16'h1527E,4);
TASK_PP(16'h1527F,4);
TASK_PP(16'h15280,4);
TASK_PP(16'h15281,4);
TASK_PP(16'h15282,4);
TASK_PP(16'h15283,4);
TASK_PP(16'h15284,4);
TASK_PP(16'h15285,4);
TASK_PP(16'h15286,4);
TASK_PP(16'h15287,4);
TASK_PP(16'h15288,4);
TASK_PP(16'h15289,4);
TASK_PP(16'h1528A,4);
TASK_PP(16'h1528B,4);
TASK_PP(16'h1528C,4);
TASK_PP(16'h1528D,4);
TASK_PP(16'h1528E,4);
TASK_PP(16'h1528F,4);
TASK_PP(16'h15290,4);
TASK_PP(16'h15291,4);
TASK_PP(16'h15292,4);
TASK_PP(16'h15293,4);
TASK_PP(16'h15294,4);
TASK_PP(16'h15295,4);
TASK_PP(16'h15296,4);
TASK_PP(16'h15297,4);
TASK_PP(16'h15298,4);
TASK_PP(16'h15299,4);
TASK_PP(16'h1529A,4);
TASK_PP(16'h1529B,4);
TASK_PP(16'h1529C,4);
TASK_PP(16'h1529D,4);
TASK_PP(16'h1529E,4);
TASK_PP(16'h1529F,4);
TASK_PP(16'h152A0,4);
TASK_PP(16'h152A1,4);
TASK_PP(16'h152A2,4);
TASK_PP(16'h152A3,4);
TASK_PP(16'h152A4,4);
TASK_PP(16'h152A5,4);
TASK_PP(16'h152A6,4);
TASK_PP(16'h152A7,4);
TASK_PP(16'h152A8,4);
TASK_PP(16'h152A9,4);
TASK_PP(16'h152AA,4);
TASK_PP(16'h152AB,4);
TASK_PP(16'h152AC,4);
TASK_PP(16'h152AD,4);
TASK_PP(16'h152AE,4);
TASK_PP(16'h152AF,4);
TASK_PP(16'h152B0,4);
TASK_PP(16'h152B1,4);
TASK_PP(16'h152B2,4);
TASK_PP(16'h152B3,4);
TASK_PP(16'h152B4,4);
TASK_PP(16'h152B5,4);
TASK_PP(16'h152B6,4);
TASK_PP(16'h152B7,4);
TASK_PP(16'h152B8,4);
TASK_PP(16'h152B9,4);
TASK_PP(16'h152BA,4);
TASK_PP(16'h152BB,4);
TASK_PP(16'h152BC,4);
TASK_PP(16'h152BD,4);
TASK_PP(16'h152BE,4);
TASK_PP(16'h152BF,4);
TASK_PP(16'h152C0,4);
TASK_PP(16'h152C1,4);
TASK_PP(16'h152C2,4);
TASK_PP(16'h152C3,4);
TASK_PP(16'h152C4,4);
TASK_PP(16'h152C5,4);
TASK_PP(16'h152C6,4);
TASK_PP(16'h152C7,4);
TASK_PP(16'h152C8,4);
TASK_PP(16'h152C9,4);
TASK_PP(16'h152CA,4);
TASK_PP(16'h152CB,4);
TASK_PP(16'h152CC,4);
TASK_PP(16'h152CD,4);
TASK_PP(16'h152CE,4);
TASK_PP(16'h152CF,4);
TASK_PP(16'h152D0,4);
TASK_PP(16'h152D1,4);
TASK_PP(16'h152D2,4);
TASK_PP(16'h152D3,4);
TASK_PP(16'h152D4,4);
TASK_PP(16'h152D5,4);
TASK_PP(16'h152D6,4);
TASK_PP(16'h152D7,4);
TASK_PP(16'h152D8,4);
TASK_PP(16'h152D9,4);
TASK_PP(16'h152DA,4);
TASK_PP(16'h152DB,4);
TASK_PP(16'h152DC,4);
TASK_PP(16'h152DD,4);
TASK_PP(16'h152DE,4);
TASK_PP(16'h152DF,4);
TASK_PP(16'h152E0,4);
TASK_PP(16'h152E1,4);
TASK_PP(16'h152E2,4);
TASK_PP(16'h152E3,4);
TASK_PP(16'h152E4,4);
TASK_PP(16'h152E5,4);
TASK_PP(16'h152E6,4);
TASK_PP(16'h152E7,4);
TASK_PP(16'h152E8,4);
TASK_PP(16'h152E9,4);
TASK_PP(16'h152EA,4);
TASK_PP(16'h152EB,4);
TASK_PP(16'h152EC,4);
TASK_PP(16'h152ED,4);
TASK_PP(16'h152EE,4);
TASK_PP(16'h152EF,4);
TASK_PP(16'h152F0,4);
TASK_PP(16'h152F1,4);
TASK_PP(16'h152F2,4);
TASK_PP(16'h152F3,4);
TASK_PP(16'h152F4,4);
TASK_PP(16'h152F5,4);
TASK_PP(16'h152F6,4);
TASK_PP(16'h152F7,4);
TASK_PP(16'h152F8,4);
TASK_PP(16'h152F9,4);
TASK_PP(16'h152FA,4);
TASK_PP(16'h152FB,4);
TASK_PP(16'h152FC,4);
TASK_PP(16'h152FD,4);
TASK_PP(16'h152FE,4);
TASK_PP(16'h152FF,4);
TASK_PP(16'h15300,4);
TASK_PP(16'h15301,4);
TASK_PP(16'h15302,4);
TASK_PP(16'h15303,4);
TASK_PP(16'h15304,4);
TASK_PP(16'h15305,4);
TASK_PP(16'h15306,4);
TASK_PP(16'h15307,4);
TASK_PP(16'h15308,4);
TASK_PP(16'h15309,4);
TASK_PP(16'h1530A,4);
TASK_PP(16'h1530B,4);
TASK_PP(16'h1530C,4);
TASK_PP(16'h1530D,4);
TASK_PP(16'h1530E,4);
TASK_PP(16'h1530F,4);
TASK_PP(16'h15310,4);
TASK_PP(16'h15311,4);
TASK_PP(16'h15312,4);
TASK_PP(16'h15313,4);
TASK_PP(16'h15314,4);
TASK_PP(16'h15315,4);
TASK_PP(16'h15316,4);
TASK_PP(16'h15317,4);
TASK_PP(16'h15318,4);
TASK_PP(16'h15319,4);
TASK_PP(16'h1531A,4);
TASK_PP(16'h1531B,4);
TASK_PP(16'h1531C,4);
TASK_PP(16'h1531D,4);
TASK_PP(16'h1531E,4);
TASK_PP(16'h1531F,4);
TASK_PP(16'h15320,4);
TASK_PP(16'h15321,4);
TASK_PP(16'h15322,4);
TASK_PP(16'h15323,4);
TASK_PP(16'h15324,4);
TASK_PP(16'h15325,4);
TASK_PP(16'h15326,4);
TASK_PP(16'h15327,4);
TASK_PP(16'h15328,4);
TASK_PP(16'h15329,4);
TASK_PP(16'h1532A,4);
TASK_PP(16'h1532B,4);
TASK_PP(16'h1532C,4);
TASK_PP(16'h1532D,4);
TASK_PP(16'h1532E,4);
TASK_PP(16'h1532F,4);
TASK_PP(16'h15330,4);
TASK_PP(16'h15331,4);
TASK_PP(16'h15332,4);
TASK_PP(16'h15333,4);
TASK_PP(16'h15334,4);
TASK_PP(16'h15335,4);
TASK_PP(16'h15336,4);
TASK_PP(16'h15337,4);
TASK_PP(16'h15338,4);
TASK_PP(16'h15339,4);
TASK_PP(16'h1533A,4);
TASK_PP(16'h1533B,4);
TASK_PP(16'h1533C,4);
TASK_PP(16'h1533D,4);
TASK_PP(16'h1533E,4);
TASK_PP(16'h1533F,4);
TASK_PP(16'h15340,4);
TASK_PP(16'h15341,4);
TASK_PP(16'h15342,4);
TASK_PP(16'h15343,4);
TASK_PP(16'h15344,4);
TASK_PP(16'h15345,4);
TASK_PP(16'h15346,4);
TASK_PP(16'h15347,4);
TASK_PP(16'h15348,4);
TASK_PP(16'h15349,4);
TASK_PP(16'h1534A,4);
TASK_PP(16'h1534B,4);
TASK_PP(16'h1534C,4);
TASK_PP(16'h1534D,4);
TASK_PP(16'h1534E,4);
TASK_PP(16'h1534F,4);
TASK_PP(16'h15350,4);
TASK_PP(16'h15351,4);
TASK_PP(16'h15352,4);
TASK_PP(16'h15353,4);
TASK_PP(16'h15354,4);
TASK_PP(16'h15355,4);
TASK_PP(16'h15356,4);
TASK_PP(16'h15357,4);
TASK_PP(16'h15358,4);
TASK_PP(16'h15359,4);
TASK_PP(16'h1535A,4);
TASK_PP(16'h1535B,4);
TASK_PP(16'h1535C,4);
TASK_PP(16'h1535D,4);
TASK_PP(16'h1535E,4);
TASK_PP(16'h1535F,4);
TASK_PP(16'h15360,4);
TASK_PP(16'h15361,4);
TASK_PP(16'h15362,4);
TASK_PP(16'h15363,4);
TASK_PP(16'h15364,4);
TASK_PP(16'h15365,4);
TASK_PP(16'h15366,4);
TASK_PP(16'h15367,4);
TASK_PP(16'h15368,4);
TASK_PP(16'h15369,4);
TASK_PP(16'h1536A,4);
TASK_PP(16'h1536B,4);
TASK_PP(16'h1536C,4);
TASK_PP(16'h1536D,4);
TASK_PP(16'h1536E,4);
TASK_PP(16'h1536F,4);
TASK_PP(16'h15370,4);
TASK_PP(16'h15371,4);
TASK_PP(16'h15372,4);
TASK_PP(16'h15373,4);
TASK_PP(16'h15374,4);
TASK_PP(16'h15375,4);
TASK_PP(16'h15376,4);
TASK_PP(16'h15377,4);
TASK_PP(16'h15378,4);
TASK_PP(16'h15379,4);
TASK_PP(16'h1537A,4);
TASK_PP(16'h1537B,4);
TASK_PP(16'h1537C,4);
TASK_PP(16'h1537D,4);
TASK_PP(16'h1537E,4);
TASK_PP(16'h1537F,4);
TASK_PP(16'h15380,4);
TASK_PP(16'h15381,4);
TASK_PP(16'h15382,4);
TASK_PP(16'h15383,4);
TASK_PP(16'h15384,4);
TASK_PP(16'h15385,4);
TASK_PP(16'h15386,4);
TASK_PP(16'h15387,4);
TASK_PP(16'h15388,4);
TASK_PP(16'h15389,4);
TASK_PP(16'h1538A,4);
TASK_PP(16'h1538B,4);
TASK_PP(16'h1538C,4);
TASK_PP(16'h1538D,4);
TASK_PP(16'h1538E,4);
TASK_PP(16'h1538F,4);
TASK_PP(16'h15390,4);
TASK_PP(16'h15391,4);
TASK_PP(16'h15392,4);
TASK_PP(16'h15393,4);
TASK_PP(16'h15394,4);
TASK_PP(16'h15395,4);
TASK_PP(16'h15396,4);
TASK_PP(16'h15397,4);
TASK_PP(16'h15398,4);
TASK_PP(16'h15399,4);
TASK_PP(16'h1539A,4);
TASK_PP(16'h1539B,4);
TASK_PP(16'h1539C,4);
TASK_PP(16'h1539D,4);
TASK_PP(16'h1539E,4);
TASK_PP(16'h1539F,4);
TASK_PP(16'h153A0,4);
TASK_PP(16'h153A1,4);
TASK_PP(16'h153A2,4);
TASK_PP(16'h153A3,4);
TASK_PP(16'h153A4,4);
TASK_PP(16'h153A5,4);
TASK_PP(16'h153A6,4);
TASK_PP(16'h153A7,4);
TASK_PP(16'h153A8,4);
TASK_PP(16'h153A9,4);
TASK_PP(16'h153AA,4);
TASK_PP(16'h153AB,4);
TASK_PP(16'h153AC,4);
TASK_PP(16'h153AD,4);
TASK_PP(16'h153AE,4);
TASK_PP(16'h153AF,4);
TASK_PP(16'h153B0,4);
TASK_PP(16'h153B1,4);
TASK_PP(16'h153B2,4);
TASK_PP(16'h153B3,4);
TASK_PP(16'h153B4,4);
TASK_PP(16'h153B5,4);
TASK_PP(16'h153B6,4);
TASK_PP(16'h153B7,4);
TASK_PP(16'h153B8,4);
TASK_PP(16'h153B9,4);
TASK_PP(16'h153BA,4);
TASK_PP(16'h153BB,4);
TASK_PP(16'h153BC,4);
TASK_PP(16'h153BD,4);
TASK_PP(16'h153BE,4);
TASK_PP(16'h153BF,4);
TASK_PP(16'h153C0,4);
TASK_PP(16'h153C1,4);
TASK_PP(16'h153C2,4);
TASK_PP(16'h153C3,4);
TASK_PP(16'h153C4,4);
TASK_PP(16'h153C5,4);
TASK_PP(16'h153C6,4);
TASK_PP(16'h153C7,4);
TASK_PP(16'h153C8,4);
TASK_PP(16'h153C9,4);
TASK_PP(16'h153CA,4);
TASK_PP(16'h153CB,4);
TASK_PP(16'h153CC,4);
TASK_PP(16'h153CD,4);
TASK_PP(16'h153CE,4);
TASK_PP(16'h153CF,4);
TASK_PP(16'h153D0,4);
TASK_PP(16'h153D1,4);
TASK_PP(16'h153D2,4);
TASK_PP(16'h153D3,4);
TASK_PP(16'h153D4,4);
TASK_PP(16'h153D5,4);
TASK_PP(16'h153D6,4);
TASK_PP(16'h153D7,4);
TASK_PP(16'h153D8,4);
TASK_PP(16'h153D9,4);
TASK_PP(16'h153DA,4);
TASK_PP(16'h153DB,4);
TASK_PP(16'h153DC,4);
TASK_PP(16'h153DD,4);
TASK_PP(16'h153DE,4);
TASK_PP(16'h153DF,4);
TASK_PP(16'h153E0,4);
TASK_PP(16'h153E1,4);
TASK_PP(16'h153E2,4);
TASK_PP(16'h153E3,4);
TASK_PP(16'h153E4,4);
TASK_PP(16'h153E5,4);
TASK_PP(16'h153E6,4);
TASK_PP(16'h153E7,4);
TASK_PP(16'h153E8,4);
TASK_PP(16'h153E9,4);
TASK_PP(16'h153EA,4);
TASK_PP(16'h153EB,4);
TASK_PP(16'h153EC,4);
TASK_PP(16'h153ED,4);
TASK_PP(16'h153EE,4);
TASK_PP(16'h153EF,4);
TASK_PP(16'h153F0,4);
TASK_PP(16'h153F1,4);
TASK_PP(16'h153F2,4);
TASK_PP(16'h153F3,4);
TASK_PP(16'h153F4,4);
TASK_PP(16'h153F5,4);
TASK_PP(16'h153F6,4);
TASK_PP(16'h153F7,4);
TASK_PP(16'h153F8,4);
TASK_PP(16'h153F9,4);
TASK_PP(16'h153FA,4);
TASK_PP(16'h153FB,4);
TASK_PP(16'h153FC,4);
TASK_PP(16'h153FD,4);
TASK_PP(16'h153FE,4);
TASK_PP(16'h153FF,4);
TASK_PP(16'h15400,4);
TASK_PP(16'h15401,4);
TASK_PP(16'h15402,4);
TASK_PP(16'h15403,4);
TASK_PP(16'h15404,4);
TASK_PP(16'h15405,4);
TASK_PP(16'h15406,4);
TASK_PP(16'h15407,4);
TASK_PP(16'h15408,4);
TASK_PP(16'h15409,4);
TASK_PP(16'h1540A,4);
TASK_PP(16'h1540B,4);
TASK_PP(16'h1540C,4);
TASK_PP(16'h1540D,4);
TASK_PP(16'h1540E,4);
TASK_PP(16'h1540F,4);
TASK_PP(16'h15410,4);
TASK_PP(16'h15411,4);
TASK_PP(16'h15412,4);
TASK_PP(16'h15413,4);
TASK_PP(16'h15414,4);
TASK_PP(16'h15415,4);
TASK_PP(16'h15416,4);
TASK_PP(16'h15417,4);
TASK_PP(16'h15418,4);
TASK_PP(16'h15419,4);
TASK_PP(16'h1541A,4);
TASK_PP(16'h1541B,4);
TASK_PP(16'h1541C,4);
TASK_PP(16'h1541D,4);
TASK_PP(16'h1541E,4);
TASK_PP(16'h1541F,4);
TASK_PP(16'h15420,4);
TASK_PP(16'h15421,4);
TASK_PP(16'h15422,4);
TASK_PP(16'h15423,4);
TASK_PP(16'h15424,4);
TASK_PP(16'h15425,4);
TASK_PP(16'h15426,4);
TASK_PP(16'h15427,4);
TASK_PP(16'h15428,4);
TASK_PP(16'h15429,4);
TASK_PP(16'h1542A,4);
TASK_PP(16'h1542B,4);
TASK_PP(16'h1542C,4);
TASK_PP(16'h1542D,4);
TASK_PP(16'h1542E,4);
TASK_PP(16'h1542F,4);
TASK_PP(16'h15430,4);
TASK_PP(16'h15431,4);
TASK_PP(16'h15432,4);
TASK_PP(16'h15433,4);
TASK_PP(16'h15434,4);
TASK_PP(16'h15435,4);
TASK_PP(16'h15436,4);
TASK_PP(16'h15437,4);
TASK_PP(16'h15438,4);
TASK_PP(16'h15439,4);
TASK_PP(16'h1543A,4);
TASK_PP(16'h1543B,4);
TASK_PP(16'h1543C,4);
TASK_PP(16'h1543D,4);
TASK_PP(16'h1543E,4);
TASK_PP(16'h1543F,4);
TASK_PP(16'h15440,4);
TASK_PP(16'h15441,4);
TASK_PP(16'h15442,4);
TASK_PP(16'h15443,4);
TASK_PP(16'h15444,4);
TASK_PP(16'h15445,4);
TASK_PP(16'h15446,4);
TASK_PP(16'h15447,4);
TASK_PP(16'h15448,4);
TASK_PP(16'h15449,4);
TASK_PP(16'h1544A,4);
TASK_PP(16'h1544B,4);
TASK_PP(16'h1544C,4);
TASK_PP(16'h1544D,4);
TASK_PP(16'h1544E,4);
TASK_PP(16'h1544F,4);
TASK_PP(16'h15450,4);
TASK_PP(16'h15451,4);
TASK_PP(16'h15452,4);
TASK_PP(16'h15453,4);
TASK_PP(16'h15454,4);
TASK_PP(16'h15455,4);
TASK_PP(16'h15456,4);
TASK_PP(16'h15457,4);
TASK_PP(16'h15458,4);
TASK_PP(16'h15459,4);
TASK_PP(16'h1545A,4);
TASK_PP(16'h1545B,4);
TASK_PP(16'h1545C,4);
TASK_PP(16'h1545D,4);
TASK_PP(16'h1545E,4);
TASK_PP(16'h1545F,4);
TASK_PP(16'h15460,4);
TASK_PP(16'h15461,4);
TASK_PP(16'h15462,4);
TASK_PP(16'h15463,4);
TASK_PP(16'h15464,4);
TASK_PP(16'h15465,4);
TASK_PP(16'h15466,4);
TASK_PP(16'h15467,4);
TASK_PP(16'h15468,4);
TASK_PP(16'h15469,4);
TASK_PP(16'h1546A,4);
TASK_PP(16'h1546B,4);
TASK_PP(16'h1546C,4);
TASK_PP(16'h1546D,4);
TASK_PP(16'h1546E,4);
TASK_PP(16'h1546F,4);
TASK_PP(16'h15470,4);
TASK_PP(16'h15471,4);
TASK_PP(16'h15472,4);
TASK_PP(16'h15473,4);
TASK_PP(16'h15474,4);
TASK_PP(16'h15475,4);
TASK_PP(16'h15476,4);
TASK_PP(16'h15477,4);
TASK_PP(16'h15478,4);
TASK_PP(16'h15479,4);
TASK_PP(16'h1547A,4);
TASK_PP(16'h1547B,4);
TASK_PP(16'h1547C,4);
TASK_PP(16'h1547D,4);
TASK_PP(16'h1547E,4);
TASK_PP(16'h1547F,4);
TASK_PP(16'h15480,4);
TASK_PP(16'h15481,4);
TASK_PP(16'h15482,4);
TASK_PP(16'h15483,4);
TASK_PP(16'h15484,4);
TASK_PP(16'h15485,4);
TASK_PP(16'h15486,4);
TASK_PP(16'h15487,4);
TASK_PP(16'h15488,4);
TASK_PP(16'h15489,4);
TASK_PP(16'h1548A,4);
TASK_PP(16'h1548B,4);
TASK_PP(16'h1548C,4);
TASK_PP(16'h1548D,4);
TASK_PP(16'h1548E,4);
TASK_PP(16'h1548F,4);
TASK_PP(16'h15490,4);
TASK_PP(16'h15491,4);
TASK_PP(16'h15492,4);
TASK_PP(16'h15493,4);
TASK_PP(16'h15494,4);
TASK_PP(16'h15495,4);
TASK_PP(16'h15496,4);
TASK_PP(16'h15497,4);
TASK_PP(16'h15498,4);
TASK_PP(16'h15499,4);
TASK_PP(16'h1549A,4);
TASK_PP(16'h1549B,4);
TASK_PP(16'h1549C,4);
TASK_PP(16'h1549D,4);
TASK_PP(16'h1549E,4);
TASK_PP(16'h1549F,4);
TASK_PP(16'h154A0,4);
TASK_PP(16'h154A1,4);
TASK_PP(16'h154A2,4);
TASK_PP(16'h154A3,4);
TASK_PP(16'h154A4,4);
TASK_PP(16'h154A5,4);
TASK_PP(16'h154A6,4);
TASK_PP(16'h154A7,4);
TASK_PP(16'h154A8,4);
TASK_PP(16'h154A9,4);
TASK_PP(16'h154AA,4);
TASK_PP(16'h154AB,4);
TASK_PP(16'h154AC,4);
TASK_PP(16'h154AD,4);
TASK_PP(16'h154AE,4);
TASK_PP(16'h154AF,4);
TASK_PP(16'h154B0,4);
TASK_PP(16'h154B1,4);
TASK_PP(16'h154B2,4);
TASK_PP(16'h154B3,4);
TASK_PP(16'h154B4,4);
TASK_PP(16'h154B5,4);
TASK_PP(16'h154B6,4);
TASK_PP(16'h154B7,4);
TASK_PP(16'h154B8,4);
TASK_PP(16'h154B9,4);
TASK_PP(16'h154BA,4);
TASK_PP(16'h154BB,4);
TASK_PP(16'h154BC,4);
TASK_PP(16'h154BD,4);
TASK_PP(16'h154BE,4);
TASK_PP(16'h154BF,4);
TASK_PP(16'h154C0,4);
TASK_PP(16'h154C1,4);
TASK_PP(16'h154C2,4);
TASK_PP(16'h154C3,4);
TASK_PP(16'h154C4,4);
TASK_PP(16'h154C5,4);
TASK_PP(16'h154C6,4);
TASK_PP(16'h154C7,4);
TASK_PP(16'h154C8,4);
TASK_PP(16'h154C9,4);
TASK_PP(16'h154CA,4);
TASK_PP(16'h154CB,4);
TASK_PP(16'h154CC,4);
TASK_PP(16'h154CD,4);
TASK_PP(16'h154CE,4);
TASK_PP(16'h154CF,4);
TASK_PP(16'h154D0,4);
TASK_PP(16'h154D1,4);
TASK_PP(16'h154D2,4);
TASK_PP(16'h154D3,4);
TASK_PP(16'h154D4,4);
TASK_PP(16'h154D5,4);
TASK_PP(16'h154D6,4);
TASK_PP(16'h154D7,4);
TASK_PP(16'h154D8,4);
TASK_PP(16'h154D9,4);
TASK_PP(16'h154DA,4);
TASK_PP(16'h154DB,4);
TASK_PP(16'h154DC,4);
TASK_PP(16'h154DD,4);
TASK_PP(16'h154DE,4);
TASK_PP(16'h154DF,4);
TASK_PP(16'h154E0,4);
TASK_PP(16'h154E1,4);
TASK_PP(16'h154E2,4);
TASK_PP(16'h154E3,4);
TASK_PP(16'h154E4,4);
TASK_PP(16'h154E5,4);
TASK_PP(16'h154E6,4);
TASK_PP(16'h154E7,4);
TASK_PP(16'h154E8,4);
TASK_PP(16'h154E9,4);
TASK_PP(16'h154EA,4);
TASK_PP(16'h154EB,4);
TASK_PP(16'h154EC,4);
TASK_PP(16'h154ED,4);
TASK_PP(16'h154EE,4);
TASK_PP(16'h154EF,4);
TASK_PP(16'h154F0,4);
TASK_PP(16'h154F1,4);
TASK_PP(16'h154F2,4);
TASK_PP(16'h154F3,4);
TASK_PP(16'h154F4,4);
TASK_PP(16'h154F5,4);
TASK_PP(16'h154F6,4);
TASK_PP(16'h154F7,4);
TASK_PP(16'h154F8,4);
TASK_PP(16'h154F9,4);
TASK_PP(16'h154FA,4);
TASK_PP(16'h154FB,4);
TASK_PP(16'h154FC,4);
TASK_PP(16'h154FD,4);
TASK_PP(16'h154FE,4);
TASK_PP(16'h154FF,4);
TASK_PP(16'h15500,4);
TASK_PP(16'h15501,4);
TASK_PP(16'h15502,4);
TASK_PP(16'h15503,4);
TASK_PP(16'h15504,4);
TASK_PP(16'h15505,4);
TASK_PP(16'h15506,4);
TASK_PP(16'h15507,4);
TASK_PP(16'h15508,4);
TASK_PP(16'h15509,4);
TASK_PP(16'h1550A,4);
TASK_PP(16'h1550B,4);
TASK_PP(16'h1550C,4);
TASK_PP(16'h1550D,4);
TASK_PP(16'h1550E,4);
TASK_PP(16'h1550F,4);
TASK_PP(16'h15510,4);
TASK_PP(16'h15511,4);
TASK_PP(16'h15512,4);
TASK_PP(16'h15513,4);
TASK_PP(16'h15514,4);
TASK_PP(16'h15515,4);
TASK_PP(16'h15516,4);
TASK_PP(16'h15517,4);
TASK_PP(16'h15518,4);
TASK_PP(16'h15519,4);
TASK_PP(16'h1551A,4);
TASK_PP(16'h1551B,4);
TASK_PP(16'h1551C,4);
TASK_PP(16'h1551D,4);
TASK_PP(16'h1551E,4);
TASK_PP(16'h1551F,4);
TASK_PP(16'h15520,4);
TASK_PP(16'h15521,4);
TASK_PP(16'h15522,4);
TASK_PP(16'h15523,4);
TASK_PP(16'h15524,4);
TASK_PP(16'h15525,4);
TASK_PP(16'h15526,4);
TASK_PP(16'h15527,4);
TASK_PP(16'h15528,4);
TASK_PP(16'h15529,4);
TASK_PP(16'h1552A,4);
TASK_PP(16'h1552B,4);
TASK_PP(16'h1552C,4);
TASK_PP(16'h1552D,4);
TASK_PP(16'h1552E,4);
TASK_PP(16'h1552F,4);
TASK_PP(16'h15530,4);
TASK_PP(16'h15531,4);
TASK_PP(16'h15532,4);
TASK_PP(16'h15533,4);
TASK_PP(16'h15534,4);
TASK_PP(16'h15535,4);
TASK_PP(16'h15536,4);
TASK_PP(16'h15537,4);
TASK_PP(16'h15538,4);
TASK_PP(16'h15539,4);
TASK_PP(16'h1553A,4);
TASK_PP(16'h1553B,4);
TASK_PP(16'h1553C,4);
TASK_PP(16'h1553D,4);
TASK_PP(16'h1553E,4);
TASK_PP(16'h1553F,4);
TASK_PP(16'h15540,4);
TASK_PP(16'h15541,4);
TASK_PP(16'h15542,4);
TASK_PP(16'h15543,4);
TASK_PP(16'h15544,4);
TASK_PP(16'h15545,4);
TASK_PP(16'h15546,4);
TASK_PP(16'h15547,4);
TASK_PP(16'h15548,4);
TASK_PP(16'h15549,4);
TASK_PP(16'h1554A,4);
TASK_PP(16'h1554B,4);
TASK_PP(16'h1554C,4);
TASK_PP(16'h1554D,4);
TASK_PP(16'h1554E,4);
TASK_PP(16'h1554F,4);
TASK_PP(16'h15550,4);
TASK_PP(16'h15551,4);
TASK_PP(16'h15552,4);
TASK_PP(16'h15553,4);
TASK_PP(16'h15554,4);
TASK_PP(16'h15555,4);
TASK_PP(16'h15556,4);
TASK_PP(16'h15557,4);
TASK_PP(16'h15558,4);
TASK_PP(16'h15559,4);
TASK_PP(16'h1555A,4);
TASK_PP(16'h1555B,4);
TASK_PP(16'h1555C,4);
TASK_PP(16'h1555D,4);
TASK_PP(16'h1555E,4);
TASK_PP(16'h1555F,4);
TASK_PP(16'h15560,4);
TASK_PP(16'h15561,4);
TASK_PP(16'h15562,4);
TASK_PP(16'h15563,4);
TASK_PP(16'h15564,4);
TASK_PP(16'h15565,4);
TASK_PP(16'h15566,4);
TASK_PP(16'h15567,4);
TASK_PP(16'h15568,4);
TASK_PP(16'h15569,4);
TASK_PP(16'h1556A,4);
TASK_PP(16'h1556B,4);
TASK_PP(16'h1556C,4);
TASK_PP(16'h1556D,4);
TASK_PP(16'h1556E,4);
TASK_PP(16'h1556F,4);
TASK_PP(16'h15570,4);
TASK_PP(16'h15571,4);
TASK_PP(16'h15572,4);
TASK_PP(16'h15573,4);
TASK_PP(16'h15574,4);
TASK_PP(16'h15575,4);
TASK_PP(16'h15576,4);
TASK_PP(16'h15577,4);
TASK_PP(16'h15578,4);
TASK_PP(16'h15579,4);
TASK_PP(16'h1557A,4);
TASK_PP(16'h1557B,4);
TASK_PP(16'h1557C,4);
TASK_PP(16'h1557D,4);
TASK_PP(16'h1557E,4);
TASK_PP(16'h1557F,4);
TASK_PP(16'h15580,4);
TASK_PP(16'h15581,4);
TASK_PP(16'h15582,4);
TASK_PP(16'h15583,4);
TASK_PP(16'h15584,4);
TASK_PP(16'h15585,4);
TASK_PP(16'h15586,4);
TASK_PP(16'h15587,4);
TASK_PP(16'h15588,4);
TASK_PP(16'h15589,4);
TASK_PP(16'h1558A,4);
TASK_PP(16'h1558B,4);
TASK_PP(16'h1558C,4);
TASK_PP(16'h1558D,4);
TASK_PP(16'h1558E,4);
TASK_PP(16'h1558F,4);
TASK_PP(16'h15590,4);
TASK_PP(16'h15591,4);
TASK_PP(16'h15592,4);
TASK_PP(16'h15593,4);
TASK_PP(16'h15594,4);
TASK_PP(16'h15595,4);
TASK_PP(16'h15596,4);
TASK_PP(16'h15597,4);
TASK_PP(16'h15598,4);
TASK_PP(16'h15599,4);
TASK_PP(16'h1559A,4);
TASK_PP(16'h1559B,4);
TASK_PP(16'h1559C,4);
TASK_PP(16'h1559D,4);
TASK_PP(16'h1559E,4);
TASK_PP(16'h1559F,4);
TASK_PP(16'h155A0,4);
TASK_PP(16'h155A1,4);
TASK_PP(16'h155A2,4);
TASK_PP(16'h155A3,4);
TASK_PP(16'h155A4,4);
TASK_PP(16'h155A5,4);
TASK_PP(16'h155A6,4);
TASK_PP(16'h155A7,4);
TASK_PP(16'h155A8,4);
TASK_PP(16'h155A9,4);
TASK_PP(16'h155AA,4);
TASK_PP(16'h155AB,4);
TASK_PP(16'h155AC,4);
TASK_PP(16'h155AD,4);
TASK_PP(16'h155AE,4);
TASK_PP(16'h155AF,4);
TASK_PP(16'h155B0,4);
TASK_PP(16'h155B1,4);
TASK_PP(16'h155B2,4);
TASK_PP(16'h155B3,4);
TASK_PP(16'h155B4,4);
TASK_PP(16'h155B5,4);
TASK_PP(16'h155B6,4);
TASK_PP(16'h155B7,4);
TASK_PP(16'h155B8,4);
TASK_PP(16'h155B9,4);
TASK_PP(16'h155BA,4);
TASK_PP(16'h155BB,4);
TASK_PP(16'h155BC,4);
TASK_PP(16'h155BD,4);
TASK_PP(16'h155BE,4);
TASK_PP(16'h155BF,4);
TASK_PP(16'h155C0,4);
TASK_PP(16'h155C1,4);
TASK_PP(16'h155C2,4);
TASK_PP(16'h155C3,4);
TASK_PP(16'h155C4,4);
TASK_PP(16'h155C5,4);
TASK_PP(16'h155C6,4);
TASK_PP(16'h155C7,4);
TASK_PP(16'h155C8,4);
TASK_PP(16'h155C9,4);
TASK_PP(16'h155CA,4);
TASK_PP(16'h155CB,4);
TASK_PP(16'h155CC,4);
TASK_PP(16'h155CD,4);
TASK_PP(16'h155CE,4);
TASK_PP(16'h155CF,4);
TASK_PP(16'h155D0,4);
TASK_PP(16'h155D1,4);
TASK_PP(16'h155D2,4);
TASK_PP(16'h155D3,4);
TASK_PP(16'h155D4,4);
TASK_PP(16'h155D5,4);
TASK_PP(16'h155D6,4);
TASK_PP(16'h155D7,4);
TASK_PP(16'h155D8,4);
TASK_PP(16'h155D9,4);
TASK_PP(16'h155DA,4);
TASK_PP(16'h155DB,4);
TASK_PP(16'h155DC,4);
TASK_PP(16'h155DD,4);
TASK_PP(16'h155DE,4);
TASK_PP(16'h155DF,4);
TASK_PP(16'h155E0,4);
TASK_PP(16'h155E1,4);
TASK_PP(16'h155E2,4);
TASK_PP(16'h155E3,4);
TASK_PP(16'h155E4,4);
TASK_PP(16'h155E5,4);
TASK_PP(16'h155E6,4);
TASK_PP(16'h155E7,4);
TASK_PP(16'h155E8,4);
TASK_PP(16'h155E9,4);
TASK_PP(16'h155EA,4);
TASK_PP(16'h155EB,4);
TASK_PP(16'h155EC,4);
TASK_PP(16'h155ED,4);
TASK_PP(16'h155EE,4);
TASK_PP(16'h155EF,4);
TASK_PP(16'h155F0,4);
TASK_PP(16'h155F1,4);
TASK_PP(16'h155F2,4);
TASK_PP(16'h155F3,4);
TASK_PP(16'h155F4,4);
TASK_PP(16'h155F5,4);
TASK_PP(16'h155F6,4);
TASK_PP(16'h155F7,4);
TASK_PP(16'h155F8,4);
TASK_PP(16'h155F9,4);
TASK_PP(16'h155FA,4);
TASK_PP(16'h155FB,4);
TASK_PP(16'h155FC,4);
TASK_PP(16'h155FD,4);
TASK_PP(16'h155FE,4);
TASK_PP(16'h155FF,4);
TASK_PP(16'h15600,4);
TASK_PP(16'h15601,4);
TASK_PP(16'h15602,4);
TASK_PP(16'h15603,4);
TASK_PP(16'h15604,4);
TASK_PP(16'h15605,4);
TASK_PP(16'h15606,4);
TASK_PP(16'h15607,4);
TASK_PP(16'h15608,4);
TASK_PP(16'h15609,4);
TASK_PP(16'h1560A,4);
TASK_PP(16'h1560B,4);
TASK_PP(16'h1560C,4);
TASK_PP(16'h1560D,4);
TASK_PP(16'h1560E,4);
TASK_PP(16'h1560F,4);
TASK_PP(16'h15610,4);
TASK_PP(16'h15611,4);
TASK_PP(16'h15612,4);
TASK_PP(16'h15613,4);
TASK_PP(16'h15614,4);
TASK_PP(16'h15615,4);
TASK_PP(16'h15616,4);
TASK_PP(16'h15617,4);
TASK_PP(16'h15618,4);
TASK_PP(16'h15619,4);
TASK_PP(16'h1561A,4);
TASK_PP(16'h1561B,4);
TASK_PP(16'h1561C,4);
TASK_PP(16'h1561D,4);
TASK_PP(16'h1561E,4);
TASK_PP(16'h1561F,4);
TASK_PP(16'h15620,4);
TASK_PP(16'h15621,4);
TASK_PP(16'h15622,4);
TASK_PP(16'h15623,4);
TASK_PP(16'h15624,4);
TASK_PP(16'h15625,4);
TASK_PP(16'h15626,4);
TASK_PP(16'h15627,4);
TASK_PP(16'h15628,4);
TASK_PP(16'h15629,4);
TASK_PP(16'h1562A,4);
TASK_PP(16'h1562B,4);
TASK_PP(16'h1562C,4);
TASK_PP(16'h1562D,4);
TASK_PP(16'h1562E,4);
TASK_PP(16'h1562F,4);
TASK_PP(16'h15630,4);
TASK_PP(16'h15631,4);
TASK_PP(16'h15632,4);
TASK_PP(16'h15633,4);
TASK_PP(16'h15634,4);
TASK_PP(16'h15635,4);
TASK_PP(16'h15636,4);
TASK_PP(16'h15637,4);
TASK_PP(16'h15638,4);
TASK_PP(16'h15639,4);
TASK_PP(16'h1563A,4);
TASK_PP(16'h1563B,4);
TASK_PP(16'h1563C,4);
TASK_PP(16'h1563D,4);
TASK_PP(16'h1563E,4);
TASK_PP(16'h1563F,4);
TASK_PP(16'h15640,4);
TASK_PP(16'h15641,4);
TASK_PP(16'h15642,4);
TASK_PP(16'h15643,4);
TASK_PP(16'h15644,4);
TASK_PP(16'h15645,4);
TASK_PP(16'h15646,4);
TASK_PP(16'h15647,4);
TASK_PP(16'h15648,4);
TASK_PP(16'h15649,4);
TASK_PP(16'h1564A,4);
TASK_PP(16'h1564B,4);
TASK_PP(16'h1564C,4);
TASK_PP(16'h1564D,4);
TASK_PP(16'h1564E,4);
TASK_PP(16'h1564F,4);
TASK_PP(16'h15650,4);
TASK_PP(16'h15651,4);
TASK_PP(16'h15652,4);
TASK_PP(16'h15653,4);
TASK_PP(16'h15654,4);
TASK_PP(16'h15655,4);
TASK_PP(16'h15656,4);
TASK_PP(16'h15657,4);
TASK_PP(16'h15658,4);
TASK_PP(16'h15659,4);
TASK_PP(16'h1565A,4);
TASK_PP(16'h1565B,4);
TASK_PP(16'h1565C,4);
TASK_PP(16'h1565D,4);
TASK_PP(16'h1565E,4);
TASK_PP(16'h1565F,4);
TASK_PP(16'h15660,4);
TASK_PP(16'h15661,4);
TASK_PP(16'h15662,4);
TASK_PP(16'h15663,4);
TASK_PP(16'h15664,4);
TASK_PP(16'h15665,4);
TASK_PP(16'h15666,4);
TASK_PP(16'h15667,4);
TASK_PP(16'h15668,4);
TASK_PP(16'h15669,4);
TASK_PP(16'h1566A,4);
TASK_PP(16'h1566B,4);
TASK_PP(16'h1566C,4);
TASK_PP(16'h1566D,4);
TASK_PP(16'h1566E,4);
TASK_PP(16'h1566F,4);
TASK_PP(16'h15670,4);
TASK_PP(16'h15671,4);
TASK_PP(16'h15672,4);
TASK_PP(16'h15673,4);
TASK_PP(16'h15674,4);
TASK_PP(16'h15675,4);
TASK_PP(16'h15676,4);
TASK_PP(16'h15677,4);
TASK_PP(16'h15678,4);
TASK_PP(16'h15679,4);
TASK_PP(16'h1567A,4);
TASK_PP(16'h1567B,4);
TASK_PP(16'h1567C,4);
TASK_PP(16'h1567D,4);
TASK_PP(16'h1567E,4);
TASK_PP(16'h1567F,4);
TASK_PP(16'h15680,4);
TASK_PP(16'h15681,4);
TASK_PP(16'h15682,4);
TASK_PP(16'h15683,4);
TASK_PP(16'h15684,4);
TASK_PP(16'h15685,4);
TASK_PP(16'h15686,4);
TASK_PP(16'h15687,4);
TASK_PP(16'h15688,4);
TASK_PP(16'h15689,4);
TASK_PP(16'h1568A,4);
TASK_PP(16'h1568B,4);
TASK_PP(16'h1568C,4);
TASK_PP(16'h1568D,4);
TASK_PP(16'h1568E,4);
TASK_PP(16'h1568F,4);
TASK_PP(16'h15690,4);
TASK_PP(16'h15691,4);
TASK_PP(16'h15692,4);
TASK_PP(16'h15693,4);
TASK_PP(16'h15694,4);
TASK_PP(16'h15695,4);
TASK_PP(16'h15696,4);
TASK_PP(16'h15697,4);
TASK_PP(16'h15698,4);
TASK_PP(16'h15699,4);
TASK_PP(16'h1569A,4);
TASK_PP(16'h1569B,4);
TASK_PP(16'h1569C,4);
TASK_PP(16'h1569D,4);
TASK_PP(16'h1569E,4);
TASK_PP(16'h1569F,4);
TASK_PP(16'h156A0,4);
TASK_PP(16'h156A1,4);
TASK_PP(16'h156A2,4);
TASK_PP(16'h156A3,4);
TASK_PP(16'h156A4,4);
TASK_PP(16'h156A5,4);
TASK_PP(16'h156A6,4);
TASK_PP(16'h156A7,4);
TASK_PP(16'h156A8,4);
TASK_PP(16'h156A9,4);
TASK_PP(16'h156AA,4);
TASK_PP(16'h156AB,4);
TASK_PP(16'h156AC,4);
TASK_PP(16'h156AD,4);
TASK_PP(16'h156AE,4);
TASK_PP(16'h156AF,4);
TASK_PP(16'h156B0,4);
TASK_PP(16'h156B1,4);
TASK_PP(16'h156B2,4);
TASK_PP(16'h156B3,4);
TASK_PP(16'h156B4,4);
TASK_PP(16'h156B5,4);
TASK_PP(16'h156B6,4);
TASK_PP(16'h156B7,4);
TASK_PP(16'h156B8,4);
TASK_PP(16'h156B9,4);
TASK_PP(16'h156BA,4);
TASK_PP(16'h156BB,4);
TASK_PP(16'h156BC,4);
TASK_PP(16'h156BD,4);
TASK_PP(16'h156BE,4);
TASK_PP(16'h156BF,4);
TASK_PP(16'h156C0,4);
TASK_PP(16'h156C1,4);
TASK_PP(16'h156C2,4);
TASK_PP(16'h156C3,4);
TASK_PP(16'h156C4,4);
TASK_PP(16'h156C5,4);
TASK_PP(16'h156C6,4);
TASK_PP(16'h156C7,4);
TASK_PP(16'h156C8,4);
TASK_PP(16'h156C9,4);
TASK_PP(16'h156CA,4);
TASK_PP(16'h156CB,4);
TASK_PP(16'h156CC,4);
TASK_PP(16'h156CD,4);
TASK_PP(16'h156CE,4);
TASK_PP(16'h156CF,4);
TASK_PP(16'h156D0,4);
TASK_PP(16'h156D1,4);
TASK_PP(16'h156D2,4);
TASK_PP(16'h156D3,4);
TASK_PP(16'h156D4,4);
TASK_PP(16'h156D5,4);
TASK_PP(16'h156D6,4);
TASK_PP(16'h156D7,4);
TASK_PP(16'h156D8,4);
TASK_PP(16'h156D9,4);
TASK_PP(16'h156DA,4);
TASK_PP(16'h156DB,4);
TASK_PP(16'h156DC,4);
TASK_PP(16'h156DD,4);
TASK_PP(16'h156DE,4);
TASK_PP(16'h156DF,4);
TASK_PP(16'h156E0,4);
TASK_PP(16'h156E1,4);
TASK_PP(16'h156E2,4);
TASK_PP(16'h156E3,4);
TASK_PP(16'h156E4,4);
TASK_PP(16'h156E5,4);
TASK_PP(16'h156E6,4);
TASK_PP(16'h156E7,4);
TASK_PP(16'h156E8,4);
TASK_PP(16'h156E9,4);
TASK_PP(16'h156EA,4);
TASK_PP(16'h156EB,4);
TASK_PP(16'h156EC,4);
TASK_PP(16'h156ED,4);
TASK_PP(16'h156EE,4);
TASK_PP(16'h156EF,4);
TASK_PP(16'h156F0,4);
TASK_PP(16'h156F1,4);
TASK_PP(16'h156F2,4);
TASK_PP(16'h156F3,4);
TASK_PP(16'h156F4,4);
TASK_PP(16'h156F5,4);
TASK_PP(16'h156F6,4);
TASK_PP(16'h156F7,4);
TASK_PP(16'h156F8,4);
TASK_PP(16'h156F9,4);
TASK_PP(16'h156FA,4);
TASK_PP(16'h156FB,4);
TASK_PP(16'h156FC,4);
TASK_PP(16'h156FD,4);
TASK_PP(16'h156FE,4);
TASK_PP(16'h156FF,4);
TASK_PP(16'h15700,4);
TASK_PP(16'h15701,4);
TASK_PP(16'h15702,4);
TASK_PP(16'h15703,4);
TASK_PP(16'h15704,4);
TASK_PP(16'h15705,4);
TASK_PP(16'h15706,4);
TASK_PP(16'h15707,4);
TASK_PP(16'h15708,4);
TASK_PP(16'h15709,4);
TASK_PP(16'h1570A,4);
TASK_PP(16'h1570B,4);
TASK_PP(16'h1570C,4);
TASK_PP(16'h1570D,4);
TASK_PP(16'h1570E,4);
TASK_PP(16'h1570F,4);
TASK_PP(16'h15710,4);
TASK_PP(16'h15711,4);
TASK_PP(16'h15712,4);
TASK_PP(16'h15713,4);
TASK_PP(16'h15714,4);
TASK_PP(16'h15715,4);
TASK_PP(16'h15716,4);
TASK_PP(16'h15717,4);
TASK_PP(16'h15718,4);
TASK_PP(16'h15719,4);
TASK_PP(16'h1571A,4);
TASK_PP(16'h1571B,4);
TASK_PP(16'h1571C,4);
TASK_PP(16'h1571D,4);
TASK_PP(16'h1571E,4);
TASK_PP(16'h1571F,4);
TASK_PP(16'h15720,4);
TASK_PP(16'h15721,4);
TASK_PP(16'h15722,4);
TASK_PP(16'h15723,4);
TASK_PP(16'h15724,4);
TASK_PP(16'h15725,4);
TASK_PP(16'h15726,4);
TASK_PP(16'h15727,4);
TASK_PP(16'h15728,4);
TASK_PP(16'h15729,4);
TASK_PP(16'h1572A,4);
TASK_PP(16'h1572B,4);
TASK_PP(16'h1572C,4);
TASK_PP(16'h1572D,4);
TASK_PP(16'h1572E,4);
TASK_PP(16'h1572F,4);
TASK_PP(16'h15730,4);
TASK_PP(16'h15731,4);
TASK_PP(16'h15732,4);
TASK_PP(16'h15733,4);
TASK_PP(16'h15734,4);
TASK_PP(16'h15735,4);
TASK_PP(16'h15736,4);
TASK_PP(16'h15737,4);
TASK_PP(16'h15738,4);
TASK_PP(16'h15739,4);
TASK_PP(16'h1573A,4);
TASK_PP(16'h1573B,4);
TASK_PP(16'h1573C,4);
TASK_PP(16'h1573D,4);
TASK_PP(16'h1573E,4);
TASK_PP(16'h1573F,4);
TASK_PP(16'h15740,4);
TASK_PP(16'h15741,4);
TASK_PP(16'h15742,4);
TASK_PP(16'h15743,4);
TASK_PP(16'h15744,4);
TASK_PP(16'h15745,4);
TASK_PP(16'h15746,4);
TASK_PP(16'h15747,4);
TASK_PP(16'h15748,4);
TASK_PP(16'h15749,4);
TASK_PP(16'h1574A,4);
TASK_PP(16'h1574B,4);
TASK_PP(16'h1574C,4);
TASK_PP(16'h1574D,4);
TASK_PP(16'h1574E,4);
TASK_PP(16'h1574F,4);
TASK_PP(16'h15750,4);
TASK_PP(16'h15751,4);
TASK_PP(16'h15752,4);
TASK_PP(16'h15753,4);
TASK_PP(16'h15754,4);
TASK_PP(16'h15755,4);
TASK_PP(16'h15756,4);
TASK_PP(16'h15757,4);
TASK_PP(16'h15758,4);
TASK_PP(16'h15759,4);
TASK_PP(16'h1575A,4);
TASK_PP(16'h1575B,4);
TASK_PP(16'h1575C,4);
TASK_PP(16'h1575D,4);
TASK_PP(16'h1575E,4);
TASK_PP(16'h1575F,4);
TASK_PP(16'h15760,4);
TASK_PP(16'h15761,4);
TASK_PP(16'h15762,4);
TASK_PP(16'h15763,4);
TASK_PP(16'h15764,4);
TASK_PP(16'h15765,4);
TASK_PP(16'h15766,4);
TASK_PP(16'h15767,4);
TASK_PP(16'h15768,4);
TASK_PP(16'h15769,4);
TASK_PP(16'h1576A,4);
TASK_PP(16'h1576B,4);
TASK_PP(16'h1576C,4);
TASK_PP(16'h1576D,4);
TASK_PP(16'h1576E,4);
TASK_PP(16'h1576F,4);
TASK_PP(16'h15770,4);
TASK_PP(16'h15771,4);
TASK_PP(16'h15772,4);
TASK_PP(16'h15773,4);
TASK_PP(16'h15774,4);
TASK_PP(16'h15775,4);
TASK_PP(16'h15776,4);
TASK_PP(16'h15777,4);
TASK_PP(16'h15778,4);
TASK_PP(16'h15779,4);
TASK_PP(16'h1577A,4);
TASK_PP(16'h1577B,4);
TASK_PP(16'h1577C,4);
TASK_PP(16'h1577D,4);
TASK_PP(16'h1577E,4);
TASK_PP(16'h1577F,4);
TASK_PP(16'h15780,4);
TASK_PP(16'h15781,4);
TASK_PP(16'h15782,4);
TASK_PP(16'h15783,4);
TASK_PP(16'h15784,4);
TASK_PP(16'h15785,4);
TASK_PP(16'h15786,4);
TASK_PP(16'h15787,4);
TASK_PP(16'h15788,4);
TASK_PP(16'h15789,4);
TASK_PP(16'h1578A,4);
TASK_PP(16'h1578B,4);
TASK_PP(16'h1578C,4);
TASK_PP(16'h1578D,4);
TASK_PP(16'h1578E,4);
TASK_PP(16'h1578F,4);
TASK_PP(16'h15790,4);
TASK_PP(16'h15791,4);
TASK_PP(16'h15792,4);
TASK_PP(16'h15793,4);
TASK_PP(16'h15794,4);
TASK_PP(16'h15795,4);
TASK_PP(16'h15796,4);
TASK_PP(16'h15797,4);
TASK_PP(16'h15798,4);
TASK_PP(16'h15799,4);
TASK_PP(16'h1579A,4);
TASK_PP(16'h1579B,4);
TASK_PP(16'h1579C,4);
TASK_PP(16'h1579D,4);
TASK_PP(16'h1579E,4);
TASK_PP(16'h1579F,4);
TASK_PP(16'h157A0,4);
TASK_PP(16'h157A1,4);
TASK_PP(16'h157A2,4);
TASK_PP(16'h157A3,4);
TASK_PP(16'h157A4,4);
TASK_PP(16'h157A5,4);
TASK_PP(16'h157A6,4);
TASK_PP(16'h157A7,4);
TASK_PP(16'h157A8,4);
TASK_PP(16'h157A9,4);
TASK_PP(16'h157AA,4);
TASK_PP(16'h157AB,4);
TASK_PP(16'h157AC,4);
TASK_PP(16'h157AD,4);
TASK_PP(16'h157AE,4);
TASK_PP(16'h157AF,4);
TASK_PP(16'h157B0,4);
TASK_PP(16'h157B1,4);
TASK_PP(16'h157B2,4);
TASK_PP(16'h157B3,4);
TASK_PP(16'h157B4,4);
TASK_PP(16'h157B5,4);
TASK_PP(16'h157B6,4);
TASK_PP(16'h157B7,4);
TASK_PP(16'h157B8,4);
TASK_PP(16'h157B9,4);
TASK_PP(16'h157BA,4);
TASK_PP(16'h157BB,4);
TASK_PP(16'h157BC,4);
TASK_PP(16'h157BD,4);
TASK_PP(16'h157BE,4);
TASK_PP(16'h157BF,4);
TASK_PP(16'h157C0,4);
TASK_PP(16'h157C1,4);
TASK_PP(16'h157C2,4);
TASK_PP(16'h157C3,4);
TASK_PP(16'h157C4,4);
TASK_PP(16'h157C5,4);
TASK_PP(16'h157C6,4);
TASK_PP(16'h157C7,4);
TASK_PP(16'h157C8,4);
TASK_PP(16'h157C9,4);
TASK_PP(16'h157CA,4);
TASK_PP(16'h157CB,4);
TASK_PP(16'h157CC,4);
TASK_PP(16'h157CD,4);
TASK_PP(16'h157CE,4);
TASK_PP(16'h157CF,4);
TASK_PP(16'h157D0,4);
TASK_PP(16'h157D1,4);
TASK_PP(16'h157D2,4);
TASK_PP(16'h157D3,4);
TASK_PP(16'h157D4,4);
TASK_PP(16'h157D5,4);
TASK_PP(16'h157D6,4);
TASK_PP(16'h157D7,4);
TASK_PP(16'h157D8,4);
TASK_PP(16'h157D9,4);
TASK_PP(16'h157DA,4);
TASK_PP(16'h157DB,4);
TASK_PP(16'h157DC,4);
TASK_PP(16'h157DD,4);
TASK_PP(16'h157DE,4);
TASK_PP(16'h157DF,4);
TASK_PP(16'h157E0,4);
TASK_PP(16'h157E1,4);
TASK_PP(16'h157E2,4);
TASK_PP(16'h157E3,4);
TASK_PP(16'h157E4,4);
TASK_PP(16'h157E5,4);
TASK_PP(16'h157E6,4);
TASK_PP(16'h157E7,4);
TASK_PP(16'h157E8,4);
TASK_PP(16'h157E9,4);
TASK_PP(16'h157EA,4);
TASK_PP(16'h157EB,4);
TASK_PP(16'h157EC,4);
TASK_PP(16'h157ED,4);
TASK_PP(16'h157EE,4);
TASK_PP(16'h157EF,4);
TASK_PP(16'h157F0,4);
TASK_PP(16'h157F1,4);
TASK_PP(16'h157F2,4);
TASK_PP(16'h157F3,4);
TASK_PP(16'h157F4,4);
TASK_PP(16'h157F5,4);
TASK_PP(16'h157F6,4);
TASK_PP(16'h157F7,4);
TASK_PP(16'h157F8,4);
TASK_PP(16'h157F9,4);
TASK_PP(16'h157FA,4);
TASK_PP(16'h157FB,4);
TASK_PP(16'h157FC,4);
TASK_PP(16'h157FD,4);
TASK_PP(16'h157FE,4);
TASK_PP(16'h157FF,4);
TASK_PP(16'h15800,4);
TASK_PP(16'h15801,4);
TASK_PP(16'h15802,4);
TASK_PP(16'h15803,4);
TASK_PP(16'h15804,4);
TASK_PP(16'h15805,4);
TASK_PP(16'h15806,4);
TASK_PP(16'h15807,4);
TASK_PP(16'h15808,4);
TASK_PP(16'h15809,4);
TASK_PP(16'h1580A,4);
TASK_PP(16'h1580B,4);
TASK_PP(16'h1580C,4);
TASK_PP(16'h1580D,4);
TASK_PP(16'h1580E,4);
TASK_PP(16'h1580F,4);
TASK_PP(16'h15810,4);
TASK_PP(16'h15811,4);
TASK_PP(16'h15812,4);
TASK_PP(16'h15813,4);
TASK_PP(16'h15814,4);
TASK_PP(16'h15815,4);
TASK_PP(16'h15816,4);
TASK_PP(16'h15817,4);
TASK_PP(16'h15818,4);
TASK_PP(16'h15819,4);
TASK_PP(16'h1581A,4);
TASK_PP(16'h1581B,4);
TASK_PP(16'h1581C,4);
TASK_PP(16'h1581D,4);
TASK_PP(16'h1581E,4);
TASK_PP(16'h1581F,4);
TASK_PP(16'h15820,4);
TASK_PP(16'h15821,4);
TASK_PP(16'h15822,4);
TASK_PP(16'h15823,4);
TASK_PP(16'h15824,4);
TASK_PP(16'h15825,4);
TASK_PP(16'h15826,4);
TASK_PP(16'h15827,4);
TASK_PP(16'h15828,4);
TASK_PP(16'h15829,4);
TASK_PP(16'h1582A,4);
TASK_PP(16'h1582B,4);
TASK_PP(16'h1582C,4);
TASK_PP(16'h1582D,4);
TASK_PP(16'h1582E,4);
TASK_PP(16'h1582F,4);
TASK_PP(16'h15830,4);
TASK_PP(16'h15831,4);
TASK_PP(16'h15832,4);
TASK_PP(16'h15833,4);
TASK_PP(16'h15834,4);
TASK_PP(16'h15835,4);
TASK_PP(16'h15836,4);
TASK_PP(16'h15837,4);
TASK_PP(16'h15838,4);
TASK_PP(16'h15839,4);
TASK_PP(16'h1583A,4);
TASK_PP(16'h1583B,4);
TASK_PP(16'h1583C,4);
TASK_PP(16'h1583D,4);
TASK_PP(16'h1583E,4);
TASK_PP(16'h1583F,4);
TASK_PP(16'h15840,4);
TASK_PP(16'h15841,4);
TASK_PP(16'h15842,4);
TASK_PP(16'h15843,4);
TASK_PP(16'h15844,4);
TASK_PP(16'h15845,4);
TASK_PP(16'h15846,4);
TASK_PP(16'h15847,4);
TASK_PP(16'h15848,4);
TASK_PP(16'h15849,4);
TASK_PP(16'h1584A,4);
TASK_PP(16'h1584B,4);
TASK_PP(16'h1584C,4);
TASK_PP(16'h1584D,4);
TASK_PP(16'h1584E,4);
TASK_PP(16'h1584F,4);
TASK_PP(16'h15850,4);
TASK_PP(16'h15851,4);
TASK_PP(16'h15852,4);
TASK_PP(16'h15853,4);
TASK_PP(16'h15854,4);
TASK_PP(16'h15855,4);
TASK_PP(16'h15856,4);
TASK_PP(16'h15857,4);
TASK_PP(16'h15858,4);
TASK_PP(16'h15859,4);
TASK_PP(16'h1585A,4);
TASK_PP(16'h1585B,4);
TASK_PP(16'h1585C,4);
TASK_PP(16'h1585D,4);
TASK_PP(16'h1585E,4);
TASK_PP(16'h1585F,4);
TASK_PP(16'h15860,4);
TASK_PP(16'h15861,4);
TASK_PP(16'h15862,4);
TASK_PP(16'h15863,4);
TASK_PP(16'h15864,4);
TASK_PP(16'h15865,4);
TASK_PP(16'h15866,4);
TASK_PP(16'h15867,4);
TASK_PP(16'h15868,4);
TASK_PP(16'h15869,4);
TASK_PP(16'h1586A,4);
TASK_PP(16'h1586B,4);
TASK_PP(16'h1586C,4);
TASK_PP(16'h1586D,4);
TASK_PP(16'h1586E,4);
TASK_PP(16'h1586F,4);
TASK_PP(16'h15870,4);
TASK_PP(16'h15871,4);
TASK_PP(16'h15872,4);
TASK_PP(16'h15873,4);
TASK_PP(16'h15874,4);
TASK_PP(16'h15875,4);
TASK_PP(16'h15876,4);
TASK_PP(16'h15877,4);
TASK_PP(16'h15878,4);
TASK_PP(16'h15879,4);
TASK_PP(16'h1587A,4);
TASK_PP(16'h1587B,4);
TASK_PP(16'h1587C,4);
TASK_PP(16'h1587D,4);
TASK_PP(16'h1587E,4);
TASK_PP(16'h1587F,4);
TASK_PP(16'h15880,4);
TASK_PP(16'h15881,4);
TASK_PP(16'h15882,4);
TASK_PP(16'h15883,4);
TASK_PP(16'h15884,4);
TASK_PP(16'h15885,4);
TASK_PP(16'h15886,4);
TASK_PP(16'h15887,4);
TASK_PP(16'h15888,4);
TASK_PP(16'h15889,4);
TASK_PP(16'h1588A,4);
TASK_PP(16'h1588B,4);
TASK_PP(16'h1588C,4);
TASK_PP(16'h1588D,4);
TASK_PP(16'h1588E,4);
TASK_PP(16'h1588F,4);
TASK_PP(16'h15890,4);
TASK_PP(16'h15891,4);
TASK_PP(16'h15892,4);
TASK_PP(16'h15893,4);
TASK_PP(16'h15894,4);
TASK_PP(16'h15895,4);
TASK_PP(16'h15896,4);
TASK_PP(16'h15897,4);
TASK_PP(16'h15898,4);
TASK_PP(16'h15899,4);
TASK_PP(16'h1589A,4);
TASK_PP(16'h1589B,4);
TASK_PP(16'h1589C,4);
TASK_PP(16'h1589D,4);
TASK_PP(16'h1589E,4);
TASK_PP(16'h1589F,4);
TASK_PP(16'h158A0,4);
TASK_PP(16'h158A1,4);
TASK_PP(16'h158A2,4);
TASK_PP(16'h158A3,4);
TASK_PP(16'h158A4,4);
TASK_PP(16'h158A5,4);
TASK_PP(16'h158A6,4);
TASK_PP(16'h158A7,4);
TASK_PP(16'h158A8,4);
TASK_PP(16'h158A9,4);
TASK_PP(16'h158AA,4);
TASK_PP(16'h158AB,4);
TASK_PP(16'h158AC,4);
TASK_PP(16'h158AD,4);
TASK_PP(16'h158AE,4);
TASK_PP(16'h158AF,4);
TASK_PP(16'h158B0,4);
TASK_PP(16'h158B1,4);
TASK_PP(16'h158B2,4);
TASK_PP(16'h158B3,4);
TASK_PP(16'h158B4,4);
TASK_PP(16'h158B5,4);
TASK_PP(16'h158B6,4);
TASK_PP(16'h158B7,4);
TASK_PP(16'h158B8,4);
TASK_PP(16'h158B9,4);
TASK_PP(16'h158BA,4);
TASK_PP(16'h158BB,4);
TASK_PP(16'h158BC,4);
TASK_PP(16'h158BD,4);
TASK_PP(16'h158BE,4);
TASK_PP(16'h158BF,4);
TASK_PP(16'h158C0,4);
TASK_PP(16'h158C1,4);
TASK_PP(16'h158C2,4);
TASK_PP(16'h158C3,4);
TASK_PP(16'h158C4,4);
TASK_PP(16'h158C5,4);
TASK_PP(16'h158C6,4);
TASK_PP(16'h158C7,4);
TASK_PP(16'h158C8,4);
TASK_PP(16'h158C9,4);
TASK_PP(16'h158CA,4);
TASK_PP(16'h158CB,4);
TASK_PP(16'h158CC,4);
TASK_PP(16'h158CD,4);
TASK_PP(16'h158CE,4);
TASK_PP(16'h158CF,4);
TASK_PP(16'h158D0,4);
TASK_PP(16'h158D1,4);
TASK_PP(16'h158D2,4);
TASK_PP(16'h158D3,4);
TASK_PP(16'h158D4,4);
TASK_PP(16'h158D5,4);
TASK_PP(16'h158D6,4);
TASK_PP(16'h158D7,4);
TASK_PP(16'h158D8,4);
TASK_PP(16'h158D9,4);
TASK_PP(16'h158DA,4);
TASK_PP(16'h158DB,4);
TASK_PP(16'h158DC,4);
TASK_PP(16'h158DD,4);
TASK_PP(16'h158DE,4);
TASK_PP(16'h158DF,4);
TASK_PP(16'h158E0,4);
TASK_PP(16'h158E1,4);
TASK_PP(16'h158E2,4);
TASK_PP(16'h158E3,4);
TASK_PP(16'h158E4,4);
TASK_PP(16'h158E5,4);
TASK_PP(16'h158E6,4);
TASK_PP(16'h158E7,4);
TASK_PP(16'h158E8,4);
TASK_PP(16'h158E9,4);
TASK_PP(16'h158EA,4);
TASK_PP(16'h158EB,4);
TASK_PP(16'h158EC,4);
TASK_PP(16'h158ED,4);
TASK_PP(16'h158EE,4);
TASK_PP(16'h158EF,4);
TASK_PP(16'h158F0,4);
TASK_PP(16'h158F1,4);
TASK_PP(16'h158F2,4);
TASK_PP(16'h158F3,4);
TASK_PP(16'h158F4,4);
TASK_PP(16'h158F5,4);
TASK_PP(16'h158F6,4);
TASK_PP(16'h158F7,4);
TASK_PP(16'h158F8,4);
TASK_PP(16'h158F9,4);
TASK_PP(16'h158FA,4);
TASK_PP(16'h158FB,4);
TASK_PP(16'h158FC,4);
TASK_PP(16'h158FD,4);
TASK_PP(16'h158FE,4);
TASK_PP(16'h158FF,4);
TASK_PP(16'h15900,4);
TASK_PP(16'h15901,4);
TASK_PP(16'h15902,4);
TASK_PP(16'h15903,4);
TASK_PP(16'h15904,4);
TASK_PP(16'h15905,4);
TASK_PP(16'h15906,4);
TASK_PP(16'h15907,4);
TASK_PP(16'h15908,4);
TASK_PP(16'h15909,4);
TASK_PP(16'h1590A,4);
TASK_PP(16'h1590B,4);
TASK_PP(16'h1590C,4);
TASK_PP(16'h1590D,4);
TASK_PP(16'h1590E,4);
TASK_PP(16'h1590F,4);
TASK_PP(16'h15910,4);
TASK_PP(16'h15911,4);
TASK_PP(16'h15912,4);
TASK_PP(16'h15913,4);
TASK_PP(16'h15914,4);
TASK_PP(16'h15915,4);
TASK_PP(16'h15916,4);
TASK_PP(16'h15917,4);
TASK_PP(16'h15918,4);
TASK_PP(16'h15919,4);
TASK_PP(16'h1591A,4);
TASK_PP(16'h1591B,4);
TASK_PP(16'h1591C,4);
TASK_PP(16'h1591D,4);
TASK_PP(16'h1591E,4);
TASK_PP(16'h1591F,4);
TASK_PP(16'h15920,4);
TASK_PP(16'h15921,4);
TASK_PP(16'h15922,4);
TASK_PP(16'h15923,4);
TASK_PP(16'h15924,4);
TASK_PP(16'h15925,4);
TASK_PP(16'h15926,4);
TASK_PP(16'h15927,4);
TASK_PP(16'h15928,4);
TASK_PP(16'h15929,4);
TASK_PP(16'h1592A,4);
TASK_PP(16'h1592B,4);
TASK_PP(16'h1592C,4);
TASK_PP(16'h1592D,4);
TASK_PP(16'h1592E,4);
TASK_PP(16'h1592F,4);
TASK_PP(16'h15930,4);
TASK_PP(16'h15931,4);
TASK_PP(16'h15932,4);
TASK_PP(16'h15933,4);
TASK_PP(16'h15934,4);
TASK_PP(16'h15935,4);
TASK_PP(16'h15936,4);
TASK_PP(16'h15937,4);
TASK_PP(16'h15938,4);
TASK_PP(16'h15939,4);
TASK_PP(16'h1593A,4);
TASK_PP(16'h1593B,4);
TASK_PP(16'h1593C,4);
TASK_PP(16'h1593D,4);
TASK_PP(16'h1593E,4);
TASK_PP(16'h1593F,4);
TASK_PP(16'h15940,4);
TASK_PP(16'h15941,4);
TASK_PP(16'h15942,4);
TASK_PP(16'h15943,4);
TASK_PP(16'h15944,4);
TASK_PP(16'h15945,4);
TASK_PP(16'h15946,4);
TASK_PP(16'h15947,4);
TASK_PP(16'h15948,4);
TASK_PP(16'h15949,4);
TASK_PP(16'h1594A,4);
TASK_PP(16'h1594B,4);
TASK_PP(16'h1594C,4);
TASK_PP(16'h1594D,4);
TASK_PP(16'h1594E,4);
TASK_PP(16'h1594F,4);
TASK_PP(16'h15950,4);
TASK_PP(16'h15951,4);
TASK_PP(16'h15952,4);
TASK_PP(16'h15953,4);
TASK_PP(16'h15954,4);
TASK_PP(16'h15955,4);
TASK_PP(16'h15956,4);
TASK_PP(16'h15957,4);
TASK_PP(16'h15958,4);
TASK_PP(16'h15959,4);
TASK_PP(16'h1595A,4);
TASK_PP(16'h1595B,4);
TASK_PP(16'h1595C,4);
TASK_PP(16'h1595D,4);
TASK_PP(16'h1595E,4);
TASK_PP(16'h1595F,4);
TASK_PP(16'h15960,4);
TASK_PP(16'h15961,4);
TASK_PP(16'h15962,4);
TASK_PP(16'h15963,4);
TASK_PP(16'h15964,4);
TASK_PP(16'h15965,4);
TASK_PP(16'h15966,4);
TASK_PP(16'h15967,4);
TASK_PP(16'h15968,4);
TASK_PP(16'h15969,4);
TASK_PP(16'h1596A,4);
TASK_PP(16'h1596B,4);
TASK_PP(16'h1596C,4);
TASK_PP(16'h1596D,4);
TASK_PP(16'h1596E,4);
TASK_PP(16'h1596F,4);
TASK_PP(16'h15970,4);
TASK_PP(16'h15971,4);
TASK_PP(16'h15972,4);
TASK_PP(16'h15973,4);
TASK_PP(16'h15974,4);
TASK_PP(16'h15975,4);
TASK_PP(16'h15976,4);
TASK_PP(16'h15977,4);
TASK_PP(16'h15978,4);
TASK_PP(16'h15979,4);
TASK_PP(16'h1597A,4);
TASK_PP(16'h1597B,4);
TASK_PP(16'h1597C,4);
TASK_PP(16'h1597D,4);
TASK_PP(16'h1597E,4);
TASK_PP(16'h1597F,4);
TASK_PP(16'h15980,4);
TASK_PP(16'h15981,4);
TASK_PP(16'h15982,4);
TASK_PP(16'h15983,4);
TASK_PP(16'h15984,4);
TASK_PP(16'h15985,4);
TASK_PP(16'h15986,4);
TASK_PP(16'h15987,4);
TASK_PP(16'h15988,4);
TASK_PP(16'h15989,4);
TASK_PP(16'h1598A,4);
TASK_PP(16'h1598B,4);
TASK_PP(16'h1598C,4);
TASK_PP(16'h1598D,4);
TASK_PP(16'h1598E,4);
TASK_PP(16'h1598F,4);
TASK_PP(16'h15990,4);
TASK_PP(16'h15991,4);
TASK_PP(16'h15992,4);
TASK_PP(16'h15993,4);
TASK_PP(16'h15994,4);
TASK_PP(16'h15995,4);
TASK_PP(16'h15996,4);
TASK_PP(16'h15997,4);
TASK_PP(16'h15998,4);
TASK_PP(16'h15999,4);
TASK_PP(16'h1599A,4);
TASK_PP(16'h1599B,4);
TASK_PP(16'h1599C,4);
TASK_PP(16'h1599D,4);
TASK_PP(16'h1599E,4);
TASK_PP(16'h1599F,4);
TASK_PP(16'h159A0,4);
TASK_PP(16'h159A1,4);
TASK_PP(16'h159A2,4);
TASK_PP(16'h159A3,4);
TASK_PP(16'h159A4,4);
TASK_PP(16'h159A5,4);
TASK_PP(16'h159A6,4);
TASK_PP(16'h159A7,4);
TASK_PP(16'h159A8,4);
TASK_PP(16'h159A9,4);
TASK_PP(16'h159AA,4);
TASK_PP(16'h159AB,4);
TASK_PP(16'h159AC,4);
TASK_PP(16'h159AD,4);
TASK_PP(16'h159AE,4);
TASK_PP(16'h159AF,4);
TASK_PP(16'h159B0,4);
TASK_PP(16'h159B1,4);
TASK_PP(16'h159B2,4);
TASK_PP(16'h159B3,4);
TASK_PP(16'h159B4,4);
TASK_PP(16'h159B5,4);
TASK_PP(16'h159B6,4);
TASK_PP(16'h159B7,4);
TASK_PP(16'h159B8,4);
TASK_PP(16'h159B9,4);
TASK_PP(16'h159BA,4);
TASK_PP(16'h159BB,4);
TASK_PP(16'h159BC,4);
TASK_PP(16'h159BD,4);
TASK_PP(16'h159BE,4);
TASK_PP(16'h159BF,4);
TASK_PP(16'h159C0,4);
TASK_PP(16'h159C1,4);
TASK_PP(16'h159C2,4);
TASK_PP(16'h159C3,4);
TASK_PP(16'h159C4,4);
TASK_PP(16'h159C5,4);
TASK_PP(16'h159C6,4);
TASK_PP(16'h159C7,4);
TASK_PP(16'h159C8,4);
TASK_PP(16'h159C9,4);
TASK_PP(16'h159CA,4);
TASK_PP(16'h159CB,4);
TASK_PP(16'h159CC,4);
TASK_PP(16'h159CD,4);
TASK_PP(16'h159CE,4);
TASK_PP(16'h159CF,4);
TASK_PP(16'h159D0,4);
TASK_PP(16'h159D1,4);
TASK_PP(16'h159D2,4);
TASK_PP(16'h159D3,4);
TASK_PP(16'h159D4,4);
TASK_PP(16'h159D5,4);
TASK_PP(16'h159D6,4);
TASK_PP(16'h159D7,4);
TASK_PP(16'h159D8,4);
TASK_PP(16'h159D9,4);
TASK_PP(16'h159DA,4);
TASK_PP(16'h159DB,4);
TASK_PP(16'h159DC,4);
TASK_PP(16'h159DD,4);
TASK_PP(16'h159DE,4);
TASK_PP(16'h159DF,4);
TASK_PP(16'h159E0,4);
TASK_PP(16'h159E1,4);
TASK_PP(16'h159E2,4);
TASK_PP(16'h159E3,4);
TASK_PP(16'h159E4,4);
TASK_PP(16'h159E5,4);
TASK_PP(16'h159E6,4);
TASK_PP(16'h159E7,4);
TASK_PP(16'h159E8,4);
TASK_PP(16'h159E9,4);
TASK_PP(16'h159EA,4);
TASK_PP(16'h159EB,4);
TASK_PP(16'h159EC,4);
TASK_PP(16'h159ED,4);
TASK_PP(16'h159EE,4);
TASK_PP(16'h159EF,4);
TASK_PP(16'h159F0,4);
TASK_PP(16'h159F1,4);
TASK_PP(16'h159F2,4);
TASK_PP(16'h159F3,4);
TASK_PP(16'h159F4,4);
TASK_PP(16'h159F5,4);
TASK_PP(16'h159F6,4);
TASK_PP(16'h159F7,4);
TASK_PP(16'h159F8,4);
TASK_PP(16'h159F9,4);
TASK_PP(16'h159FA,4);
TASK_PP(16'h159FB,4);
TASK_PP(16'h159FC,4);
TASK_PP(16'h159FD,4);
TASK_PP(16'h159FE,4);
TASK_PP(16'h159FF,4);
TASK_PP(16'h15A00,4);
TASK_PP(16'h15A01,4);
TASK_PP(16'h15A02,4);
TASK_PP(16'h15A03,4);
TASK_PP(16'h15A04,4);
TASK_PP(16'h15A05,4);
TASK_PP(16'h15A06,4);
TASK_PP(16'h15A07,4);
TASK_PP(16'h15A08,4);
TASK_PP(16'h15A09,4);
TASK_PP(16'h15A0A,4);
TASK_PP(16'h15A0B,4);
TASK_PP(16'h15A0C,4);
TASK_PP(16'h15A0D,4);
TASK_PP(16'h15A0E,4);
TASK_PP(16'h15A0F,4);
TASK_PP(16'h15A10,4);
TASK_PP(16'h15A11,4);
TASK_PP(16'h15A12,4);
TASK_PP(16'h15A13,4);
TASK_PP(16'h15A14,4);
TASK_PP(16'h15A15,4);
TASK_PP(16'h15A16,4);
TASK_PP(16'h15A17,4);
TASK_PP(16'h15A18,4);
TASK_PP(16'h15A19,4);
TASK_PP(16'h15A1A,4);
TASK_PP(16'h15A1B,4);
TASK_PP(16'h15A1C,4);
TASK_PP(16'h15A1D,4);
TASK_PP(16'h15A1E,4);
TASK_PP(16'h15A1F,4);
TASK_PP(16'h15A20,4);
TASK_PP(16'h15A21,4);
TASK_PP(16'h15A22,4);
TASK_PP(16'h15A23,4);
TASK_PP(16'h15A24,4);
TASK_PP(16'h15A25,4);
TASK_PP(16'h15A26,4);
TASK_PP(16'h15A27,4);
TASK_PP(16'h15A28,4);
TASK_PP(16'h15A29,4);
TASK_PP(16'h15A2A,4);
TASK_PP(16'h15A2B,4);
TASK_PP(16'h15A2C,4);
TASK_PP(16'h15A2D,4);
TASK_PP(16'h15A2E,4);
TASK_PP(16'h15A2F,4);
TASK_PP(16'h15A30,4);
TASK_PP(16'h15A31,4);
TASK_PP(16'h15A32,4);
TASK_PP(16'h15A33,4);
TASK_PP(16'h15A34,4);
TASK_PP(16'h15A35,4);
TASK_PP(16'h15A36,4);
TASK_PP(16'h15A37,4);
TASK_PP(16'h15A38,4);
TASK_PP(16'h15A39,4);
TASK_PP(16'h15A3A,4);
TASK_PP(16'h15A3B,4);
TASK_PP(16'h15A3C,4);
TASK_PP(16'h15A3D,4);
TASK_PP(16'h15A3E,4);
TASK_PP(16'h15A3F,4);
TASK_PP(16'h15A40,4);
TASK_PP(16'h15A41,4);
TASK_PP(16'h15A42,4);
TASK_PP(16'h15A43,4);
TASK_PP(16'h15A44,4);
TASK_PP(16'h15A45,4);
TASK_PP(16'h15A46,4);
TASK_PP(16'h15A47,4);
TASK_PP(16'h15A48,4);
TASK_PP(16'h15A49,4);
TASK_PP(16'h15A4A,4);
TASK_PP(16'h15A4B,4);
TASK_PP(16'h15A4C,4);
TASK_PP(16'h15A4D,4);
TASK_PP(16'h15A4E,4);
TASK_PP(16'h15A4F,4);
TASK_PP(16'h15A50,4);
TASK_PP(16'h15A51,4);
TASK_PP(16'h15A52,4);
TASK_PP(16'h15A53,4);
TASK_PP(16'h15A54,4);
TASK_PP(16'h15A55,4);
TASK_PP(16'h15A56,4);
TASK_PP(16'h15A57,4);
TASK_PP(16'h15A58,4);
TASK_PP(16'h15A59,4);
TASK_PP(16'h15A5A,4);
TASK_PP(16'h15A5B,4);
TASK_PP(16'h15A5C,4);
TASK_PP(16'h15A5D,4);
TASK_PP(16'h15A5E,4);
TASK_PP(16'h15A5F,4);
TASK_PP(16'h15A60,4);
TASK_PP(16'h15A61,4);
TASK_PP(16'h15A62,4);
TASK_PP(16'h15A63,4);
TASK_PP(16'h15A64,4);
TASK_PP(16'h15A65,4);
TASK_PP(16'h15A66,4);
TASK_PP(16'h15A67,4);
TASK_PP(16'h15A68,4);
TASK_PP(16'h15A69,4);
TASK_PP(16'h15A6A,4);
TASK_PP(16'h15A6B,4);
TASK_PP(16'h15A6C,4);
TASK_PP(16'h15A6D,4);
TASK_PP(16'h15A6E,4);
TASK_PP(16'h15A6F,4);
TASK_PP(16'h15A70,4);
TASK_PP(16'h15A71,4);
TASK_PP(16'h15A72,4);
TASK_PP(16'h15A73,4);
TASK_PP(16'h15A74,4);
TASK_PP(16'h15A75,4);
TASK_PP(16'h15A76,4);
TASK_PP(16'h15A77,4);
TASK_PP(16'h15A78,4);
TASK_PP(16'h15A79,4);
TASK_PP(16'h15A7A,4);
TASK_PP(16'h15A7B,4);
TASK_PP(16'h15A7C,4);
TASK_PP(16'h15A7D,4);
TASK_PP(16'h15A7E,4);
TASK_PP(16'h15A7F,4);
TASK_PP(16'h15A80,4);
TASK_PP(16'h15A81,4);
TASK_PP(16'h15A82,4);
TASK_PP(16'h15A83,4);
TASK_PP(16'h15A84,4);
TASK_PP(16'h15A85,4);
TASK_PP(16'h15A86,4);
TASK_PP(16'h15A87,4);
TASK_PP(16'h15A88,4);
TASK_PP(16'h15A89,4);
TASK_PP(16'h15A8A,4);
TASK_PP(16'h15A8B,4);
TASK_PP(16'h15A8C,4);
TASK_PP(16'h15A8D,4);
TASK_PP(16'h15A8E,4);
TASK_PP(16'h15A8F,4);
TASK_PP(16'h15A90,4);
TASK_PP(16'h15A91,4);
TASK_PP(16'h15A92,4);
TASK_PP(16'h15A93,4);
TASK_PP(16'h15A94,4);
TASK_PP(16'h15A95,4);
TASK_PP(16'h15A96,4);
TASK_PP(16'h15A97,4);
TASK_PP(16'h15A98,4);
TASK_PP(16'h15A99,4);
TASK_PP(16'h15A9A,4);
TASK_PP(16'h15A9B,4);
TASK_PP(16'h15A9C,4);
TASK_PP(16'h15A9D,4);
TASK_PP(16'h15A9E,4);
TASK_PP(16'h15A9F,4);
TASK_PP(16'h15AA0,4);
TASK_PP(16'h15AA1,4);
TASK_PP(16'h15AA2,4);
TASK_PP(16'h15AA3,4);
TASK_PP(16'h15AA4,4);
TASK_PP(16'h15AA5,4);
TASK_PP(16'h15AA6,4);
TASK_PP(16'h15AA7,4);
TASK_PP(16'h15AA8,4);
TASK_PP(16'h15AA9,4);
TASK_PP(16'h15AAA,4);
TASK_PP(16'h15AAB,4);
TASK_PP(16'h15AAC,4);
TASK_PP(16'h15AAD,4);
TASK_PP(16'h15AAE,4);
TASK_PP(16'h15AAF,4);
TASK_PP(16'h15AB0,4);
TASK_PP(16'h15AB1,4);
TASK_PP(16'h15AB2,4);
TASK_PP(16'h15AB3,4);
TASK_PP(16'h15AB4,4);
TASK_PP(16'h15AB5,4);
TASK_PP(16'h15AB6,4);
TASK_PP(16'h15AB7,4);
TASK_PP(16'h15AB8,4);
TASK_PP(16'h15AB9,4);
TASK_PP(16'h15ABA,4);
TASK_PP(16'h15ABB,4);
TASK_PP(16'h15ABC,4);
TASK_PP(16'h15ABD,4);
TASK_PP(16'h15ABE,4);
TASK_PP(16'h15ABF,4);
TASK_PP(16'h15AC0,4);
TASK_PP(16'h15AC1,4);
TASK_PP(16'h15AC2,4);
TASK_PP(16'h15AC3,4);
TASK_PP(16'h15AC4,4);
TASK_PP(16'h15AC5,4);
TASK_PP(16'h15AC6,4);
TASK_PP(16'h15AC7,4);
TASK_PP(16'h15AC8,4);
TASK_PP(16'h15AC9,4);
TASK_PP(16'h15ACA,4);
TASK_PP(16'h15ACB,4);
TASK_PP(16'h15ACC,4);
TASK_PP(16'h15ACD,4);
TASK_PP(16'h15ACE,4);
TASK_PP(16'h15ACF,4);
TASK_PP(16'h15AD0,4);
TASK_PP(16'h15AD1,4);
TASK_PP(16'h15AD2,4);
TASK_PP(16'h15AD3,4);
TASK_PP(16'h15AD4,4);
TASK_PP(16'h15AD5,4);
TASK_PP(16'h15AD6,4);
TASK_PP(16'h15AD7,4);
TASK_PP(16'h15AD8,4);
TASK_PP(16'h15AD9,4);
TASK_PP(16'h15ADA,4);
TASK_PP(16'h15ADB,4);
TASK_PP(16'h15ADC,4);
TASK_PP(16'h15ADD,4);
TASK_PP(16'h15ADE,4);
TASK_PP(16'h15ADF,4);
TASK_PP(16'h15AE0,4);
TASK_PP(16'h15AE1,4);
TASK_PP(16'h15AE2,4);
TASK_PP(16'h15AE3,4);
TASK_PP(16'h15AE4,4);
TASK_PP(16'h15AE5,4);
TASK_PP(16'h15AE6,4);
TASK_PP(16'h15AE7,4);
TASK_PP(16'h15AE8,4);
TASK_PP(16'h15AE9,4);
TASK_PP(16'h15AEA,4);
TASK_PP(16'h15AEB,4);
TASK_PP(16'h15AEC,4);
TASK_PP(16'h15AED,4);
TASK_PP(16'h15AEE,4);
TASK_PP(16'h15AEF,4);
TASK_PP(16'h15AF0,4);
TASK_PP(16'h15AF1,4);
TASK_PP(16'h15AF2,4);
TASK_PP(16'h15AF3,4);
TASK_PP(16'h15AF4,4);
TASK_PP(16'h15AF5,4);
TASK_PP(16'h15AF6,4);
TASK_PP(16'h15AF7,4);
TASK_PP(16'h15AF8,4);
TASK_PP(16'h15AF9,4);
TASK_PP(16'h15AFA,4);
TASK_PP(16'h15AFB,4);
TASK_PP(16'h15AFC,4);
TASK_PP(16'h15AFD,4);
TASK_PP(16'h15AFE,4);
TASK_PP(16'h15AFF,4);
TASK_PP(16'h15B00,4);
TASK_PP(16'h15B01,4);
TASK_PP(16'h15B02,4);
TASK_PP(16'h15B03,4);
TASK_PP(16'h15B04,4);
TASK_PP(16'h15B05,4);
TASK_PP(16'h15B06,4);
TASK_PP(16'h15B07,4);
TASK_PP(16'h15B08,4);
TASK_PP(16'h15B09,4);
TASK_PP(16'h15B0A,4);
TASK_PP(16'h15B0B,4);
TASK_PP(16'h15B0C,4);
TASK_PP(16'h15B0D,4);
TASK_PP(16'h15B0E,4);
TASK_PP(16'h15B0F,4);
TASK_PP(16'h15B10,4);
TASK_PP(16'h15B11,4);
TASK_PP(16'h15B12,4);
TASK_PP(16'h15B13,4);
TASK_PP(16'h15B14,4);
TASK_PP(16'h15B15,4);
TASK_PP(16'h15B16,4);
TASK_PP(16'h15B17,4);
TASK_PP(16'h15B18,4);
TASK_PP(16'h15B19,4);
TASK_PP(16'h15B1A,4);
TASK_PP(16'h15B1B,4);
TASK_PP(16'h15B1C,4);
TASK_PP(16'h15B1D,4);
TASK_PP(16'h15B1E,4);
TASK_PP(16'h15B1F,4);
TASK_PP(16'h15B20,4);
TASK_PP(16'h15B21,4);
TASK_PP(16'h15B22,4);
TASK_PP(16'h15B23,4);
TASK_PP(16'h15B24,4);
TASK_PP(16'h15B25,4);
TASK_PP(16'h15B26,4);
TASK_PP(16'h15B27,4);
TASK_PP(16'h15B28,4);
TASK_PP(16'h15B29,4);
TASK_PP(16'h15B2A,4);
TASK_PP(16'h15B2B,4);
TASK_PP(16'h15B2C,4);
TASK_PP(16'h15B2D,4);
TASK_PP(16'h15B2E,4);
TASK_PP(16'h15B2F,4);
TASK_PP(16'h15B30,4);
TASK_PP(16'h15B31,4);
TASK_PP(16'h15B32,4);
TASK_PP(16'h15B33,4);
TASK_PP(16'h15B34,4);
TASK_PP(16'h15B35,4);
TASK_PP(16'h15B36,4);
TASK_PP(16'h15B37,4);
TASK_PP(16'h15B38,4);
TASK_PP(16'h15B39,4);
TASK_PP(16'h15B3A,4);
TASK_PP(16'h15B3B,4);
TASK_PP(16'h15B3C,4);
TASK_PP(16'h15B3D,4);
TASK_PP(16'h15B3E,4);
TASK_PP(16'h15B3F,4);
TASK_PP(16'h15B40,4);
TASK_PP(16'h15B41,4);
TASK_PP(16'h15B42,4);
TASK_PP(16'h15B43,4);
TASK_PP(16'h15B44,4);
TASK_PP(16'h15B45,4);
TASK_PP(16'h15B46,4);
TASK_PP(16'h15B47,4);
TASK_PP(16'h15B48,4);
TASK_PP(16'h15B49,4);
TASK_PP(16'h15B4A,4);
TASK_PP(16'h15B4B,4);
TASK_PP(16'h15B4C,4);
TASK_PP(16'h15B4D,4);
TASK_PP(16'h15B4E,4);
TASK_PP(16'h15B4F,4);
TASK_PP(16'h15B50,4);
TASK_PP(16'h15B51,4);
TASK_PP(16'h15B52,4);
TASK_PP(16'h15B53,4);
TASK_PP(16'h15B54,4);
TASK_PP(16'h15B55,4);
TASK_PP(16'h15B56,4);
TASK_PP(16'h15B57,4);
TASK_PP(16'h15B58,4);
TASK_PP(16'h15B59,4);
TASK_PP(16'h15B5A,4);
TASK_PP(16'h15B5B,4);
TASK_PP(16'h15B5C,4);
TASK_PP(16'h15B5D,4);
TASK_PP(16'h15B5E,4);
TASK_PP(16'h15B5F,4);
TASK_PP(16'h15B60,4);
TASK_PP(16'h15B61,4);
TASK_PP(16'h15B62,4);
TASK_PP(16'h15B63,4);
TASK_PP(16'h15B64,4);
TASK_PP(16'h15B65,4);
TASK_PP(16'h15B66,4);
TASK_PP(16'h15B67,4);
TASK_PP(16'h15B68,4);
TASK_PP(16'h15B69,4);
TASK_PP(16'h15B6A,4);
TASK_PP(16'h15B6B,4);
TASK_PP(16'h15B6C,4);
TASK_PP(16'h15B6D,4);
TASK_PP(16'h15B6E,4);
TASK_PP(16'h15B6F,4);
TASK_PP(16'h15B70,4);
TASK_PP(16'h15B71,4);
TASK_PP(16'h15B72,4);
TASK_PP(16'h15B73,4);
TASK_PP(16'h15B74,4);
TASK_PP(16'h15B75,4);
TASK_PP(16'h15B76,4);
TASK_PP(16'h15B77,4);
TASK_PP(16'h15B78,4);
TASK_PP(16'h15B79,4);
TASK_PP(16'h15B7A,4);
TASK_PP(16'h15B7B,4);
TASK_PP(16'h15B7C,4);
TASK_PP(16'h15B7D,4);
TASK_PP(16'h15B7E,4);
TASK_PP(16'h15B7F,4);
TASK_PP(16'h15B80,4);
TASK_PP(16'h15B81,4);
TASK_PP(16'h15B82,4);
TASK_PP(16'h15B83,4);
TASK_PP(16'h15B84,4);
TASK_PP(16'h15B85,4);
TASK_PP(16'h15B86,4);
TASK_PP(16'h15B87,4);
TASK_PP(16'h15B88,4);
TASK_PP(16'h15B89,4);
TASK_PP(16'h15B8A,4);
TASK_PP(16'h15B8B,4);
TASK_PP(16'h15B8C,4);
TASK_PP(16'h15B8D,4);
TASK_PP(16'h15B8E,4);
TASK_PP(16'h15B8F,4);
TASK_PP(16'h15B90,4);
TASK_PP(16'h15B91,4);
TASK_PP(16'h15B92,4);
TASK_PP(16'h15B93,4);
TASK_PP(16'h15B94,4);
TASK_PP(16'h15B95,4);
TASK_PP(16'h15B96,4);
TASK_PP(16'h15B97,4);
TASK_PP(16'h15B98,4);
TASK_PP(16'h15B99,4);
TASK_PP(16'h15B9A,4);
TASK_PP(16'h15B9B,4);
TASK_PP(16'h15B9C,4);
TASK_PP(16'h15B9D,4);
TASK_PP(16'h15B9E,4);
TASK_PP(16'h15B9F,4);
TASK_PP(16'h15BA0,4);
TASK_PP(16'h15BA1,4);
TASK_PP(16'h15BA2,4);
TASK_PP(16'h15BA3,4);
TASK_PP(16'h15BA4,4);
TASK_PP(16'h15BA5,4);
TASK_PP(16'h15BA6,4);
TASK_PP(16'h15BA7,4);
TASK_PP(16'h15BA8,4);
TASK_PP(16'h15BA9,4);
TASK_PP(16'h15BAA,4);
TASK_PP(16'h15BAB,4);
TASK_PP(16'h15BAC,4);
TASK_PP(16'h15BAD,4);
TASK_PP(16'h15BAE,4);
TASK_PP(16'h15BAF,4);
TASK_PP(16'h15BB0,4);
TASK_PP(16'h15BB1,4);
TASK_PP(16'h15BB2,4);
TASK_PP(16'h15BB3,4);
TASK_PP(16'h15BB4,4);
TASK_PP(16'h15BB5,4);
TASK_PP(16'h15BB6,4);
TASK_PP(16'h15BB7,4);
TASK_PP(16'h15BB8,4);
TASK_PP(16'h15BB9,4);
TASK_PP(16'h15BBA,4);
TASK_PP(16'h15BBB,4);
TASK_PP(16'h15BBC,4);
TASK_PP(16'h15BBD,4);
TASK_PP(16'h15BBE,4);
TASK_PP(16'h15BBF,4);
TASK_PP(16'h15BC0,4);
TASK_PP(16'h15BC1,4);
TASK_PP(16'h15BC2,4);
TASK_PP(16'h15BC3,4);
TASK_PP(16'h15BC4,4);
TASK_PP(16'h15BC5,4);
TASK_PP(16'h15BC6,4);
TASK_PP(16'h15BC7,4);
TASK_PP(16'h15BC8,4);
TASK_PP(16'h15BC9,4);
TASK_PP(16'h15BCA,4);
TASK_PP(16'h15BCB,4);
TASK_PP(16'h15BCC,4);
TASK_PP(16'h15BCD,4);
TASK_PP(16'h15BCE,4);
TASK_PP(16'h15BCF,4);
TASK_PP(16'h15BD0,4);
TASK_PP(16'h15BD1,4);
TASK_PP(16'h15BD2,4);
TASK_PP(16'h15BD3,4);
TASK_PP(16'h15BD4,4);
TASK_PP(16'h15BD5,4);
TASK_PP(16'h15BD6,4);
TASK_PP(16'h15BD7,4);
TASK_PP(16'h15BD8,4);
TASK_PP(16'h15BD9,4);
TASK_PP(16'h15BDA,4);
TASK_PP(16'h15BDB,4);
TASK_PP(16'h15BDC,4);
TASK_PP(16'h15BDD,4);
TASK_PP(16'h15BDE,4);
TASK_PP(16'h15BDF,4);
TASK_PP(16'h15BE0,4);
TASK_PP(16'h15BE1,4);
TASK_PP(16'h15BE2,4);
TASK_PP(16'h15BE3,4);
TASK_PP(16'h15BE4,4);
TASK_PP(16'h15BE5,4);
TASK_PP(16'h15BE6,4);
TASK_PP(16'h15BE7,4);
TASK_PP(16'h15BE8,4);
TASK_PP(16'h15BE9,4);
TASK_PP(16'h15BEA,4);
TASK_PP(16'h15BEB,4);
TASK_PP(16'h15BEC,4);
TASK_PP(16'h15BED,4);
TASK_PP(16'h15BEE,4);
TASK_PP(16'h15BEF,4);
TASK_PP(16'h15BF0,4);
TASK_PP(16'h15BF1,4);
TASK_PP(16'h15BF2,4);
TASK_PP(16'h15BF3,4);
TASK_PP(16'h15BF4,4);
TASK_PP(16'h15BF5,4);
TASK_PP(16'h15BF6,4);
TASK_PP(16'h15BF7,4);
TASK_PP(16'h15BF8,4);
TASK_PP(16'h15BF9,4);
TASK_PP(16'h15BFA,4);
TASK_PP(16'h15BFB,4);
TASK_PP(16'h15BFC,4);
TASK_PP(16'h15BFD,4);
TASK_PP(16'h15BFE,4);
TASK_PP(16'h15BFF,4);
TASK_PP(16'h15C00,4);
TASK_PP(16'h15C01,4);
TASK_PP(16'h15C02,4);
TASK_PP(16'h15C03,4);
TASK_PP(16'h15C04,4);
TASK_PP(16'h15C05,4);
TASK_PP(16'h15C06,4);
TASK_PP(16'h15C07,4);
TASK_PP(16'h15C08,4);
TASK_PP(16'h15C09,4);
TASK_PP(16'h15C0A,4);
TASK_PP(16'h15C0B,4);
TASK_PP(16'h15C0C,4);
TASK_PP(16'h15C0D,4);
TASK_PP(16'h15C0E,4);
TASK_PP(16'h15C0F,4);
TASK_PP(16'h15C10,4);
TASK_PP(16'h15C11,4);
TASK_PP(16'h15C12,4);
TASK_PP(16'h15C13,4);
TASK_PP(16'h15C14,4);
TASK_PP(16'h15C15,4);
TASK_PP(16'h15C16,4);
TASK_PP(16'h15C17,4);
TASK_PP(16'h15C18,4);
TASK_PP(16'h15C19,4);
TASK_PP(16'h15C1A,4);
TASK_PP(16'h15C1B,4);
TASK_PP(16'h15C1C,4);
TASK_PP(16'h15C1D,4);
TASK_PP(16'h15C1E,4);
TASK_PP(16'h15C1F,4);
TASK_PP(16'h15C20,4);
TASK_PP(16'h15C21,4);
TASK_PP(16'h15C22,4);
TASK_PP(16'h15C23,4);
TASK_PP(16'h15C24,4);
TASK_PP(16'h15C25,4);
TASK_PP(16'h15C26,4);
TASK_PP(16'h15C27,4);
TASK_PP(16'h15C28,4);
TASK_PP(16'h15C29,4);
TASK_PP(16'h15C2A,4);
TASK_PP(16'h15C2B,4);
TASK_PP(16'h15C2C,4);
TASK_PP(16'h15C2D,4);
TASK_PP(16'h15C2E,4);
TASK_PP(16'h15C2F,4);
TASK_PP(16'h15C30,4);
TASK_PP(16'h15C31,4);
TASK_PP(16'h15C32,4);
TASK_PP(16'h15C33,4);
TASK_PP(16'h15C34,4);
TASK_PP(16'h15C35,4);
TASK_PP(16'h15C36,4);
TASK_PP(16'h15C37,4);
TASK_PP(16'h15C38,4);
TASK_PP(16'h15C39,4);
TASK_PP(16'h15C3A,4);
TASK_PP(16'h15C3B,4);
TASK_PP(16'h15C3C,4);
TASK_PP(16'h15C3D,4);
TASK_PP(16'h15C3E,4);
TASK_PP(16'h15C3F,4);
TASK_PP(16'h15C40,4);
TASK_PP(16'h15C41,4);
TASK_PP(16'h15C42,4);
TASK_PP(16'h15C43,4);
TASK_PP(16'h15C44,4);
TASK_PP(16'h15C45,4);
TASK_PP(16'h15C46,4);
TASK_PP(16'h15C47,4);
TASK_PP(16'h15C48,4);
TASK_PP(16'h15C49,4);
TASK_PP(16'h15C4A,4);
TASK_PP(16'h15C4B,4);
TASK_PP(16'h15C4C,4);
TASK_PP(16'h15C4D,4);
TASK_PP(16'h15C4E,4);
TASK_PP(16'h15C4F,4);
TASK_PP(16'h15C50,4);
TASK_PP(16'h15C51,4);
TASK_PP(16'h15C52,4);
TASK_PP(16'h15C53,4);
TASK_PP(16'h15C54,4);
TASK_PP(16'h15C55,4);
TASK_PP(16'h15C56,4);
TASK_PP(16'h15C57,4);
TASK_PP(16'h15C58,4);
TASK_PP(16'h15C59,4);
TASK_PP(16'h15C5A,4);
TASK_PP(16'h15C5B,4);
TASK_PP(16'h15C5C,4);
TASK_PP(16'h15C5D,4);
TASK_PP(16'h15C5E,4);
TASK_PP(16'h15C5F,4);
TASK_PP(16'h15C60,4);
TASK_PP(16'h15C61,4);
TASK_PP(16'h15C62,4);
TASK_PP(16'h15C63,4);
TASK_PP(16'h15C64,4);
TASK_PP(16'h15C65,4);
TASK_PP(16'h15C66,4);
TASK_PP(16'h15C67,4);
TASK_PP(16'h15C68,4);
TASK_PP(16'h15C69,4);
TASK_PP(16'h15C6A,4);
TASK_PP(16'h15C6B,4);
TASK_PP(16'h15C6C,4);
TASK_PP(16'h15C6D,4);
TASK_PP(16'h15C6E,4);
TASK_PP(16'h15C6F,4);
TASK_PP(16'h15C70,4);
TASK_PP(16'h15C71,4);
TASK_PP(16'h15C72,4);
TASK_PP(16'h15C73,4);
TASK_PP(16'h15C74,4);
TASK_PP(16'h15C75,4);
TASK_PP(16'h15C76,4);
TASK_PP(16'h15C77,4);
TASK_PP(16'h15C78,4);
TASK_PP(16'h15C79,4);
TASK_PP(16'h15C7A,4);
TASK_PP(16'h15C7B,4);
TASK_PP(16'h15C7C,4);
TASK_PP(16'h15C7D,4);
TASK_PP(16'h15C7E,4);
TASK_PP(16'h15C7F,4);
TASK_PP(16'h15C80,4);
TASK_PP(16'h15C81,4);
TASK_PP(16'h15C82,4);
TASK_PP(16'h15C83,4);
TASK_PP(16'h15C84,4);
TASK_PP(16'h15C85,4);
TASK_PP(16'h15C86,4);
TASK_PP(16'h15C87,4);
TASK_PP(16'h15C88,4);
TASK_PP(16'h15C89,4);
TASK_PP(16'h15C8A,4);
TASK_PP(16'h15C8B,4);
TASK_PP(16'h15C8C,4);
TASK_PP(16'h15C8D,4);
TASK_PP(16'h15C8E,4);
TASK_PP(16'h15C8F,4);
TASK_PP(16'h15C90,4);
TASK_PP(16'h15C91,4);
TASK_PP(16'h15C92,4);
TASK_PP(16'h15C93,4);
TASK_PP(16'h15C94,4);
TASK_PP(16'h15C95,4);
TASK_PP(16'h15C96,4);
TASK_PP(16'h15C97,4);
TASK_PP(16'h15C98,4);
TASK_PP(16'h15C99,4);
TASK_PP(16'h15C9A,4);
TASK_PP(16'h15C9B,4);
TASK_PP(16'h15C9C,4);
TASK_PP(16'h15C9D,4);
TASK_PP(16'h15C9E,4);
TASK_PP(16'h15C9F,4);
TASK_PP(16'h15CA0,4);
TASK_PP(16'h15CA1,4);
TASK_PP(16'h15CA2,4);
TASK_PP(16'h15CA3,4);
TASK_PP(16'h15CA4,4);
TASK_PP(16'h15CA5,4);
TASK_PP(16'h15CA6,4);
TASK_PP(16'h15CA7,4);
TASK_PP(16'h15CA8,4);
TASK_PP(16'h15CA9,4);
TASK_PP(16'h15CAA,4);
TASK_PP(16'h15CAB,4);
TASK_PP(16'h15CAC,4);
TASK_PP(16'h15CAD,4);
TASK_PP(16'h15CAE,4);
TASK_PP(16'h15CAF,4);
TASK_PP(16'h15CB0,4);
TASK_PP(16'h15CB1,4);
TASK_PP(16'h15CB2,4);
TASK_PP(16'h15CB3,4);
TASK_PP(16'h15CB4,4);
TASK_PP(16'h15CB5,4);
TASK_PP(16'h15CB6,4);
TASK_PP(16'h15CB7,4);
TASK_PP(16'h15CB8,4);
TASK_PP(16'h15CB9,4);
TASK_PP(16'h15CBA,4);
TASK_PP(16'h15CBB,4);
TASK_PP(16'h15CBC,4);
TASK_PP(16'h15CBD,4);
TASK_PP(16'h15CBE,4);
TASK_PP(16'h15CBF,4);
TASK_PP(16'h15CC0,4);
TASK_PP(16'h15CC1,4);
TASK_PP(16'h15CC2,4);
TASK_PP(16'h15CC3,4);
TASK_PP(16'h15CC4,4);
TASK_PP(16'h15CC5,4);
TASK_PP(16'h15CC6,4);
TASK_PP(16'h15CC7,4);
TASK_PP(16'h15CC8,4);
TASK_PP(16'h15CC9,4);
TASK_PP(16'h15CCA,4);
TASK_PP(16'h15CCB,4);
TASK_PP(16'h15CCC,4);
TASK_PP(16'h15CCD,4);
TASK_PP(16'h15CCE,4);
TASK_PP(16'h15CCF,4);
TASK_PP(16'h15CD0,4);
TASK_PP(16'h15CD1,4);
TASK_PP(16'h15CD2,4);
TASK_PP(16'h15CD3,4);
TASK_PP(16'h15CD4,4);
TASK_PP(16'h15CD5,4);
TASK_PP(16'h15CD6,4);
TASK_PP(16'h15CD7,4);
TASK_PP(16'h15CD8,4);
TASK_PP(16'h15CD9,4);
TASK_PP(16'h15CDA,4);
TASK_PP(16'h15CDB,4);
TASK_PP(16'h15CDC,4);
TASK_PP(16'h15CDD,4);
TASK_PP(16'h15CDE,4);
TASK_PP(16'h15CDF,4);
TASK_PP(16'h15CE0,4);
TASK_PP(16'h15CE1,4);
TASK_PP(16'h15CE2,4);
TASK_PP(16'h15CE3,4);
TASK_PP(16'h15CE4,4);
TASK_PP(16'h15CE5,4);
TASK_PP(16'h15CE6,4);
TASK_PP(16'h15CE7,4);
TASK_PP(16'h15CE8,4);
TASK_PP(16'h15CE9,4);
TASK_PP(16'h15CEA,4);
TASK_PP(16'h15CEB,4);
TASK_PP(16'h15CEC,4);
TASK_PP(16'h15CED,4);
TASK_PP(16'h15CEE,4);
TASK_PP(16'h15CEF,4);
TASK_PP(16'h15CF0,4);
TASK_PP(16'h15CF1,4);
TASK_PP(16'h15CF2,4);
TASK_PP(16'h15CF3,4);
TASK_PP(16'h15CF4,4);
TASK_PP(16'h15CF5,4);
TASK_PP(16'h15CF6,4);
TASK_PP(16'h15CF7,4);
TASK_PP(16'h15CF8,4);
TASK_PP(16'h15CF9,4);
TASK_PP(16'h15CFA,4);
TASK_PP(16'h15CFB,4);
TASK_PP(16'h15CFC,4);
TASK_PP(16'h15CFD,4);
TASK_PP(16'h15CFE,4);
TASK_PP(16'h15CFF,4);
TASK_PP(16'h15D00,4);
TASK_PP(16'h15D01,4);
TASK_PP(16'h15D02,4);
TASK_PP(16'h15D03,4);
TASK_PP(16'h15D04,4);
TASK_PP(16'h15D05,4);
TASK_PP(16'h15D06,4);
TASK_PP(16'h15D07,4);
TASK_PP(16'h15D08,4);
TASK_PP(16'h15D09,4);
TASK_PP(16'h15D0A,4);
TASK_PP(16'h15D0B,4);
TASK_PP(16'h15D0C,4);
TASK_PP(16'h15D0D,4);
TASK_PP(16'h15D0E,4);
TASK_PP(16'h15D0F,4);
TASK_PP(16'h15D10,4);
TASK_PP(16'h15D11,4);
TASK_PP(16'h15D12,4);
TASK_PP(16'h15D13,4);
TASK_PP(16'h15D14,4);
TASK_PP(16'h15D15,4);
TASK_PP(16'h15D16,4);
TASK_PP(16'h15D17,4);
TASK_PP(16'h15D18,4);
TASK_PP(16'h15D19,4);
TASK_PP(16'h15D1A,4);
TASK_PP(16'h15D1B,4);
TASK_PP(16'h15D1C,4);
TASK_PP(16'h15D1D,4);
TASK_PP(16'h15D1E,4);
TASK_PP(16'h15D1F,4);
TASK_PP(16'h15D20,4);
TASK_PP(16'h15D21,4);
TASK_PP(16'h15D22,4);
TASK_PP(16'h15D23,4);
TASK_PP(16'h15D24,4);
TASK_PP(16'h15D25,4);
TASK_PP(16'h15D26,4);
TASK_PP(16'h15D27,4);
TASK_PP(16'h15D28,4);
TASK_PP(16'h15D29,4);
TASK_PP(16'h15D2A,4);
TASK_PP(16'h15D2B,4);
TASK_PP(16'h15D2C,4);
TASK_PP(16'h15D2D,4);
TASK_PP(16'h15D2E,4);
TASK_PP(16'h15D2F,4);
TASK_PP(16'h15D30,4);
TASK_PP(16'h15D31,4);
TASK_PP(16'h15D32,4);
TASK_PP(16'h15D33,4);
TASK_PP(16'h15D34,4);
TASK_PP(16'h15D35,4);
TASK_PP(16'h15D36,4);
TASK_PP(16'h15D37,4);
TASK_PP(16'h15D38,4);
TASK_PP(16'h15D39,4);
TASK_PP(16'h15D3A,4);
TASK_PP(16'h15D3B,4);
TASK_PP(16'h15D3C,4);
TASK_PP(16'h15D3D,4);
TASK_PP(16'h15D3E,4);
TASK_PP(16'h15D3F,4);
TASK_PP(16'h15D40,4);
TASK_PP(16'h15D41,4);
TASK_PP(16'h15D42,4);
TASK_PP(16'h15D43,4);
TASK_PP(16'h15D44,4);
TASK_PP(16'h15D45,4);
TASK_PP(16'h15D46,4);
TASK_PP(16'h15D47,4);
TASK_PP(16'h15D48,4);
TASK_PP(16'h15D49,4);
TASK_PP(16'h15D4A,4);
TASK_PP(16'h15D4B,4);
TASK_PP(16'h15D4C,4);
TASK_PP(16'h15D4D,4);
TASK_PP(16'h15D4E,4);
TASK_PP(16'h15D4F,4);
TASK_PP(16'h15D50,4);
TASK_PP(16'h15D51,4);
TASK_PP(16'h15D52,4);
TASK_PP(16'h15D53,4);
TASK_PP(16'h15D54,4);
TASK_PP(16'h15D55,4);
TASK_PP(16'h15D56,4);
TASK_PP(16'h15D57,4);
TASK_PP(16'h15D58,4);
TASK_PP(16'h15D59,4);
TASK_PP(16'h15D5A,4);
TASK_PP(16'h15D5B,4);
TASK_PP(16'h15D5C,4);
TASK_PP(16'h15D5D,4);
TASK_PP(16'h15D5E,4);
TASK_PP(16'h15D5F,4);
TASK_PP(16'h15D60,4);
TASK_PP(16'h15D61,4);
TASK_PP(16'h15D62,4);
TASK_PP(16'h15D63,4);
TASK_PP(16'h15D64,4);
TASK_PP(16'h15D65,4);
TASK_PP(16'h15D66,4);
TASK_PP(16'h15D67,4);
TASK_PP(16'h15D68,4);
TASK_PP(16'h15D69,4);
TASK_PP(16'h15D6A,4);
TASK_PP(16'h15D6B,4);
TASK_PP(16'h15D6C,4);
TASK_PP(16'h15D6D,4);
TASK_PP(16'h15D6E,4);
TASK_PP(16'h15D6F,4);
TASK_PP(16'h15D70,4);
TASK_PP(16'h15D71,4);
TASK_PP(16'h15D72,4);
TASK_PP(16'h15D73,4);
TASK_PP(16'h15D74,4);
TASK_PP(16'h15D75,4);
TASK_PP(16'h15D76,4);
TASK_PP(16'h15D77,4);
TASK_PP(16'h15D78,4);
TASK_PP(16'h15D79,4);
TASK_PP(16'h15D7A,4);
TASK_PP(16'h15D7B,4);
TASK_PP(16'h15D7C,4);
TASK_PP(16'h15D7D,4);
TASK_PP(16'h15D7E,4);
TASK_PP(16'h15D7F,4);
TASK_PP(16'h15D80,4);
TASK_PP(16'h15D81,4);
TASK_PP(16'h15D82,4);
TASK_PP(16'h15D83,4);
TASK_PP(16'h15D84,4);
TASK_PP(16'h15D85,4);
TASK_PP(16'h15D86,4);
TASK_PP(16'h15D87,4);
TASK_PP(16'h15D88,4);
TASK_PP(16'h15D89,4);
TASK_PP(16'h15D8A,4);
TASK_PP(16'h15D8B,4);
TASK_PP(16'h15D8C,4);
TASK_PP(16'h15D8D,4);
TASK_PP(16'h15D8E,4);
TASK_PP(16'h15D8F,4);
TASK_PP(16'h15D90,4);
TASK_PP(16'h15D91,4);
TASK_PP(16'h15D92,4);
TASK_PP(16'h15D93,4);
TASK_PP(16'h15D94,4);
TASK_PP(16'h15D95,4);
TASK_PP(16'h15D96,4);
TASK_PP(16'h15D97,4);
TASK_PP(16'h15D98,4);
TASK_PP(16'h15D99,4);
TASK_PP(16'h15D9A,4);
TASK_PP(16'h15D9B,4);
TASK_PP(16'h15D9C,4);
TASK_PP(16'h15D9D,4);
TASK_PP(16'h15D9E,4);
TASK_PP(16'h15D9F,4);
TASK_PP(16'h15DA0,4);
TASK_PP(16'h15DA1,4);
TASK_PP(16'h15DA2,4);
TASK_PP(16'h15DA3,4);
TASK_PP(16'h15DA4,4);
TASK_PP(16'h15DA5,4);
TASK_PP(16'h15DA6,4);
TASK_PP(16'h15DA7,4);
TASK_PP(16'h15DA8,4);
TASK_PP(16'h15DA9,4);
TASK_PP(16'h15DAA,4);
TASK_PP(16'h15DAB,4);
TASK_PP(16'h15DAC,4);
TASK_PP(16'h15DAD,4);
TASK_PP(16'h15DAE,4);
TASK_PP(16'h15DAF,4);
TASK_PP(16'h15DB0,4);
TASK_PP(16'h15DB1,4);
TASK_PP(16'h15DB2,4);
TASK_PP(16'h15DB3,4);
TASK_PP(16'h15DB4,4);
TASK_PP(16'h15DB5,4);
TASK_PP(16'h15DB6,4);
TASK_PP(16'h15DB7,4);
TASK_PP(16'h15DB8,4);
TASK_PP(16'h15DB9,4);
TASK_PP(16'h15DBA,4);
TASK_PP(16'h15DBB,4);
TASK_PP(16'h15DBC,4);
TASK_PP(16'h15DBD,4);
TASK_PP(16'h15DBE,4);
TASK_PP(16'h15DBF,4);
TASK_PP(16'h15DC0,4);
TASK_PP(16'h15DC1,4);
TASK_PP(16'h15DC2,4);
TASK_PP(16'h15DC3,4);
TASK_PP(16'h15DC4,4);
TASK_PP(16'h15DC5,4);
TASK_PP(16'h15DC6,4);
TASK_PP(16'h15DC7,4);
TASK_PP(16'h15DC8,4);
TASK_PP(16'h15DC9,4);
TASK_PP(16'h15DCA,4);
TASK_PP(16'h15DCB,4);
TASK_PP(16'h15DCC,4);
TASK_PP(16'h15DCD,4);
TASK_PP(16'h15DCE,4);
TASK_PP(16'h15DCF,4);
TASK_PP(16'h15DD0,4);
TASK_PP(16'h15DD1,4);
TASK_PP(16'h15DD2,4);
TASK_PP(16'h15DD3,4);
TASK_PP(16'h15DD4,4);
TASK_PP(16'h15DD5,4);
TASK_PP(16'h15DD6,4);
TASK_PP(16'h15DD7,4);
TASK_PP(16'h15DD8,4);
TASK_PP(16'h15DD9,4);
TASK_PP(16'h15DDA,4);
TASK_PP(16'h15DDB,4);
TASK_PP(16'h15DDC,4);
TASK_PP(16'h15DDD,4);
TASK_PP(16'h15DDE,4);
TASK_PP(16'h15DDF,4);
TASK_PP(16'h15DE0,4);
TASK_PP(16'h15DE1,4);
TASK_PP(16'h15DE2,4);
TASK_PP(16'h15DE3,4);
TASK_PP(16'h15DE4,4);
TASK_PP(16'h15DE5,4);
TASK_PP(16'h15DE6,4);
TASK_PP(16'h15DE7,4);
TASK_PP(16'h15DE8,4);
TASK_PP(16'h15DE9,4);
TASK_PP(16'h15DEA,4);
TASK_PP(16'h15DEB,4);
TASK_PP(16'h15DEC,4);
TASK_PP(16'h15DED,4);
TASK_PP(16'h15DEE,4);
TASK_PP(16'h15DEF,4);
TASK_PP(16'h15DF0,4);
TASK_PP(16'h15DF1,4);
TASK_PP(16'h15DF2,4);
TASK_PP(16'h15DF3,4);
TASK_PP(16'h15DF4,4);
TASK_PP(16'h15DF5,4);
TASK_PP(16'h15DF6,4);
TASK_PP(16'h15DF7,4);
TASK_PP(16'h15DF8,4);
TASK_PP(16'h15DF9,4);
TASK_PP(16'h15DFA,4);
TASK_PP(16'h15DFB,4);
TASK_PP(16'h15DFC,4);
TASK_PP(16'h15DFD,4);
TASK_PP(16'h15DFE,4);
TASK_PP(16'h15DFF,4);
TASK_PP(16'h15E00,4);
TASK_PP(16'h15E01,4);
TASK_PP(16'h15E02,4);
TASK_PP(16'h15E03,4);
TASK_PP(16'h15E04,4);
TASK_PP(16'h15E05,4);
TASK_PP(16'h15E06,4);
TASK_PP(16'h15E07,4);
TASK_PP(16'h15E08,4);
TASK_PP(16'h15E09,4);
TASK_PP(16'h15E0A,4);
TASK_PP(16'h15E0B,4);
TASK_PP(16'h15E0C,4);
TASK_PP(16'h15E0D,4);
TASK_PP(16'h15E0E,4);
TASK_PP(16'h15E0F,4);
TASK_PP(16'h15E10,4);
TASK_PP(16'h15E11,4);
TASK_PP(16'h15E12,4);
TASK_PP(16'h15E13,4);
TASK_PP(16'h15E14,4);
TASK_PP(16'h15E15,4);
TASK_PP(16'h15E16,4);
TASK_PP(16'h15E17,4);
TASK_PP(16'h15E18,4);
TASK_PP(16'h15E19,4);
TASK_PP(16'h15E1A,4);
TASK_PP(16'h15E1B,4);
TASK_PP(16'h15E1C,4);
TASK_PP(16'h15E1D,4);
TASK_PP(16'h15E1E,4);
TASK_PP(16'h15E1F,4);
TASK_PP(16'h15E20,4);
TASK_PP(16'h15E21,4);
TASK_PP(16'h15E22,4);
TASK_PP(16'h15E23,4);
TASK_PP(16'h15E24,4);
TASK_PP(16'h15E25,4);
TASK_PP(16'h15E26,4);
TASK_PP(16'h15E27,4);
TASK_PP(16'h15E28,4);
TASK_PP(16'h15E29,4);
TASK_PP(16'h15E2A,4);
TASK_PP(16'h15E2B,4);
TASK_PP(16'h15E2C,4);
TASK_PP(16'h15E2D,4);
TASK_PP(16'h15E2E,4);
TASK_PP(16'h15E2F,4);
TASK_PP(16'h15E30,4);
TASK_PP(16'h15E31,4);
TASK_PP(16'h15E32,4);
TASK_PP(16'h15E33,4);
TASK_PP(16'h15E34,4);
TASK_PP(16'h15E35,4);
TASK_PP(16'h15E36,4);
TASK_PP(16'h15E37,4);
TASK_PP(16'h15E38,4);
TASK_PP(16'h15E39,4);
TASK_PP(16'h15E3A,4);
TASK_PP(16'h15E3B,4);
TASK_PP(16'h15E3C,4);
TASK_PP(16'h15E3D,4);
TASK_PP(16'h15E3E,4);
TASK_PP(16'h15E3F,4);
TASK_PP(16'h15E40,4);
TASK_PP(16'h15E41,4);
TASK_PP(16'h15E42,4);
TASK_PP(16'h15E43,4);
TASK_PP(16'h15E44,4);
TASK_PP(16'h15E45,4);
TASK_PP(16'h15E46,4);
TASK_PP(16'h15E47,4);
TASK_PP(16'h15E48,4);
TASK_PP(16'h15E49,4);
TASK_PP(16'h15E4A,4);
TASK_PP(16'h15E4B,4);
TASK_PP(16'h15E4C,4);
TASK_PP(16'h15E4D,4);
TASK_PP(16'h15E4E,4);
TASK_PP(16'h15E4F,4);
TASK_PP(16'h15E50,4);
TASK_PP(16'h15E51,4);
TASK_PP(16'h15E52,4);
TASK_PP(16'h15E53,4);
TASK_PP(16'h15E54,4);
TASK_PP(16'h15E55,4);
TASK_PP(16'h15E56,4);
TASK_PP(16'h15E57,4);
TASK_PP(16'h15E58,4);
TASK_PP(16'h15E59,4);
TASK_PP(16'h15E5A,4);
TASK_PP(16'h15E5B,4);
TASK_PP(16'h15E5C,4);
TASK_PP(16'h15E5D,4);
TASK_PP(16'h15E5E,4);
TASK_PP(16'h15E5F,4);
TASK_PP(16'h15E60,4);
TASK_PP(16'h15E61,4);
TASK_PP(16'h15E62,4);
TASK_PP(16'h15E63,4);
TASK_PP(16'h15E64,4);
TASK_PP(16'h15E65,4);
TASK_PP(16'h15E66,4);
TASK_PP(16'h15E67,4);
TASK_PP(16'h15E68,4);
TASK_PP(16'h15E69,4);
TASK_PP(16'h15E6A,4);
TASK_PP(16'h15E6B,4);
TASK_PP(16'h15E6C,4);
TASK_PP(16'h15E6D,4);
TASK_PP(16'h15E6E,4);
TASK_PP(16'h15E6F,4);
TASK_PP(16'h15E70,4);
TASK_PP(16'h15E71,4);
TASK_PP(16'h15E72,4);
TASK_PP(16'h15E73,4);
TASK_PP(16'h15E74,4);
TASK_PP(16'h15E75,4);
TASK_PP(16'h15E76,4);
TASK_PP(16'h15E77,4);
TASK_PP(16'h15E78,4);
TASK_PP(16'h15E79,4);
TASK_PP(16'h15E7A,4);
TASK_PP(16'h15E7B,4);
TASK_PP(16'h15E7C,4);
TASK_PP(16'h15E7D,4);
TASK_PP(16'h15E7E,4);
TASK_PP(16'h15E7F,4);
TASK_PP(16'h15E80,4);
TASK_PP(16'h15E81,4);
TASK_PP(16'h15E82,4);
TASK_PP(16'h15E83,4);
TASK_PP(16'h15E84,4);
TASK_PP(16'h15E85,4);
TASK_PP(16'h15E86,4);
TASK_PP(16'h15E87,4);
TASK_PP(16'h15E88,4);
TASK_PP(16'h15E89,4);
TASK_PP(16'h15E8A,4);
TASK_PP(16'h15E8B,4);
TASK_PP(16'h15E8C,4);
TASK_PP(16'h15E8D,4);
TASK_PP(16'h15E8E,4);
TASK_PP(16'h15E8F,4);
TASK_PP(16'h15E90,4);
TASK_PP(16'h15E91,4);
TASK_PP(16'h15E92,4);
TASK_PP(16'h15E93,4);
TASK_PP(16'h15E94,4);
TASK_PP(16'h15E95,4);
TASK_PP(16'h15E96,4);
TASK_PP(16'h15E97,4);
TASK_PP(16'h15E98,4);
TASK_PP(16'h15E99,4);
TASK_PP(16'h15E9A,4);
TASK_PP(16'h15E9B,4);
TASK_PP(16'h15E9C,4);
TASK_PP(16'h15E9D,4);
TASK_PP(16'h15E9E,4);
TASK_PP(16'h15E9F,4);
TASK_PP(16'h15EA0,4);
TASK_PP(16'h15EA1,4);
TASK_PP(16'h15EA2,4);
TASK_PP(16'h15EA3,4);
TASK_PP(16'h15EA4,4);
TASK_PP(16'h15EA5,4);
TASK_PP(16'h15EA6,4);
TASK_PP(16'h15EA7,4);
TASK_PP(16'h15EA8,4);
TASK_PP(16'h15EA9,4);
TASK_PP(16'h15EAA,4);
TASK_PP(16'h15EAB,4);
TASK_PP(16'h15EAC,4);
TASK_PP(16'h15EAD,4);
TASK_PP(16'h15EAE,4);
TASK_PP(16'h15EAF,4);
TASK_PP(16'h15EB0,4);
TASK_PP(16'h15EB1,4);
TASK_PP(16'h15EB2,4);
TASK_PP(16'h15EB3,4);
TASK_PP(16'h15EB4,4);
TASK_PP(16'h15EB5,4);
TASK_PP(16'h15EB6,4);
TASK_PP(16'h15EB7,4);
TASK_PP(16'h15EB8,4);
TASK_PP(16'h15EB9,4);
TASK_PP(16'h15EBA,4);
TASK_PP(16'h15EBB,4);
TASK_PP(16'h15EBC,4);
TASK_PP(16'h15EBD,4);
TASK_PP(16'h15EBE,4);
TASK_PP(16'h15EBF,4);
TASK_PP(16'h15EC0,4);
TASK_PP(16'h15EC1,4);
TASK_PP(16'h15EC2,4);
TASK_PP(16'h15EC3,4);
TASK_PP(16'h15EC4,4);
TASK_PP(16'h15EC5,4);
TASK_PP(16'h15EC6,4);
TASK_PP(16'h15EC7,4);
TASK_PP(16'h15EC8,4);
TASK_PP(16'h15EC9,4);
TASK_PP(16'h15ECA,4);
TASK_PP(16'h15ECB,4);
TASK_PP(16'h15ECC,4);
TASK_PP(16'h15ECD,4);
TASK_PP(16'h15ECE,4);
TASK_PP(16'h15ECF,4);
TASK_PP(16'h15ED0,4);
TASK_PP(16'h15ED1,4);
TASK_PP(16'h15ED2,4);
TASK_PP(16'h15ED3,4);
TASK_PP(16'h15ED4,4);
TASK_PP(16'h15ED5,4);
TASK_PP(16'h15ED6,4);
TASK_PP(16'h15ED7,4);
TASK_PP(16'h15ED8,4);
TASK_PP(16'h15ED9,4);
TASK_PP(16'h15EDA,4);
TASK_PP(16'h15EDB,4);
TASK_PP(16'h15EDC,4);
TASK_PP(16'h15EDD,4);
TASK_PP(16'h15EDE,4);
TASK_PP(16'h15EDF,4);
TASK_PP(16'h15EE0,4);
TASK_PP(16'h15EE1,4);
TASK_PP(16'h15EE2,4);
TASK_PP(16'h15EE3,4);
TASK_PP(16'h15EE4,4);
TASK_PP(16'h15EE5,4);
TASK_PP(16'h15EE6,4);
TASK_PP(16'h15EE7,4);
TASK_PP(16'h15EE8,4);
TASK_PP(16'h15EE9,4);
TASK_PP(16'h15EEA,4);
TASK_PP(16'h15EEB,4);
TASK_PP(16'h15EEC,4);
TASK_PP(16'h15EED,4);
TASK_PP(16'h15EEE,4);
TASK_PP(16'h15EEF,4);
TASK_PP(16'h15EF0,4);
TASK_PP(16'h15EF1,4);
TASK_PP(16'h15EF2,4);
TASK_PP(16'h15EF3,4);
TASK_PP(16'h15EF4,4);
TASK_PP(16'h15EF5,4);
TASK_PP(16'h15EF6,4);
TASK_PP(16'h15EF7,4);
TASK_PP(16'h15EF8,4);
TASK_PP(16'h15EF9,4);
TASK_PP(16'h15EFA,4);
TASK_PP(16'h15EFB,4);
TASK_PP(16'h15EFC,4);
TASK_PP(16'h15EFD,4);
TASK_PP(16'h15EFE,4);
TASK_PP(16'h15EFF,4);
TASK_PP(16'h15F00,4);
TASK_PP(16'h15F01,4);
TASK_PP(16'h15F02,4);
TASK_PP(16'h15F03,4);
TASK_PP(16'h15F04,4);
TASK_PP(16'h15F05,4);
TASK_PP(16'h15F06,4);
TASK_PP(16'h15F07,4);
TASK_PP(16'h15F08,4);
TASK_PP(16'h15F09,4);
TASK_PP(16'h15F0A,4);
TASK_PP(16'h15F0B,4);
TASK_PP(16'h15F0C,4);
TASK_PP(16'h15F0D,4);
TASK_PP(16'h15F0E,4);
TASK_PP(16'h15F0F,4);
TASK_PP(16'h15F10,4);
TASK_PP(16'h15F11,4);
TASK_PP(16'h15F12,4);
TASK_PP(16'h15F13,4);
TASK_PP(16'h15F14,4);
TASK_PP(16'h15F15,4);
TASK_PP(16'h15F16,4);
TASK_PP(16'h15F17,4);
TASK_PP(16'h15F18,4);
TASK_PP(16'h15F19,4);
TASK_PP(16'h15F1A,4);
TASK_PP(16'h15F1B,4);
TASK_PP(16'h15F1C,4);
TASK_PP(16'h15F1D,4);
TASK_PP(16'h15F1E,4);
TASK_PP(16'h15F1F,4);
TASK_PP(16'h15F20,4);
TASK_PP(16'h15F21,4);
TASK_PP(16'h15F22,4);
TASK_PP(16'h15F23,4);
TASK_PP(16'h15F24,4);
TASK_PP(16'h15F25,4);
TASK_PP(16'h15F26,4);
TASK_PP(16'h15F27,4);
TASK_PP(16'h15F28,4);
TASK_PP(16'h15F29,4);
TASK_PP(16'h15F2A,4);
TASK_PP(16'h15F2B,4);
TASK_PP(16'h15F2C,4);
TASK_PP(16'h15F2D,4);
TASK_PP(16'h15F2E,4);
TASK_PP(16'h15F2F,4);
TASK_PP(16'h15F30,4);
TASK_PP(16'h15F31,4);
TASK_PP(16'h15F32,4);
TASK_PP(16'h15F33,4);
TASK_PP(16'h15F34,4);
TASK_PP(16'h15F35,4);
TASK_PP(16'h15F36,4);
TASK_PP(16'h15F37,4);
TASK_PP(16'h15F38,4);
TASK_PP(16'h15F39,4);
TASK_PP(16'h15F3A,4);
TASK_PP(16'h15F3B,4);
TASK_PP(16'h15F3C,4);
TASK_PP(16'h15F3D,4);
TASK_PP(16'h15F3E,4);
TASK_PP(16'h15F3F,4);
TASK_PP(16'h15F40,4);
TASK_PP(16'h15F41,4);
TASK_PP(16'h15F42,4);
TASK_PP(16'h15F43,4);
TASK_PP(16'h15F44,4);
TASK_PP(16'h15F45,4);
TASK_PP(16'h15F46,4);
TASK_PP(16'h15F47,4);
TASK_PP(16'h15F48,4);
TASK_PP(16'h15F49,4);
TASK_PP(16'h15F4A,4);
TASK_PP(16'h15F4B,4);
TASK_PP(16'h15F4C,4);
TASK_PP(16'h15F4D,4);
TASK_PP(16'h15F4E,4);
TASK_PP(16'h15F4F,4);
TASK_PP(16'h15F50,4);
TASK_PP(16'h15F51,4);
TASK_PP(16'h15F52,4);
TASK_PP(16'h15F53,4);
TASK_PP(16'h15F54,4);
TASK_PP(16'h15F55,4);
TASK_PP(16'h15F56,4);
TASK_PP(16'h15F57,4);
TASK_PP(16'h15F58,4);
TASK_PP(16'h15F59,4);
TASK_PP(16'h15F5A,4);
TASK_PP(16'h15F5B,4);
TASK_PP(16'h15F5C,4);
TASK_PP(16'h15F5D,4);
TASK_PP(16'h15F5E,4);
TASK_PP(16'h15F5F,4);
TASK_PP(16'h15F60,4);
TASK_PP(16'h15F61,4);
TASK_PP(16'h15F62,4);
TASK_PP(16'h15F63,4);
TASK_PP(16'h15F64,4);
TASK_PP(16'h15F65,4);
TASK_PP(16'h15F66,4);
TASK_PP(16'h15F67,4);
TASK_PP(16'h15F68,4);
TASK_PP(16'h15F69,4);
TASK_PP(16'h15F6A,4);
TASK_PP(16'h15F6B,4);
TASK_PP(16'h15F6C,4);
TASK_PP(16'h15F6D,4);
TASK_PP(16'h15F6E,4);
TASK_PP(16'h15F6F,4);
TASK_PP(16'h15F70,4);
TASK_PP(16'h15F71,4);
TASK_PP(16'h15F72,4);
TASK_PP(16'h15F73,4);
TASK_PP(16'h15F74,4);
TASK_PP(16'h15F75,4);
TASK_PP(16'h15F76,4);
TASK_PP(16'h15F77,4);
TASK_PP(16'h15F78,4);
TASK_PP(16'h15F79,4);
TASK_PP(16'h15F7A,4);
TASK_PP(16'h15F7B,4);
TASK_PP(16'h15F7C,4);
TASK_PP(16'h15F7D,4);
TASK_PP(16'h15F7E,4);
TASK_PP(16'h15F7F,4);
TASK_PP(16'h15F80,4);
TASK_PP(16'h15F81,4);
TASK_PP(16'h15F82,4);
TASK_PP(16'h15F83,4);
TASK_PP(16'h15F84,4);
TASK_PP(16'h15F85,4);
TASK_PP(16'h15F86,4);
TASK_PP(16'h15F87,4);
TASK_PP(16'h15F88,4);
TASK_PP(16'h15F89,4);
TASK_PP(16'h15F8A,4);
TASK_PP(16'h15F8B,4);
TASK_PP(16'h15F8C,4);
TASK_PP(16'h15F8D,4);
TASK_PP(16'h15F8E,4);
TASK_PP(16'h15F8F,4);
TASK_PP(16'h15F90,4);
TASK_PP(16'h15F91,4);
TASK_PP(16'h15F92,4);
TASK_PP(16'h15F93,4);
TASK_PP(16'h15F94,4);
TASK_PP(16'h15F95,4);
TASK_PP(16'h15F96,4);
TASK_PP(16'h15F97,4);
TASK_PP(16'h15F98,4);
TASK_PP(16'h15F99,4);
TASK_PP(16'h15F9A,4);
TASK_PP(16'h15F9B,4);
TASK_PP(16'h15F9C,4);
TASK_PP(16'h15F9D,4);
TASK_PP(16'h15F9E,4);
TASK_PP(16'h15F9F,4);
TASK_PP(16'h15FA0,4);
TASK_PP(16'h15FA1,4);
TASK_PP(16'h15FA2,4);
TASK_PP(16'h15FA3,4);
TASK_PP(16'h15FA4,4);
TASK_PP(16'h15FA5,4);
TASK_PP(16'h15FA6,4);
TASK_PP(16'h15FA7,4);
TASK_PP(16'h15FA8,4);
TASK_PP(16'h15FA9,4);
TASK_PP(16'h15FAA,4);
TASK_PP(16'h15FAB,4);
TASK_PP(16'h15FAC,4);
TASK_PP(16'h15FAD,4);
TASK_PP(16'h15FAE,4);
TASK_PP(16'h15FAF,4);
TASK_PP(16'h15FB0,4);
TASK_PP(16'h15FB1,4);
TASK_PP(16'h15FB2,4);
TASK_PP(16'h15FB3,4);
TASK_PP(16'h15FB4,4);
TASK_PP(16'h15FB5,4);
TASK_PP(16'h15FB6,4);
TASK_PP(16'h15FB7,4);
TASK_PP(16'h15FB8,4);
TASK_PP(16'h15FB9,4);
TASK_PP(16'h15FBA,4);
TASK_PP(16'h15FBB,4);
TASK_PP(16'h15FBC,4);
TASK_PP(16'h15FBD,4);
TASK_PP(16'h15FBE,4);
TASK_PP(16'h15FBF,4);
TASK_PP(16'h15FC0,4);
TASK_PP(16'h15FC1,4);
TASK_PP(16'h15FC2,4);
TASK_PP(16'h15FC3,4);
TASK_PP(16'h15FC4,4);
TASK_PP(16'h15FC5,4);
TASK_PP(16'h15FC6,4);
TASK_PP(16'h15FC7,4);
TASK_PP(16'h15FC8,4);
TASK_PP(16'h15FC9,4);
TASK_PP(16'h15FCA,4);
TASK_PP(16'h15FCB,4);
TASK_PP(16'h15FCC,4);
TASK_PP(16'h15FCD,4);
TASK_PP(16'h15FCE,4);
TASK_PP(16'h15FCF,4);
TASK_PP(16'h15FD0,4);
TASK_PP(16'h15FD1,4);
TASK_PP(16'h15FD2,4);
TASK_PP(16'h15FD3,4);
TASK_PP(16'h15FD4,4);
TASK_PP(16'h15FD5,4);
TASK_PP(16'h15FD6,4);
TASK_PP(16'h15FD7,4);
TASK_PP(16'h15FD8,4);
TASK_PP(16'h15FD9,4);
TASK_PP(16'h15FDA,4);
TASK_PP(16'h15FDB,4);
TASK_PP(16'h15FDC,4);
TASK_PP(16'h15FDD,4);
TASK_PP(16'h15FDE,4);
TASK_PP(16'h15FDF,4);
TASK_PP(16'h15FE0,4);
TASK_PP(16'h15FE1,4);
TASK_PP(16'h15FE2,4);
TASK_PP(16'h15FE3,4);
TASK_PP(16'h15FE4,4);
TASK_PP(16'h15FE5,4);
TASK_PP(16'h15FE6,4);
TASK_PP(16'h15FE7,4);
TASK_PP(16'h15FE8,4);
TASK_PP(16'h15FE9,4);
TASK_PP(16'h15FEA,4);
TASK_PP(16'h15FEB,4);
TASK_PP(16'h15FEC,4);
TASK_PP(16'h15FED,4);
TASK_PP(16'h15FEE,4);
TASK_PP(16'h15FEF,4);
TASK_PP(16'h15FF0,4);
TASK_PP(16'h15FF1,4);
TASK_PP(16'h15FF2,4);
TASK_PP(16'h15FF3,4);
TASK_PP(16'h15FF4,4);
TASK_PP(16'h15FF5,4);
TASK_PP(16'h15FF6,4);
TASK_PP(16'h15FF7,4);
TASK_PP(16'h15FF8,4);
TASK_PP(16'h15FF9,4);
TASK_PP(16'h15FFA,4);
TASK_PP(16'h15FFB,4);
TASK_PP(16'h15FFC,4);
TASK_PP(16'h15FFD,4);
TASK_PP(16'h15FFE,4);
TASK_PP(16'h15FFF,4);
TASK_PP(16'h16000,4);
TASK_PP(16'h16001,4);
TASK_PP(16'h16002,4);
TASK_PP(16'h16003,4);
TASK_PP(16'h16004,4);
TASK_PP(16'h16005,4);
TASK_PP(16'h16006,4);
TASK_PP(16'h16007,4);
TASK_PP(16'h16008,4);
TASK_PP(16'h16009,4);
TASK_PP(16'h1600A,4);
TASK_PP(16'h1600B,4);
TASK_PP(16'h1600C,4);
TASK_PP(16'h1600D,4);
TASK_PP(16'h1600E,4);
TASK_PP(16'h1600F,4);
TASK_PP(16'h16010,4);
TASK_PP(16'h16011,4);
TASK_PP(16'h16012,4);
TASK_PP(16'h16013,4);
TASK_PP(16'h16014,4);
TASK_PP(16'h16015,4);
TASK_PP(16'h16016,4);
TASK_PP(16'h16017,4);
TASK_PP(16'h16018,4);
TASK_PP(16'h16019,4);
TASK_PP(16'h1601A,4);
TASK_PP(16'h1601B,4);
TASK_PP(16'h1601C,4);
TASK_PP(16'h1601D,4);
TASK_PP(16'h1601E,4);
TASK_PP(16'h1601F,4);
TASK_PP(16'h16020,4);
TASK_PP(16'h16021,4);
TASK_PP(16'h16022,4);
TASK_PP(16'h16023,4);
TASK_PP(16'h16024,4);
TASK_PP(16'h16025,4);
TASK_PP(16'h16026,4);
TASK_PP(16'h16027,4);
TASK_PP(16'h16028,4);
TASK_PP(16'h16029,4);
TASK_PP(16'h1602A,4);
TASK_PP(16'h1602B,4);
TASK_PP(16'h1602C,4);
TASK_PP(16'h1602D,4);
TASK_PP(16'h1602E,4);
TASK_PP(16'h1602F,4);
TASK_PP(16'h16030,4);
TASK_PP(16'h16031,4);
TASK_PP(16'h16032,4);
TASK_PP(16'h16033,4);
TASK_PP(16'h16034,4);
TASK_PP(16'h16035,4);
TASK_PP(16'h16036,4);
TASK_PP(16'h16037,4);
TASK_PP(16'h16038,4);
TASK_PP(16'h16039,4);
TASK_PP(16'h1603A,4);
TASK_PP(16'h1603B,4);
TASK_PP(16'h1603C,4);
TASK_PP(16'h1603D,4);
TASK_PP(16'h1603E,4);
TASK_PP(16'h1603F,4);
TASK_PP(16'h16040,4);
TASK_PP(16'h16041,4);
TASK_PP(16'h16042,4);
TASK_PP(16'h16043,4);
TASK_PP(16'h16044,4);
TASK_PP(16'h16045,4);
TASK_PP(16'h16046,4);
TASK_PP(16'h16047,4);
TASK_PP(16'h16048,4);
TASK_PP(16'h16049,4);
TASK_PP(16'h1604A,4);
TASK_PP(16'h1604B,4);
TASK_PP(16'h1604C,4);
TASK_PP(16'h1604D,4);
TASK_PP(16'h1604E,4);
TASK_PP(16'h1604F,4);
TASK_PP(16'h16050,4);
TASK_PP(16'h16051,4);
TASK_PP(16'h16052,4);
TASK_PP(16'h16053,4);
TASK_PP(16'h16054,4);
TASK_PP(16'h16055,4);
TASK_PP(16'h16056,4);
TASK_PP(16'h16057,4);
TASK_PP(16'h16058,4);
TASK_PP(16'h16059,4);
TASK_PP(16'h1605A,4);
TASK_PP(16'h1605B,4);
TASK_PP(16'h1605C,4);
TASK_PP(16'h1605D,4);
TASK_PP(16'h1605E,4);
TASK_PP(16'h1605F,4);
TASK_PP(16'h16060,4);
TASK_PP(16'h16061,4);
TASK_PP(16'h16062,4);
TASK_PP(16'h16063,4);
TASK_PP(16'h16064,4);
TASK_PP(16'h16065,4);
TASK_PP(16'h16066,4);
TASK_PP(16'h16067,4);
TASK_PP(16'h16068,4);
TASK_PP(16'h16069,4);
TASK_PP(16'h1606A,4);
TASK_PP(16'h1606B,4);
TASK_PP(16'h1606C,4);
TASK_PP(16'h1606D,4);
TASK_PP(16'h1606E,4);
TASK_PP(16'h1606F,4);
TASK_PP(16'h16070,4);
TASK_PP(16'h16071,4);
TASK_PP(16'h16072,4);
TASK_PP(16'h16073,4);
TASK_PP(16'h16074,4);
TASK_PP(16'h16075,4);
TASK_PP(16'h16076,4);
TASK_PP(16'h16077,4);
TASK_PP(16'h16078,4);
TASK_PP(16'h16079,4);
TASK_PP(16'h1607A,4);
TASK_PP(16'h1607B,4);
TASK_PP(16'h1607C,4);
TASK_PP(16'h1607D,4);
TASK_PP(16'h1607E,4);
TASK_PP(16'h1607F,4);
TASK_PP(16'h16080,4);
TASK_PP(16'h16081,4);
TASK_PP(16'h16082,4);
TASK_PP(16'h16083,4);
TASK_PP(16'h16084,4);
TASK_PP(16'h16085,4);
TASK_PP(16'h16086,4);
TASK_PP(16'h16087,4);
TASK_PP(16'h16088,4);
TASK_PP(16'h16089,4);
TASK_PP(16'h1608A,4);
TASK_PP(16'h1608B,4);
TASK_PP(16'h1608C,4);
TASK_PP(16'h1608D,4);
TASK_PP(16'h1608E,4);
TASK_PP(16'h1608F,4);
TASK_PP(16'h16090,4);
TASK_PP(16'h16091,4);
TASK_PP(16'h16092,4);
TASK_PP(16'h16093,4);
TASK_PP(16'h16094,4);
TASK_PP(16'h16095,4);
TASK_PP(16'h16096,4);
TASK_PP(16'h16097,4);
TASK_PP(16'h16098,4);
TASK_PP(16'h16099,4);
TASK_PP(16'h1609A,4);
TASK_PP(16'h1609B,4);
TASK_PP(16'h1609C,4);
TASK_PP(16'h1609D,4);
TASK_PP(16'h1609E,4);
TASK_PP(16'h1609F,4);
TASK_PP(16'h160A0,4);
TASK_PP(16'h160A1,4);
TASK_PP(16'h160A2,4);
TASK_PP(16'h160A3,4);
TASK_PP(16'h160A4,4);
TASK_PP(16'h160A5,4);
TASK_PP(16'h160A6,4);
TASK_PP(16'h160A7,4);
TASK_PP(16'h160A8,4);
TASK_PP(16'h160A9,4);
TASK_PP(16'h160AA,4);
TASK_PP(16'h160AB,4);
TASK_PP(16'h160AC,4);
TASK_PP(16'h160AD,4);
TASK_PP(16'h160AE,4);
TASK_PP(16'h160AF,4);
TASK_PP(16'h160B0,4);
TASK_PP(16'h160B1,4);
TASK_PP(16'h160B2,4);
TASK_PP(16'h160B3,4);
TASK_PP(16'h160B4,4);
TASK_PP(16'h160B5,4);
TASK_PP(16'h160B6,4);
TASK_PP(16'h160B7,4);
TASK_PP(16'h160B8,4);
TASK_PP(16'h160B9,4);
TASK_PP(16'h160BA,4);
TASK_PP(16'h160BB,4);
TASK_PP(16'h160BC,4);
TASK_PP(16'h160BD,4);
TASK_PP(16'h160BE,4);
TASK_PP(16'h160BF,4);
TASK_PP(16'h160C0,4);
TASK_PP(16'h160C1,4);
TASK_PP(16'h160C2,4);
TASK_PP(16'h160C3,4);
TASK_PP(16'h160C4,4);
TASK_PP(16'h160C5,4);
TASK_PP(16'h160C6,4);
TASK_PP(16'h160C7,4);
TASK_PP(16'h160C8,4);
TASK_PP(16'h160C9,4);
TASK_PP(16'h160CA,4);
TASK_PP(16'h160CB,4);
TASK_PP(16'h160CC,4);
TASK_PP(16'h160CD,4);
TASK_PP(16'h160CE,4);
TASK_PP(16'h160CF,4);
TASK_PP(16'h160D0,4);
TASK_PP(16'h160D1,4);
TASK_PP(16'h160D2,4);
TASK_PP(16'h160D3,4);
TASK_PP(16'h160D4,4);
TASK_PP(16'h160D5,4);
TASK_PP(16'h160D6,4);
TASK_PP(16'h160D7,4);
TASK_PP(16'h160D8,4);
TASK_PP(16'h160D9,4);
TASK_PP(16'h160DA,4);
TASK_PP(16'h160DB,4);
TASK_PP(16'h160DC,4);
TASK_PP(16'h160DD,4);
TASK_PP(16'h160DE,4);
TASK_PP(16'h160DF,4);
TASK_PP(16'h160E0,4);
TASK_PP(16'h160E1,4);
TASK_PP(16'h160E2,4);
TASK_PP(16'h160E3,4);
TASK_PP(16'h160E4,4);
TASK_PP(16'h160E5,4);
TASK_PP(16'h160E6,4);
TASK_PP(16'h160E7,4);
TASK_PP(16'h160E8,4);
TASK_PP(16'h160E9,4);
TASK_PP(16'h160EA,4);
TASK_PP(16'h160EB,4);
TASK_PP(16'h160EC,4);
TASK_PP(16'h160ED,4);
TASK_PP(16'h160EE,4);
TASK_PP(16'h160EF,4);
TASK_PP(16'h160F0,4);
TASK_PP(16'h160F1,4);
TASK_PP(16'h160F2,4);
TASK_PP(16'h160F3,4);
TASK_PP(16'h160F4,4);
TASK_PP(16'h160F5,4);
TASK_PP(16'h160F6,4);
TASK_PP(16'h160F7,4);
TASK_PP(16'h160F8,4);
TASK_PP(16'h160F9,4);
TASK_PP(16'h160FA,4);
TASK_PP(16'h160FB,4);
TASK_PP(16'h160FC,4);
TASK_PP(16'h160FD,4);
TASK_PP(16'h160FE,4);
TASK_PP(16'h160FF,4);
TASK_PP(16'h16100,4);
TASK_PP(16'h16101,4);
TASK_PP(16'h16102,4);
TASK_PP(16'h16103,4);
TASK_PP(16'h16104,4);
TASK_PP(16'h16105,4);
TASK_PP(16'h16106,4);
TASK_PP(16'h16107,4);
TASK_PP(16'h16108,4);
TASK_PP(16'h16109,4);
TASK_PP(16'h1610A,4);
TASK_PP(16'h1610B,4);
TASK_PP(16'h1610C,4);
TASK_PP(16'h1610D,4);
TASK_PP(16'h1610E,4);
TASK_PP(16'h1610F,4);
TASK_PP(16'h16110,4);
TASK_PP(16'h16111,4);
TASK_PP(16'h16112,4);
TASK_PP(16'h16113,4);
TASK_PP(16'h16114,4);
TASK_PP(16'h16115,4);
TASK_PP(16'h16116,4);
TASK_PP(16'h16117,4);
TASK_PP(16'h16118,4);
TASK_PP(16'h16119,4);
TASK_PP(16'h1611A,4);
TASK_PP(16'h1611B,4);
TASK_PP(16'h1611C,4);
TASK_PP(16'h1611D,4);
TASK_PP(16'h1611E,4);
TASK_PP(16'h1611F,4);
TASK_PP(16'h16120,4);
TASK_PP(16'h16121,4);
TASK_PP(16'h16122,4);
TASK_PP(16'h16123,4);
TASK_PP(16'h16124,4);
TASK_PP(16'h16125,4);
TASK_PP(16'h16126,4);
TASK_PP(16'h16127,4);
TASK_PP(16'h16128,4);
TASK_PP(16'h16129,4);
TASK_PP(16'h1612A,4);
TASK_PP(16'h1612B,4);
TASK_PP(16'h1612C,4);
TASK_PP(16'h1612D,4);
TASK_PP(16'h1612E,4);
TASK_PP(16'h1612F,4);
TASK_PP(16'h16130,4);
TASK_PP(16'h16131,4);
TASK_PP(16'h16132,4);
TASK_PP(16'h16133,4);
TASK_PP(16'h16134,4);
TASK_PP(16'h16135,4);
TASK_PP(16'h16136,4);
TASK_PP(16'h16137,4);
TASK_PP(16'h16138,4);
TASK_PP(16'h16139,4);
TASK_PP(16'h1613A,4);
TASK_PP(16'h1613B,4);
TASK_PP(16'h1613C,4);
TASK_PP(16'h1613D,4);
TASK_PP(16'h1613E,4);
TASK_PP(16'h1613F,4);
TASK_PP(16'h16140,4);
TASK_PP(16'h16141,4);
TASK_PP(16'h16142,4);
TASK_PP(16'h16143,4);
TASK_PP(16'h16144,4);
TASK_PP(16'h16145,4);
TASK_PP(16'h16146,4);
TASK_PP(16'h16147,4);
TASK_PP(16'h16148,4);
TASK_PP(16'h16149,4);
TASK_PP(16'h1614A,4);
TASK_PP(16'h1614B,4);
TASK_PP(16'h1614C,4);
TASK_PP(16'h1614D,4);
TASK_PP(16'h1614E,4);
TASK_PP(16'h1614F,4);
TASK_PP(16'h16150,4);
TASK_PP(16'h16151,4);
TASK_PP(16'h16152,4);
TASK_PP(16'h16153,4);
TASK_PP(16'h16154,4);
TASK_PP(16'h16155,4);
TASK_PP(16'h16156,4);
TASK_PP(16'h16157,4);
TASK_PP(16'h16158,4);
TASK_PP(16'h16159,4);
TASK_PP(16'h1615A,4);
TASK_PP(16'h1615B,4);
TASK_PP(16'h1615C,4);
TASK_PP(16'h1615D,4);
TASK_PP(16'h1615E,4);
TASK_PP(16'h1615F,4);
TASK_PP(16'h16160,4);
TASK_PP(16'h16161,4);
TASK_PP(16'h16162,4);
TASK_PP(16'h16163,4);
TASK_PP(16'h16164,4);
TASK_PP(16'h16165,4);
TASK_PP(16'h16166,4);
TASK_PP(16'h16167,4);
TASK_PP(16'h16168,4);
TASK_PP(16'h16169,4);
TASK_PP(16'h1616A,4);
TASK_PP(16'h1616B,4);
TASK_PP(16'h1616C,4);
TASK_PP(16'h1616D,4);
TASK_PP(16'h1616E,4);
TASK_PP(16'h1616F,4);
TASK_PP(16'h16170,4);
TASK_PP(16'h16171,4);
TASK_PP(16'h16172,4);
TASK_PP(16'h16173,4);
TASK_PP(16'h16174,4);
TASK_PP(16'h16175,4);
TASK_PP(16'h16176,4);
TASK_PP(16'h16177,4);
TASK_PP(16'h16178,4);
TASK_PP(16'h16179,4);
TASK_PP(16'h1617A,4);
TASK_PP(16'h1617B,4);
TASK_PP(16'h1617C,4);
TASK_PP(16'h1617D,4);
TASK_PP(16'h1617E,4);
TASK_PP(16'h1617F,4);
TASK_PP(16'h16180,4);
TASK_PP(16'h16181,4);
TASK_PP(16'h16182,4);
TASK_PP(16'h16183,4);
TASK_PP(16'h16184,4);
TASK_PP(16'h16185,4);
TASK_PP(16'h16186,4);
TASK_PP(16'h16187,4);
TASK_PP(16'h16188,4);
TASK_PP(16'h16189,4);
TASK_PP(16'h1618A,4);
TASK_PP(16'h1618B,4);
TASK_PP(16'h1618C,4);
TASK_PP(16'h1618D,4);
TASK_PP(16'h1618E,4);
TASK_PP(16'h1618F,4);
TASK_PP(16'h16190,4);
TASK_PP(16'h16191,4);
TASK_PP(16'h16192,4);
TASK_PP(16'h16193,4);
TASK_PP(16'h16194,4);
TASK_PP(16'h16195,4);
TASK_PP(16'h16196,4);
TASK_PP(16'h16197,4);
TASK_PP(16'h16198,4);
TASK_PP(16'h16199,4);
TASK_PP(16'h1619A,4);
TASK_PP(16'h1619B,4);
TASK_PP(16'h1619C,4);
TASK_PP(16'h1619D,4);
TASK_PP(16'h1619E,4);
TASK_PP(16'h1619F,4);
TASK_PP(16'h161A0,4);
TASK_PP(16'h161A1,4);
TASK_PP(16'h161A2,4);
TASK_PP(16'h161A3,4);
TASK_PP(16'h161A4,4);
TASK_PP(16'h161A5,4);
TASK_PP(16'h161A6,4);
TASK_PP(16'h161A7,4);
TASK_PP(16'h161A8,4);
TASK_PP(16'h161A9,4);
TASK_PP(16'h161AA,4);
TASK_PP(16'h161AB,4);
TASK_PP(16'h161AC,4);
TASK_PP(16'h161AD,4);
TASK_PP(16'h161AE,4);
TASK_PP(16'h161AF,4);
TASK_PP(16'h161B0,4);
TASK_PP(16'h161B1,4);
TASK_PP(16'h161B2,4);
TASK_PP(16'h161B3,4);
TASK_PP(16'h161B4,4);
TASK_PP(16'h161B5,4);
TASK_PP(16'h161B6,4);
TASK_PP(16'h161B7,4);
TASK_PP(16'h161B8,4);
TASK_PP(16'h161B9,4);
TASK_PP(16'h161BA,4);
TASK_PP(16'h161BB,4);
TASK_PP(16'h161BC,4);
TASK_PP(16'h161BD,4);
TASK_PP(16'h161BE,4);
TASK_PP(16'h161BF,4);
TASK_PP(16'h161C0,4);
TASK_PP(16'h161C1,4);
TASK_PP(16'h161C2,4);
TASK_PP(16'h161C3,4);
TASK_PP(16'h161C4,4);
TASK_PP(16'h161C5,4);
TASK_PP(16'h161C6,4);
TASK_PP(16'h161C7,4);
TASK_PP(16'h161C8,4);
TASK_PP(16'h161C9,4);
TASK_PP(16'h161CA,4);
TASK_PP(16'h161CB,4);
TASK_PP(16'h161CC,4);
TASK_PP(16'h161CD,4);
TASK_PP(16'h161CE,4);
TASK_PP(16'h161CF,4);
TASK_PP(16'h161D0,4);
TASK_PP(16'h161D1,4);
TASK_PP(16'h161D2,4);
TASK_PP(16'h161D3,4);
TASK_PP(16'h161D4,4);
TASK_PP(16'h161D5,4);
TASK_PP(16'h161D6,4);
TASK_PP(16'h161D7,4);
TASK_PP(16'h161D8,4);
TASK_PP(16'h161D9,4);
TASK_PP(16'h161DA,4);
TASK_PP(16'h161DB,4);
TASK_PP(16'h161DC,4);
TASK_PP(16'h161DD,4);
TASK_PP(16'h161DE,4);
TASK_PP(16'h161DF,4);
TASK_PP(16'h161E0,4);
TASK_PP(16'h161E1,4);
TASK_PP(16'h161E2,4);
TASK_PP(16'h161E3,4);
TASK_PP(16'h161E4,4);
TASK_PP(16'h161E5,4);
TASK_PP(16'h161E6,4);
TASK_PP(16'h161E7,4);
TASK_PP(16'h161E8,4);
TASK_PP(16'h161E9,4);
TASK_PP(16'h161EA,4);
TASK_PP(16'h161EB,4);
TASK_PP(16'h161EC,4);
TASK_PP(16'h161ED,4);
TASK_PP(16'h161EE,4);
TASK_PP(16'h161EF,4);
TASK_PP(16'h161F0,4);
TASK_PP(16'h161F1,4);
TASK_PP(16'h161F2,4);
TASK_PP(16'h161F3,4);
TASK_PP(16'h161F4,4);
TASK_PP(16'h161F5,4);
TASK_PP(16'h161F6,4);
TASK_PP(16'h161F7,4);
TASK_PP(16'h161F8,4);
TASK_PP(16'h161F9,4);
TASK_PP(16'h161FA,4);
TASK_PP(16'h161FB,4);
TASK_PP(16'h161FC,4);
TASK_PP(16'h161FD,4);
TASK_PP(16'h161FE,4);
TASK_PP(16'h161FF,4);
TASK_PP(16'h16200,4);
TASK_PP(16'h16201,4);
TASK_PP(16'h16202,4);
TASK_PP(16'h16203,4);
TASK_PP(16'h16204,4);
TASK_PP(16'h16205,4);
TASK_PP(16'h16206,4);
TASK_PP(16'h16207,4);
TASK_PP(16'h16208,4);
TASK_PP(16'h16209,4);
TASK_PP(16'h1620A,4);
TASK_PP(16'h1620B,4);
TASK_PP(16'h1620C,4);
TASK_PP(16'h1620D,4);
TASK_PP(16'h1620E,4);
TASK_PP(16'h1620F,4);
TASK_PP(16'h16210,4);
TASK_PP(16'h16211,4);
TASK_PP(16'h16212,4);
TASK_PP(16'h16213,4);
TASK_PP(16'h16214,4);
TASK_PP(16'h16215,4);
TASK_PP(16'h16216,4);
TASK_PP(16'h16217,4);
TASK_PP(16'h16218,4);
TASK_PP(16'h16219,4);
TASK_PP(16'h1621A,4);
TASK_PP(16'h1621B,4);
TASK_PP(16'h1621C,4);
TASK_PP(16'h1621D,4);
TASK_PP(16'h1621E,4);
TASK_PP(16'h1621F,4);
TASK_PP(16'h16220,4);
TASK_PP(16'h16221,4);
TASK_PP(16'h16222,4);
TASK_PP(16'h16223,4);
TASK_PP(16'h16224,4);
TASK_PP(16'h16225,4);
TASK_PP(16'h16226,4);
TASK_PP(16'h16227,4);
TASK_PP(16'h16228,4);
TASK_PP(16'h16229,4);
TASK_PP(16'h1622A,4);
TASK_PP(16'h1622B,4);
TASK_PP(16'h1622C,4);
TASK_PP(16'h1622D,4);
TASK_PP(16'h1622E,4);
TASK_PP(16'h1622F,4);
TASK_PP(16'h16230,4);
TASK_PP(16'h16231,4);
TASK_PP(16'h16232,4);
TASK_PP(16'h16233,4);
TASK_PP(16'h16234,4);
TASK_PP(16'h16235,4);
TASK_PP(16'h16236,4);
TASK_PP(16'h16237,4);
TASK_PP(16'h16238,4);
TASK_PP(16'h16239,4);
TASK_PP(16'h1623A,4);
TASK_PP(16'h1623B,4);
TASK_PP(16'h1623C,4);
TASK_PP(16'h1623D,4);
TASK_PP(16'h1623E,4);
TASK_PP(16'h1623F,4);
TASK_PP(16'h16240,4);
TASK_PP(16'h16241,4);
TASK_PP(16'h16242,4);
TASK_PP(16'h16243,4);
TASK_PP(16'h16244,4);
TASK_PP(16'h16245,4);
TASK_PP(16'h16246,4);
TASK_PP(16'h16247,4);
TASK_PP(16'h16248,4);
TASK_PP(16'h16249,4);
TASK_PP(16'h1624A,4);
TASK_PP(16'h1624B,4);
TASK_PP(16'h1624C,4);
TASK_PP(16'h1624D,4);
TASK_PP(16'h1624E,4);
TASK_PP(16'h1624F,4);
TASK_PP(16'h16250,4);
TASK_PP(16'h16251,4);
TASK_PP(16'h16252,4);
TASK_PP(16'h16253,4);
TASK_PP(16'h16254,4);
TASK_PP(16'h16255,4);
TASK_PP(16'h16256,4);
TASK_PP(16'h16257,4);
TASK_PP(16'h16258,4);
TASK_PP(16'h16259,4);
TASK_PP(16'h1625A,4);
TASK_PP(16'h1625B,4);
TASK_PP(16'h1625C,4);
TASK_PP(16'h1625D,4);
TASK_PP(16'h1625E,4);
TASK_PP(16'h1625F,4);
TASK_PP(16'h16260,4);
TASK_PP(16'h16261,4);
TASK_PP(16'h16262,4);
TASK_PP(16'h16263,4);
TASK_PP(16'h16264,4);
TASK_PP(16'h16265,4);
TASK_PP(16'h16266,4);
TASK_PP(16'h16267,4);
TASK_PP(16'h16268,4);
TASK_PP(16'h16269,4);
TASK_PP(16'h1626A,4);
TASK_PP(16'h1626B,4);
TASK_PP(16'h1626C,4);
TASK_PP(16'h1626D,4);
TASK_PP(16'h1626E,4);
TASK_PP(16'h1626F,4);
TASK_PP(16'h16270,4);
TASK_PP(16'h16271,4);
TASK_PP(16'h16272,4);
TASK_PP(16'h16273,4);
TASK_PP(16'h16274,4);
TASK_PP(16'h16275,4);
TASK_PP(16'h16276,4);
TASK_PP(16'h16277,4);
TASK_PP(16'h16278,4);
TASK_PP(16'h16279,4);
TASK_PP(16'h1627A,4);
TASK_PP(16'h1627B,4);
TASK_PP(16'h1627C,4);
TASK_PP(16'h1627D,4);
TASK_PP(16'h1627E,4);
TASK_PP(16'h1627F,4);
TASK_PP(16'h16280,4);
TASK_PP(16'h16281,4);
TASK_PP(16'h16282,4);
TASK_PP(16'h16283,4);
TASK_PP(16'h16284,4);
TASK_PP(16'h16285,4);
TASK_PP(16'h16286,4);
TASK_PP(16'h16287,4);
TASK_PP(16'h16288,4);
TASK_PP(16'h16289,4);
TASK_PP(16'h1628A,4);
TASK_PP(16'h1628B,4);
TASK_PP(16'h1628C,4);
TASK_PP(16'h1628D,4);
TASK_PP(16'h1628E,4);
TASK_PP(16'h1628F,4);
TASK_PP(16'h16290,4);
TASK_PP(16'h16291,4);
TASK_PP(16'h16292,4);
TASK_PP(16'h16293,4);
TASK_PP(16'h16294,4);
TASK_PP(16'h16295,4);
TASK_PP(16'h16296,4);
TASK_PP(16'h16297,4);
TASK_PP(16'h16298,4);
TASK_PP(16'h16299,4);
TASK_PP(16'h1629A,4);
TASK_PP(16'h1629B,4);
TASK_PP(16'h1629C,4);
TASK_PP(16'h1629D,4);
TASK_PP(16'h1629E,4);
TASK_PP(16'h1629F,4);
TASK_PP(16'h162A0,4);
TASK_PP(16'h162A1,4);
TASK_PP(16'h162A2,4);
TASK_PP(16'h162A3,4);
TASK_PP(16'h162A4,4);
TASK_PP(16'h162A5,4);
TASK_PP(16'h162A6,4);
TASK_PP(16'h162A7,4);
TASK_PP(16'h162A8,4);
TASK_PP(16'h162A9,4);
TASK_PP(16'h162AA,4);
TASK_PP(16'h162AB,4);
TASK_PP(16'h162AC,4);
TASK_PP(16'h162AD,4);
TASK_PP(16'h162AE,4);
TASK_PP(16'h162AF,4);
TASK_PP(16'h162B0,4);
TASK_PP(16'h162B1,4);
TASK_PP(16'h162B2,4);
TASK_PP(16'h162B3,4);
TASK_PP(16'h162B4,4);
TASK_PP(16'h162B5,4);
TASK_PP(16'h162B6,4);
TASK_PP(16'h162B7,4);
TASK_PP(16'h162B8,4);
TASK_PP(16'h162B9,4);
TASK_PP(16'h162BA,4);
TASK_PP(16'h162BB,4);
TASK_PP(16'h162BC,4);
TASK_PP(16'h162BD,4);
TASK_PP(16'h162BE,4);
TASK_PP(16'h162BF,4);
TASK_PP(16'h162C0,4);
TASK_PP(16'h162C1,4);
TASK_PP(16'h162C2,4);
TASK_PP(16'h162C3,4);
TASK_PP(16'h162C4,4);
TASK_PP(16'h162C5,4);
TASK_PP(16'h162C6,4);
TASK_PP(16'h162C7,4);
TASK_PP(16'h162C8,4);
TASK_PP(16'h162C9,4);
TASK_PP(16'h162CA,4);
TASK_PP(16'h162CB,4);
TASK_PP(16'h162CC,4);
TASK_PP(16'h162CD,4);
TASK_PP(16'h162CE,4);
TASK_PP(16'h162CF,4);
TASK_PP(16'h162D0,4);
TASK_PP(16'h162D1,4);
TASK_PP(16'h162D2,4);
TASK_PP(16'h162D3,4);
TASK_PP(16'h162D4,4);
TASK_PP(16'h162D5,4);
TASK_PP(16'h162D6,4);
TASK_PP(16'h162D7,4);
TASK_PP(16'h162D8,4);
TASK_PP(16'h162D9,4);
TASK_PP(16'h162DA,4);
TASK_PP(16'h162DB,4);
TASK_PP(16'h162DC,4);
TASK_PP(16'h162DD,4);
TASK_PP(16'h162DE,4);
TASK_PP(16'h162DF,4);
TASK_PP(16'h162E0,4);
TASK_PP(16'h162E1,4);
TASK_PP(16'h162E2,4);
TASK_PP(16'h162E3,4);
TASK_PP(16'h162E4,4);
TASK_PP(16'h162E5,4);
TASK_PP(16'h162E6,4);
TASK_PP(16'h162E7,4);
TASK_PP(16'h162E8,4);
TASK_PP(16'h162E9,4);
TASK_PP(16'h162EA,4);
TASK_PP(16'h162EB,4);
TASK_PP(16'h162EC,4);
TASK_PP(16'h162ED,4);
TASK_PP(16'h162EE,4);
TASK_PP(16'h162EF,4);
TASK_PP(16'h162F0,4);
TASK_PP(16'h162F1,4);
TASK_PP(16'h162F2,4);
TASK_PP(16'h162F3,4);
TASK_PP(16'h162F4,4);
TASK_PP(16'h162F5,4);
TASK_PP(16'h162F6,4);
TASK_PP(16'h162F7,4);
TASK_PP(16'h162F8,4);
TASK_PP(16'h162F9,4);
TASK_PP(16'h162FA,4);
TASK_PP(16'h162FB,4);
TASK_PP(16'h162FC,4);
TASK_PP(16'h162FD,4);
TASK_PP(16'h162FE,4);
TASK_PP(16'h162FF,4);
TASK_PP(16'h16300,4);
TASK_PP(16'h16301,4);
TASK_PP(16'h16302,4);
TASK_PP(16'h16303,4);
TASK_PP(16'h16304,4);
TASK_PP(16'h16305,4);
TASK_PP(16'h16306,4);
TASK_PP(16'h16307,4);
TASK_PP(16'h16308,4);
TASK_PP(16'h16309,4);
TASK_PP(16'h1630A,4);
TASK_PP(16'h1630B,4);
TASK_PP(16'h1630C,4);
TASK_PP(16'h1630D,4);
TASK_PP(16'h1630E,4);
TASK_PP(16'h1630F,4);
TASK_PP(16'h16310,4);
TASK_PP(16'h16311,4);
TASK_PP(16'h16312,4);
TASK_PP(16'h16313,4);
TASK_PP(16'h16314,4);
TASK_PP(16'h16315,4);
TASK_PP(16'h16316,4);
TASK_PP(16'h16317,4);
TASK_PP(16'h16318,4);
TASK_PP(16'h16319,4);
TASK_PP(16'h1631A,4);
TASK_PP(16'h1631B,4);
TASK_PP(16'h1631C,4);
TASK_PP(16'h1631D,4);
TASK_PP(16'h1631E,4);
TASK_PP(16'h1631F,4);
TASK_PP(16'h16320,4);
TASK_PP(16'h16321,4);
TASK_PP(16'h16322,4);
TASK_PP(16'h16323,4);
TASK_PP(16'h16324,4);
TASK_PP(16'h16325,4);
TASK_PP(16'h16326,4);
TASK_PP(16'h16327,4);
TASK_PP(16'h16328,4);
TASK_PP(16'h16329,4);
TASK_PP(16'h1632A,4);
TASK_PP(16'h1632B,4);
TASK_PP(16'h1632C,4);
TASK_PP(16'h1632D,4);
TASK_PP(16'h1632E,4);
TASK_PP(16'h1632F,4);
TASK_PP(16'h16330,4);
TASK_PP(16'h16331,4);
TASK_PP(16'h16332,4);
TASK_PP(16'h16333,4);
TASK_PP(16'h16334,4);
TASK_PP(16'h16335,4);
TASK_PP(16'h16336,4);
TASK_PP(16'h16337,4);
TASK_PP(16'h16338,4);
TASK_PP(16'h16339,4);
TASK_PP(16'h1633A,4);
TASK_PP(16'h1633B,4);
TASK_PP(16'h1633C,4);
TASK_PP(16'h1633D,4);
TASK_PP(16'h1633E,4);
TASK_PP(16'h1633F,4);
TASK_PP(16'h16340,4);
TASK_PP(16'h16341,4);
TASK_PP(16'h16342,4);
TASK_PP(16'h16343,4);
TASK_PP(16'h16344,4);
TASK_PP(16'h16345,4);
TASK_PP(16'h16346,4);
TASK_PP(16'h16347,4);
TASK_PP(16'h16348,4);
TASK_PP(16'h16349,4);
TASK_PP(16'h1634A,4);
TASK_PP(16'h1634B,4);
TASK_PP(16'h1634C,4);
TASK_PP(16'h1634D,4);
TASK_PP(16'h1634E,4);
TASK_PP(16'h1634F,4);
TASK_PP(16'h16350,4);
TASK_PP(16'h16351,4);
TASK_PP(16'h16352,4);
TASK_PP(16'h16353,4);
TASK_PP(16'h16354,4);
TASK_PP(16'h16355,4);
TASK_PP(16'h16356,4);
TASK_PP(16'h16357,4);
TASK_PP(16'h16358,4);
TASK_PP(16'h16359,4);
TASK_PP(16'h1635A,4);
TASK_PP(16'h1635B,4);
TASK_PP(16'h1635C,4);
TASK_PP(16'h1635D,4);
TASK_PP(16'h1635E,4);
TASK_PP(16'h1635F,4);
TASK_PP(16'h16360,4);
TASK_PP(16'h16361,4);
TASK_PP(16'h16362,4);
TASK_PP(16'h16363,4);
TASK_PP(16'h16364,4);
TASK_PP(16'h16365,4);
TASK_PP(16'h16366,4);
TASK_PP(16'h16367,4);
TASK_PP(16'h16368,4);
TASK_PP(16'h16369,4);
TASK_PP(16'h1636A,4);
TASK_PP(16'h1636B,4);
TASK_PP(16'h1636C,4);
TASK_PP(16'h1636D,4);
TASK_PP(16'h1636E,4);
TASK_PP(16'h1636F,4);
TASK_PP(16'h16370,4);
TASK_PP(16'h16371,4);
TASK_PP(16'h16372,4);
TASK_PP(16'h16373,4);
TASK_PP(16'h16374,4);
TASK_PP(16'h16375,4);
TASK_PP(16'h16376,4);
TASK_PP(16'h16377,4);
TASK_PP(16'h16378,4);
TASK_PP(16'h16379,4);
TASK_PP(16'h1637A,4);
TASK_PP(16'h1637B,4);
TASK_PP(16'h1637C,4);
TASK_PP(16'h1637D,4);
TASK_PP(16'h1637E,4);
TASK_PP(16'h1637F,4);
TASK_PP(16'h16380,4);
TASK_PP(16'h16381,4);
TASK_PP(16'h16382,4);
TASK_PP(16'h16383,4);
TASK_PP(16'h16384,4);
TASK_PP(16'h16385,4);
TASK_PP(16'h16386,4);
TASK_PP(16'h16387,4);
TASK_PP(16'h16388,4);
TASK_PP(16'h16389,4);
TASK_PP(16'h1638A,4);
TASK_PP(16'h1638B,4);
TASK_PP(16'h1638C,4);
TASK_PP(16'h1638D,4);
TASK_PP(16'h1638E,4);
TASK_PP(16'h1638F,4);
TASK_PP(16'h16390,4);
TASK_PP(16'h16391,4);
TASK_PP(16'h16392,4);
TASK_PP(16'h16393,4);
TASK_PP(16'h16394,4);
TASK_PP(16'h16395,4);
TASK_PP(16'h16396,4);
TASK_PP(16'h16397,4);
TASK_PP(16'h16398,4);
TASK_PP(16'h16399,4);
TASK_PP(16'h1639A,4);
TASK_PP(16'h1639B,4);
TASK_PP(16'h1639C,4);
TASK_PP(16'h1639D,4);
TASK_PP(16'h1639E,4);
TASK_PP(16'h1639F,4);
TASK_PP(16'h163A0,4);
TASK_PP(16'h163A1,4);
TASK_PP(16'h163A2,4);
TASK_PP(16'h163A3,4);
TASK_PP(16'h163A4,4);
TASK_PP(16'h163A5,4);
TASK_PP(16'h163A6,4);
TASK_PP(16'h163A7,4);
TASK_PP(16'h163A8,4);
TASK_PP(16'h163A9,4);
TASK_PP(16'h163AA,4);
TASK_PP(16'h163AB,4);
TASK_PP(16'h163AC,4);
TASK_PP(16'h163AD,4);
TASK_PP(16'h163AE,4);
TASK_PP(16'h163AF,4);
TASK_PP(16'h163B0,4);
TASK_PP(16'h163B1,4);
TASK_PP(16'h163B2,4);
TASK_PP(16'h163B3,4);
TASK_PP(16'h163B4,4);
TASK_PP(16'h163B5,4);
TASK_PP(16'h163B6,4);
TASK_PP(16'h163B7,4);
TASK_PP(16'h163B8,4);
TASK_PP(16'h163B9,4);
TASK_PP(16'h163BA,4);
TASK_PP(16'h163BB,4);
TASK_PP(16'h163BC,4);
TASK_PP(16'h163BD,4);
TASK_PP(16'h163BE,4);
TASK_PP(16'h163BF,4);
TASK_PP(16'h163C0,4);
TASK_PP(16'h163C1,4);
TASK_PP(16'h163C2,4);
TASK_PP(16'h163C3,4);
TASK_PP(16'h163C4,4);
TASK_PP(16'h163C5,4);
TASK_PP(16'h163C6,4);
TASK_PP(16'h163C7,4);
TASK_PP(16'h163C8,4);
TASK_PP(16'h163C9,4);
TASK_PP(16'h163CA,4);
TASK_PP(16'h163CB,4);
TASK_PP(16'h163CC,4);
TASK_PP(16'h163CD,4);
TASK_PP(16'h163CE,4);
TASK_PP(16'h163CF,4);
TASK_PP(16'h163D0,4);
TASK_PP(16'h163D1,4);
TASK_PP(16'h163D2,4);
TASK_PP(16'h163D3,4);
TASK_PP(16'h163D4,4);
TASK_PP(16'h163D5,4);
TASK_PP(16'h163D6,4);
TASK_PP(16'h163D7,4);
TASK_PP(16'h163D8,4);
TASK_PP(16'h163D9,4);
TASK_PP(16'h163DA,4);
TASK_PP(16'h163DB,4);
TASK_PP(16'h163DC,4);
TASK_PP(16'h163DD,4);
TASK_PP(16'h163DE,4);
TASK_PP(16'h163DF,4);
TASK_PP(16'h163E0,4);
TASK_PP(16'h163E1,4);
TASK_PP(16'h163E2,4);
TASK_PP(16'h163E3,4);
TASK_PP(16'h163E4,4);
TASK_PP(16'h163E5,4);
TASK_PP(16'h163E6,4);
TASK_PP(16'h163E7,4);
TASK_PP(16'h163E8,4);
TASK_PP(16'h163E9,4);
TASK_PP(16'h163EA,4);
TASK_PP(16'h163EB,4);
TASK_PP(16'h163EC,4);
TASK_PP(16'h163ED,4);
TASK_PP(16'h163EE,4);
TASK_PP(16'h163EF,4);
TASK_PP(16'h163F0,4);
TASK_PP(16'h163F1,4);
TASK_PP(16'h163F2,4);
TASK_PP(16'h163F3,4);
TASK_PP(16'h163F4,4);
TASK_PP(16'h163F5,4);
TASK_PP(16'h163F6,4);
TASK_PP(16'h163F7,4);
TASK_PP(16'h163F8,4);
TASK_PP(16'h163F9,4);
TASK_PP(16'h163FA,4);
TASK_PP(16'h163FB,4);
TASK_PP(16'h163FC,4);
TASK_PP(16'h163FD,4);
TASK_PP(16'h163FE,4);
TASK_PP(16'h163FF,4);
TASK_PP(16'h16400,4);
TASK_PP(16'h16401,4);
TASK_PP(16'h16402,4);
TASK_PP(16'h16403,4);
TASK_PP(16'h16404,4);
TASK_PP(16'h16405,4);
TASK_PP(16'h16406,4);
TASK_PP(16'h16407,4);
TASK_PP(16'h16408,4);
TASK_PP(16'h16409,4);
TASK_PP(16'h1640A,4);
TASK_PP(16'h1640B,4);
TASK_PP(16'h1640C,4);
TASK_PP(16'h1640D,4);
TASK_PP(16'h1640E,4);
TASK_PP(16'h1640F,4);
TASK_PP(16'h16410,4);
TASK_PP(16'h16411,4);
TASK_PP(16'h16412,4);
TASK_PP(16'h16413,4);
TASK_PP(16'h16414,4);
TASK_PP(16'h16415,4);
TASK_PP(16'h16416,4);
TASK_PP(16'h16417,4);
TASK_PP(16'h16418,4);
TASK_PP(16'h16419,4);
TASK_PP(16'h1641A,4);
TASK_PP(16'h1641B,4);
TASK_PP(16'h1641C,4);
TASK_PP(16'h1641D,4);
TASK_PP(16'h1641E,4);
TASK_PP(16'h1641F,4);
TASK_PP(16'h16420,4);
TASK_PP(16'h16421,4);
TASK_PP(16'h16422,4);
TASK_PP(16'h16423,4);
TASK_PP(16'h16424,4);
TASK_PP(16'h16425,4);
TASK_PP(16'h16426,4);
TASK_PP(16'h16427,4);
TASK_PP(16'h16428,4);
TASK_PP(16'h16429,4);
TASK_PP(16'h1642A,4);
TASK_PP(16'h1642B,4);
TASK_PP(16'h1642C,4);
TASK_PP(16'h1642D,4);
TASK_PP(16'h1642E,4);
TASK_PP(16'h1642F,4);
TASK_PP(16'h16430,4);
TASK_PP(16'h16431,4);
TASK_PP(16'h16432,4);
TASK_PP(16'h16433,4);
TASK_PP(16'h16434,4);
TASK_PP(16'h16435,4);
TASK_PP(16'h16436,4);
TASK_PP(16'h16437,4);
TASK_PP(16'h16438,4);
TASK_PP(16'h16439,4);
TASK_PP(16'h1643A,4);
TASK_PP(16'h1643B,4);
TASK_PP(16'h1643C,4);
TASK_PP(16'h1643D,4);
TASK_PP(16'h1643E,4);
TASK_PP(16'h1643F,4);
TASK_PP(16'h16440,4);
TASK_PP(16'h16441,4);
TASK_PP(16'h16442,4);
TASK_PP(16'h16443,4);
TASK_PP(16'h16444,4);
TASK_PP(16'h16445,4);
TASK_PP(16'h16446,4);
TASK_PP(16'h16447,4);
TASK_PP(16'h16448,4);
TASK_PP(16'h16449,4);
TASK_PP(16'h1644A,4);
TASK_PP(16'h1644B,4);
TASK_PP(16'h1644C,4);
TASK_PP(16'h1644D,4);
TASK_PP(16'h1644E,4);
TASK_PP(16'h1644F,4);
TASK_PP(16'h16450,4);
TASK_PP(16'h16451,4);
TASK_PP(16'h16452,4);
TASK_PP(16'h16453,4);
TASK_PP(16'h16454,4);
TASK_PP(16'h16455,4);
TASK_PP(16'h16456,4);
TASK_PP(16'h16457,4);
TASK_PP(16'h16458,4);
TASK_PP(16'h16459,4);
TASK_PP(16'h1645A,4);
TASK_PP(16'h1645B,4);
TASK_PP(16'h1645C,4);
TASK_PP(16'h1645D,4);
TASK_PP(16'h1645E,4);
TASK_PP(16'h1645F,4);
TASK_PP(16'h16460,4);
TASK_PP(16'h16461,4);
TASK_PP(16'h16462,4);
TASK_PP(16'h16463,4);
TASK_PP(16'h16464,4);
TASK_PP(16'h16465,4);
TASK_PP(16'h16466,4);
TASK_PP(16'h16467,4);
TASK_PP(16'h16468,4);
TASK_PP(16'h16469,4);
TASK_PP(16'h1646A,4);
TASK_PP(16'h1646B,4);
TASK_PP(16'h1646C,4);
TASK_PP(16'h1646D,4);
TASK_PP(16'h1646E,4);
TASK_PP(16'h1646F,4);
TASK_PP(16'h16470,4);
TASK_PP(16'h16471,4);
TASK_PP(16'h16472,4);
TASK_PP(16'h16473,4);
TASK_PP(16'h16474,4);
TASK_PP(16'h16475,4);
TASK_PP(16'h16476,4);
TASK_PP(16'h16477,4);
TASK_PP(16'h16478,4);
TASK_PP(16'h16479,4);
TASK_PP(16'h1647A,4);
TASK_PP(16'h1647B,4);
TASK_PP(16'h1647C,4);
TASK_PP(16'h1647D,4);
TASK_PP(16'h1647E,4);
TASK_PP(16'h1647F,4);
TASK_PP(16'h16480,4);
TASK_PP(16'h16481,4);
TASK_PP(16'h16482,4);
TASK_PP(16'h16483,4);
TASK_PP(16'h16484,4);
TASK_PP(16'h16485,4);
TASK_PP(16'h16486,4);
TASK_PP(16'h16487,4);
TASK_PP(16'h16488,4);
TASK_PP(16'h16489,4);
TASK_PP(16'h1648A,4);
TASK_PP(16'h1648B,4);
TASK_PP(16'h1648C,4);
TASK_PP(16'h1648D,4);
TASK_PP(16'h1648E,4);
TASK_PP(16'h1648F,4);
TASK_PP(16'h16490,4);
TASK_PP(16'h16491,4);
TASK_PP(16'h16492,4);
TASK_PP(16'h16493,4);
TASK_PP(16'h16494,4);
TASK_PP(16'h16495,4);
TASK_PP(16'h16496,4);
TASK_PP(16'h16497,4);
TASK_PP(16'h16498,4);
TASK_PP(16'h16499,4);
TASK_PP(16'h1649A,4);
TASK_PP(16'h1649B,4);
TASK_PP(16'h1649C,4);
TASK_PP(16'h1649D,4);
TASK_PP(16'h1649E,4);
TASK_PP(16'h1649F,4);
TASK_PP(16'h164A0,4);
TASK_PP(16'h164A1,4);
TASK_PP(16'h164A2,4);
TASK_PP(16'h164A3,4);
TASK_PP(16'h164A4,4);
TASK_PP(16'h164A5,4);
TASK_PP(16'h164A6,4);
TASK_PP(16'h164A7,4);
TASK_PP(16'h164A8,4);
TASK_PP(16'h164A9,4);
TASK_PP(16'h164AA,4);
TASK_PP(16'h164AB,4);
TASK_PP(16'h164AC,4);
TASK_PP(16'h164AD,4);
TASK_PP(16'h164AE,4);
TASK_PP(16'h164AF,4);
TASK_PP(16'h164B0,4);
TASK_PP(16'h164B1,4);
TASK_PP(16'h164B2,4);
TASK_PP(16'h164B3,4);
TASK_PP(16'h164B4,4);
TASK_PP(16'h164B5,4);
TASK_PP(16'h164B6,4);
TASK_PP(16'h164B7,4);
TASK_PP(16'h164B8,4);
TASK_PP(16'h164B9,4);
TASK_PP(16'h164BA,4);
TASK_PP(16'h164BB,4);
TASK_PP(16'h164BC,4);
TASK_PP(16'h164BD,4);
TASK_PP(16'h164BE,4);
TASK_PP(16'h164BF,4);
TASK_PP(16'h164C0,4);
TASK_PP(16'h164C1,4);
TASK_PP(16'h164C2,4);
TASK_PP(16'h164C3,4);
TASK_PP(16'h164C4,4);
TASK_PP(16'h164C5,4);
TASK_PP(16'h164C6,4);
TASK_PP(16'h164C7,4);
TASK_PP(16'h164C8,4);
TASK_PP(16'h164C9,4);
TASK_PP(16'h164CA,4);
TASK_PP(16'h164CB,4);
TASK_PP(16'h164CC,4);
TASK_PP(16'h164CD,4);
TASK_PP(16'h164CE,4);
TASK_PP(16'h164CF,4);
TASK_PP(16'h164D0,4);
TASK_PP(16'h164D1,4);
TASK_PP(16'h164D2,4);
TASK_PP(16'h164D3,4);
TASK_PP(16'h164D4,4);
TASK_PP(16'h164D5,4);
TASK_PP(16'h164D6,4);
TASK_PP(16'h164D7,4);
TASK_PP(16'h164D8,4);
TASK_PP(16'h164D9,4);
TASK_PP(16'h164DA,4);
TASK_PP(16'h164DB,4);
TASK_PP(16'h164DC,4);
TASK_PP(16'h164DD,4);
TASK_PP(16'h164DE,4);
TASK_PP(16'h164DF,4);
TASK_PP(16'h164E0,4);
TASK_PP(16'h164E1,4);
TASK_PP(16'h164E2,4);
TASK_PP(16'h164E3,4);
TASK_PP(16'h164E4,4);
TASK_PP(16'h164E5,4);
TASK_PP(16'h164E6,4);
TASK_PP(16'h164E7,4);
TASK_PP(16'h164E8,4);
TASK_PP(16'h164E9,4);
TASK_PP(16'h164EA,4);
TASK_PP(16'h164EB,4);
TASK_PP(16'h164EC,4);
TASK_PP(16'h164ED,4);
TASK_PP(16'h164EE,4);
TASK_PP(16'h164EF,4);
TASK_PP(16'h164F0,4);
TASK_PP(16'h164F1,4);
TASK_PP(16'h164F2,4);
TASK_PP(16'h164F3,4);
TASK_PP(16'h164F4,4);
TASK_PP(16'h164F5,4);
TASK_PP(16'h164F6,4);
TASK_PP(16'h164F7,4);
TASK_PP(16'h164F8,4);
TASK_PP(16'h164F9,4);
TASK_PP(16'h164FA,4);
TASK_PP(16'h164FB,4);
TASK_PP(16'h164FC,4);
TASK_PP(16'h164FD,4);
TASK_PP(16'h164FE,4);
TASK_PP(16'h164FF,4);
TASK_PP(16'h16500,4);
TASK_PP(16'h16501,4);
TASK_PP(16'h16502,4);
TASK_PP(16'h16503,4);
TASK_PP(16'h16504,4);
TASK_PP(16'h16505,4);
TASK_PP(16'h16506,4);
TASK_PP(16'h16507,4);
TASK_PP(16'h16508,4);
TASK_PP(16'h16509,4);
TASK_PP(16'h1650A,4);
TASK_PP(16'h1650B,4);
TASK_PP(16'h1650C,4);
TASK_PP(16'h1650D,4);
TASK_PP(16'h1650E,4);
TASK_PP(16'h1650F,4);
TASK_PP(16'h16510,4);
TASK_PP(16'h16511,4);
TASK_PP(16'h16512,4);
TASK_PP(16'h16513,4);
TASK_PP(16'h16514,4);
TASK_PP(16'h16515,4);
TASK_PP(16'h16516,4);
TASK_PP(16'h16517,4);
TASK_PP(16'h16518,4);
TASK_PP(16'h16519,4);
TASK_PP(16'h1651A,4);
TASK_PP(16'h1651B,4);
TASK_PP(16'h1651C,4);
TASK_PP(16'h1651D,4);
TASK_PP(16'h1651E,4);
TASK_PP(16'h1651F,4);
TASK_PP(16'h16520,4);
TASK_PP(16'h16521,4);
TASK_PP(16'h16522,4);
TASK_PP(16'h16523,4);
TASK_PP(16'h16524,4);
TASK_PP(16'h16525,4);
TASK_PP(16'h16526,4);
TASK_PP(16'h16527,4);
TASK_PP(16'h16528,4);
TASK_PP(16'h16529,4);
TASK_PP(16'h1652A,4);
TASK_PP(16'h1652B,4);
TASK_PP(16'h1652C,4);
TASK_PP(16'h1652D,4);
TASK_PP(16'h1652E,4);
TASK_PP(16'h1652F,4);
TASK_PP(16'h16530,4);
TASK_PP(16'h16531,4);
TASK_PP(16'h16532,4);
TASK_PP(16'h16533,4);
TASK_PP(16'h16534,4);
TASK_PP(16'h16535,4);
TASK_PP(16'h16536,4);
TASK_PP(16'h16537,4);
TASK_PP(16'h16538,4);
TASK_PP(16'h16539,4);
TASK_PP(16'h1653A,4);
TASK_PP(16'h1653B,4);
TASK_PP(16'h1653C,4);
TASK_PP(16'h1653D,4);
TASK_PP(16'h1653E,4);
TASK_PP(16'h1653F,4);
TASK_PP(16'h16540,4);
TASK_PP(16'h16541,4);
TASK_PP(16'h16542,4);
TASK_PP(16'h16543,4);
TASK_PP(16'h16544,4);
TASK_PP(16'h16545,4);
TASK_PP(16'h16546,4);
TASK_PP(16'h16547,4);
TASK_PP(16'h16548,4);
TASK_PP(16'h16549,4);
TASK_PP(16'h1654A,4);
TASK_PP(16'h1654B,4);
TASK_PP(16'h1654C,4);
TASK_PP(16'h1654D,4);
TASK_PP(16'h1654E,4);
TASK_PP(16'h1654F,4);
TASK_PP(16'h16550,4);
TASK_PP(16'h16551,4);
TASK_PP(16'h16552,4);
TASK_PP(16'h16553,4);
TASK_PP(16'h16554,4);
TASK_PP(16'h16555,4);
TASK_PP(16'h16556,4);
TASK_PP(16'h16557,4);
TASK_PP(16'h16558,4);
TASK_PP(16'h16559,4);
TASK_PP(16'h1655A,4);
TASK_PP(16'h1655B,4);
TASK_PP(16'h1655C,4);
TASK_PP(16'h1655D,4);
TASK_PP(16'h1655E,4);
TASK_PP(16'h1655F,4);
TASK_PP(16'h16560,4);
TASK_PP(16'h16561,4);
TASK_PP(16'h16562,4);
TASK_PP(16'h16563,4);
TASK_PP(16'h16564,4);
TASK_PP(16'h16565,4);
TASK_PP(16'h16566,4);
TASK_PP(16'h16567,4);
TASK_PP(16'h16568,4);
TASK_PP(16'h16569,4);
TASK_PP(16'h1656A,4);
TASK_PP(16'h1656B,4);
TASK_PP(16'h1656C,4);
TASK_PP(16'h1656D,4);
TASK_PP(16'h1656E,4);
TASK_PP(16'h1656F,4);
TASK_PP(16'h16570,4);
TASK_PP(16'h16571,4);
TASK_PP(16'h16572,4);
TASK_PP(16'h16573,4);
TASK_PP(16'h16574,4);
TASK_PP(16'h16575,4);
TASK_PP(16'h16576,4);
TASK_PP(16'h16577,4);
TASK_PP(16'h16578,4);
TASK_PP(16'h16579,4);
TASK_PP(16'h1657A,4);
TASK_PP(16'h1657B,4);
TASK_PP(16'h1657C,4);
TASK_PP(16'h1657D,4);
TASK_PP(16'h1657E,4);
TASK_PP(16'h1657F,4);
TASK_PP(16'h16580,4);
TASK_PP(16'h16581,4);
TASK_PP(16'h16582,4);
TASK_PP(16'h16583,4);
TASK_PP(16'h16584,4);
TASK_PP(16'h16585,4);
TASK_PP(16'h16586,4);
TASK_PP(16'h16587,4);
TASK_PP(16'h16588,4);
TASK_PP(16'h16589,4);
TASK_PP(16'h1658A,4);
TASK_PP(16'h1658B,4);
TASK_PP(16'h1658C,4);
TASK_PP(16'h1658D,4);
TASK_PP(16'h1658E,4);
TASK_PP(16'h1658F,4);
TASK_PP(16'h16590,4);
TASK_PP(16'h16591,4);
TASK_PP(16'h16592,4);
TASK_PP(16'h16593,4);
TASK_PP(16'h16594,4);
TASK_PP(16'h16595,4);
TASK_PP(16'h16596,4);
TASK_PP(16'h16597,4);
TASK_PP(16'h16598,4);
TASK_PP(16'h16599,4);
TASK_PP(16'h1659A,4);
TASK_PP(16'h1659B,4);
TASK_PP(16'h1659C,4);
TASK_PP(16'h1659D,4);
TASK_PP(16'h1659E,4);
TASK_PP(16'h1659F,4);
TASK_PP(16'h165A0,4);
TASK_PP(16'h165A1,4);
TASK_PP(16'h165A2,4);
TASK_PP(16'h165A3,4);
TASK_PP(16'h165A4,4);
TASK_PP(16'h165A5,4);
TASK_PP(16'h165A6,4);
TASK_PP(16'h165A7,4);
TASK_PP(16'h165A8,4);
TASK_PP(16'h165A9,4);
TASK_PP(16'h165AA,4);
TASK_PP(16'h165AB,4);
TASK_PP(16'h165AC,4);
TASK_PP(16'h165AD,4);
TASK_PP(16'h165AE,4);
TASK_PP(16'h165AF,4);
TASK_PP(16'h165B0,4);
TASK_PP(16'h165B1,4);
TASK_PP(16'h165B2,4);
TASK_PP(16'h165B3,4);
TASK_PP(16'h165B4,4);
TASK_PP(16'h165B5,4);
TASK_PP(16'h165B6,4);
TASK_PP(16'h165B7,4);
TASK_PP(16'h165B8,4);
TASK_PP(16'h165B9,4);
TASK_PP(16'h165BA,4);
TASK_PP(16'h165BB,4);
TASK_PP(16'h165BC,4);
TASK_PP(16'h165BD,4);
TASK_PP(16'h165BE,4);
TASK_PP(16'h165BF,4);
TASK_PP(16'h165C0,4);
TASK_PP(16'h165C1,4);
TASK_PP(16'h165C2,4);
TASK_PP(16'h165C3,4);
TASK_PP(16'h165C4,4);
TASK_PP(16'h165C5,4);
TASK_PP(16'h165C6,4);
TASK_PP(16'h165C7,4);
TASK_PP(16'h165C8,4);
TASK_PP(16'h165C9,4);
TASK_PP(16'h165CA,4);
TASK_PP(16'h165CB,4);
TASK_PP(16'h165CC,4);
TASK_PP(16'h165CD,4);
TASK_PP(16'h165CE,4);
TASK_PP(16'h165CF,4);
TASK_PP(16'h165D0,4);
TASK_PP(16'h165D1,4);
TASK_PP(16'h165D2,4);
TASK_PP(16'h165D3,4);
TASK_PP(16'h165D4,4);
TASK_PP(16'h165D5,4);
TASK_PP(16'h165D6,4);
TASK_PP(16'h165D7,4);
TASK_PP(16'h165D8,4);
TASK_PP(16'h165D9,4);
TASK_PP(16'h165DA,4);
TASK_PP(16'h165DB,4);
TASK_PP(16'h165DC,4);
TASK_PP(16'h165DD,4);
TASK_PP(16'h165DE,4);
TASK_PP(16'h165DF,4);
TASK_PP(16'h165E0,4);
TASK_PP(16'h165E1,4);
TASK_PP(16'h165E2,4);
TASK_PP(16'h165E3,4);
TASK_PP(16'h165E4,4);
TASK_PP(16'h165E5,4);
TASK_PP(16'h165E6,4);
TASK_PP(16'h165E7,4);
TASK_PP(16'h165E8,4);
TASK_PP(16'h165E9,4);
TASK_PP(16'h165EA,4);
TASK_PP(16'h165EB,4);
TASK_PP(16'h165EC,4);
TASK_PP(16'h165ED,4);
TASK_PP(16'h165EE,4);
TASK_PP(16'h165EF,4);
TASK_PP(16'h165F0,4);
TASK_PP(16'h165F1,4);
TASK_PP(16'h165F2,4);
TASK_PP(16'h165F3,4);
TASK_PP(16'h165F4,4);
TASK_PP(16'h165F5,4);
TASK_PP(16'h165F6,4);
TASK_PP(16'h165F7,4);
TASK_PP(16'h165F8,4);
TASK_PP(16'h165F9,4);
TASK_PP(16'h165FA,4);
TASK_PP(16'h165FB,4);
TASK_PP(16'h165FC,4);
TASK_PP(16'h165FD,4);
TASK_PP(16'h165FE,4);
TASK_PP(16'h165FF,4);
TASK_PP(16'h16600,4);
TASK_PP(16'h16601,4);
TASK_PP(16'h16602,4);
TASK_PP(16'h16603,4);
TASK_PP(16'h16604,4);
TASK_PP(16'h16605,4);
TASK_PP(16'h16606,4);
TASK_PP(16'h16607,4);
TASK_PP(16'h16608,4);
TASK_PP(16'h16609,4);
TASK_PP(16'h1660A,4);
TASK_PP(16'h1660B,4);
TASK_PP(16'h1660C,4);
TASK_PP(16'h1660D,4);
TASK_PP(16'h1660E,4);
TASK_PP(16'h1660F,4);
TASK_PP(16'h16610,4);
TASK_PP(16'h16611,4);
TASK_PP(16'h16612,4);
TASK_PP(16'h16613,4);
TASK_PP(16'h16614,4);
TASK_PP(16'h16615,4);
TASK_PP(16'h16616,4);
TASK_PP(16'h16617,4);
TASK_PP(16'h16618,4);
TASK_PP(16'h16619,4);
TASK_PP(16'h1661A,4);
TASK_PP(16'h1661B,4);
TASK_PP(16'h1661C,4);
TASK_PP(16'h1661D,4);
TASK_PP(16'h1661E,4);
TASK_PP(16'h1661F,4);
TASK_PP(16'h16620,4);
TASK_PP(16'h16621,4);
TASK_PP(16'h16622,4);
TASK_PP(16'h16623,4);
TASK_PP(16'h16624,4);
TASK_PP(16'h16625,4);
TASK_PP(16'h16626,4);
TASK_PP(16'h16627,4);
TASK_PP(16'h16628,4);
TASK_PP(16'h16629,4);
TASK_PP(16'h1662A,4);
TASK_PP(16'h1662B,4);
TASK_PP(16'h1662C,4);
TASK_PP(16'h1662D,4);
TASK_PP(16'h1662E,4);
TASK_PP(16'h1662F,4);
TASK_PP(16'h16630,4);
TASK_PP(16'h16631,4);
TASK_PP(16'h16632,4);
TASK_PP(16'h16633,4);
TASK_PP(16'h16634,4);
TASK_PP(16'h16635,4);
TASK_PP(16'h16636,4);
TASK_PP(16'h16637,4);
TASK_PP(16'h16638,4);
TASK_PP(16'h16639,4);
TASK_PP(16'h1663A,4);
TASK_PP(16'h1663B,4);
TASK_PP(16'h1663C,4);
TASK_PP(16'h1663D,4);
TASK_PP(16'h1663E,4);
TASK_PP(16'h1663F,4);
TASK_PP(16'h16640,4);
TASK_PP(16'h16641,4);
TASK_PP(16'h16642,4);
TASK_PP(16'h16643,4);
TASK_PP(16'h16644,4);
TASK_PP(16'h16645,4);
TASK_PP(16'h16646,4);
TASK_PP(16'h16647,4);
TASK_PP(16'h16648,4);
TASK_PP(16'h16649,4);
TASK_PP(16'h1664A,4);
TASK_PP(16'h1664B,4);
TASK_PP(16'h1664C,4);
TASK_PP(16'h1664D,4);
TASK_PP(16'h1664E,4);
TASK_PP(16'h1664F,4);
TASK_PP(16'h16650,4);
TASK_PP(16'h16651,4);
TASK_PP(16'h16652,4);
TASK_PP(16'h16653,4);
TASK_PP(16'h16654,4);
TASK_PP(16'h16655,4);
TASK_PP(16'h16656,4);
TASK_PP(16'h16657,4);
TASK_PP(16'h16658,4);
TASK_PP(16'h16659,4);
TASK_PP(16'h1665A,4);
TASK_PP(16'h1665B,4);
TASK_PP(16'h1665C,4);
TASK_PP(16'h1665D,4);
TASK_PP(16'h1665E,4);
TASK_PP(16'h1665F,4);
TASK_PP(16'h16660,4);
TASK_PP(16'h16661,4);
TASK_PP(16'h16662,4);
TASK_PP(16'h16663,4);
TASK_PP(16'h16664,4);
TASK_PP(16'h16665,4);
TASK_PP(16'h16666,4);
TASK_PP(16'h16667,4);
TASK_PP(16'h16668,4);
TASK_PP(16'h16669,4);
TASK_PP(16'h1666A,4);
TASK_PP(16'h1666B,4);
TASK_PP(16'h1666C,4);
TASK_PP(16'h1666D,4);
TASK_PP(16'h1666E,4);
TASK_PP(16'h1666F,4);
TASK_PP(16'h16670,4);
TASK_PP(16'h16671,4);
TASK_PP(16'h16672,4);
TASK_PP(16'h16673,4);
TASK_PP(16'h16674,4);
TASK_PP(16'h16675,4);
TASK_PP(16'h16676,4);
TASK_PP(16'h16677,4);
TASK_PP(16'h16678,4);
TASK_PP(16'h16679,4);
TASK_PP(16'h1667A,4);
TASK_PP(16'h1667B,4);
TASK_PP(16'h1667C,4);
TASK_PP(16'h1667D,4);
TASK_PP(16'h1667E,4);
TASK_PP(16'h1667F,4);
TASK_PP(16'h16680,4);
TASK_PP(16'h16681,4);
TASK_PP(16'h16682,4);
TASK_PP(16'h16683,4);
TASK_PP(16'h16684,4);
TASK_PP(16'h16685,4);
TASK_PP(16'h16686,4);
TASK_PP(16'h16687,4);
TASK_PP(16'h16688,4);
TASK_PP(16'h16689,4);
TASK_PP(16'h1668A,4);
TASK_PP(16'h1668B,4);
TASK_PP(16'h1668C,4);
TASK_PP(16'h1668D,4);
TASK_PP(16'h1668E,4);
TASK_PP(16'h1668F,4);
TASK_PP(16'h16690,4);
TASK_PP(16'h16691,4);
TASK_PP(16'h16692,4);
TASK_PP(16'h16693,4);
TASK_PP(16'h16694,4);
TASK_PP(16'h16695,4);
TASK_PP(16'h16696,4);
TASK_PP(16'h16697,4);
TASK_PP(16'h16698,4);
TASK_PP(16'h16699,4);
TASK_PP(16'h1669A,4);
TASK_PP(16'h1669B,4);
TASK_PP(16'h1669C,4);
TASK_PP(16'h1669D,4);
TASK_PP(16'h1669E,4);
TASK_PP(16'h1669F,4);
TASK_PP(16'h166A0,4);
TASK_PP(16'h166A1,4);
TASK_PP(16'h166A2,4);
TASK_PP(16'h166A3,4);
TASK_PP(16'h166A4,4);
TASK_PP(16'h166A5,4);
TASK_PP(16'h166A6,4);
TASK_PP(16'h166A7,4);
TASK_PP(16'h166A8,4);
TASK_PP(16'h166A9,4);
TASK_PP(16'h166AA,4);
TASK_PP(16'h166AB,4);
TASK_PP(16'h166AC,4);
TASK_PP(16'h166AD,4);
TASK_PP(16'h166AE,4);
TASK_PP(16'h166AF,4);
TASK_PP(16'h166B0,4);
TASK_PP(16'h166B1,4);
TASK_PP(16'h166B2,4);
TASK_PP(16'h166B3,4);
TASK_PP(16'h166B4,4);
TASK_PP(16'h166B5,4);
TASK_PP(16'h166B6,4);
TASK_PP(16'h166B7,4);
TASK_PP(16'h166B8,4);
TASK_PP(16'h166B9,4);
TASK_PP(16'h166BA,4);
TASK_PP(16'h166BB,4);
TASK_PP(16'h166BC,4);
TASK_PP(16'h166BD,4);
TASK_PP(16'h166BE,4);
TASK_PP(16'h166BF,4);
TASK_PP(16'h166C0,4);
TASK_PP(16'h166C1,4);
TASK_PP(16'h166C2,4);
TASK_PP(16'h166C3,4);
TASK_PP(16'h166C4,4);
TASK_PP(16'h166C5,4);
TASK_PP(16'h166C6,4);
TASK_PP(16'h166C7,4);
TASK_PP(16'h166C8,4);
TASK_PP(16'h166C9,4);
TASK_PP(16'h166CA,4);
TASK_PP(16'h166CB,4);
TASK_PP(16'h166CC,4);
TASK_PP(16'h166CD,4);
TASK_PP(16'h166CE,4);
TASK_PP(16'h166CF,4);
TASK_PP(16'h166D0,4);
TASK_PP(16'h166D1,4);
TASK_PP(16'h166D2,4);
TASK_PP(16'h166D3,4);
TASK_PP(16'h166D4,4);
TASK_PP(16'h166D5,4);
TASK_PP(16'h166D6,4);
TASK_PP(16'h166D7,4);
TASK_PP(16'h166D8,4);
TASK_PP(16'h166D9,4);
TASK_PP(16'h166DA,4);
TASK_PP(16'h166DB,4);
TASK_PP(16'h166DC,4);
TASK_PP(16'h166DD,4);
TASK_PP(16'h166DE,4);
TASK_PP(16'h166DF,4);
TASK_PP(16'h166E0,4);
TASK_PP(16'h166E1,4);
TASK_PP(16'h166E2,4);
TASK_PP(16'h166E3,4);
TASK_PP(16'h166E4,4);
TASK_PP(16'h166E5,4);
TASK_PP(16'h166E6,4);
TASK_PP(16'h166E7,4);
TASK_PP(16'h166E8,4);
TASK_PP(16'h166E9,4);
TASK_PP(16'h166EA,4);
TASK_PP(16'h166EB,4);
TASK_PP(16'h166EC,4);
TASK_PP(16'h166ED,4);
TASK_PP(16'h166EE,4);
TASK_PP(16'h166EF,4);
TASK_PP(16'h166F0,4);
TASK_PP(16'h166F1,4);
TASK_PP(16'h166F2,4);
TASK_PP(16'h166F3,4);
TASK_PP(16'h166F4,4);
TASK_PP(16'h166F5,4);
TASK_PP(16'h166F6,4);
TASK_PP(16'h166F7,4);
TASK_PP(16'h166F8,4);
TASK_PP(16'h166F9,4);
TASK_PP(16'h166FA,4);
TASK_PP(16'h166FB,4);
TASK_PP(16'h166FC,4);
TASK_PP(16'h166FD,4);
TASK_PP(16'h166FE,4);
TASK_PP(16'h166FF,4);
TASK_PP(16'h16700,4);
TASK_PP(16'h16701,4);
TASK_PP(16'h16702,4);
TASK_PP(16'h16703,4);
TASK_PP(16'h16704,4);
TASK_PP(16'h16705,4);
TASK_PP(16'h16706,4);
TASK_PP(16'h16707,4);
TASK_PP(16'h16708,4);
TASK_PP(16'h16709,4);
TASK_PP(16'h1670A,4);
TASK_PP(16'h1670B,4);
TASK_PP(16'h1670C,4);
TASK_PP(16'h1670D,4);
TASK_PP(16'h1670E,4);
TASK_PP(16'h1670F,4);
TASK_PP(16'h16710,4);
TASK_PP(16'h16711,4);
TASK_PP(16'h16712,4);
TASK_PP(16'h16713,4);
TASK_PP(16'h16714,4);
TASK_PP(16'h16715,4);
TASK_PP(16'h16716,4);
TASK_PP(16'h16717,4);
TASK_PP(16'h16718,4);
TASK_PP(16'h16719,4);
TASK_PP(16'h1671A,4);
TASK_PP(16'h1671B,4);
TASK_PP(16'h1671C,4);
TASK_PP(16'h1671D,4);
TASK_PP(16'h1671E,4);
TASK_PP(16'h1671F,4);
TASK_PP(16'h16720,4);
TASK_PP(16'h16721,4);
TASK_PP(16'h16722,4);
TASK_PP(16'h16723,4);
TASK_PP(16'h16724,4);
TASK_PP(16'h16725,4);
TASK_PP(16'h16726,4);
TASK_PP(16'h16727,4);
TASK_PP(16'h16728,4);
TASK_PP(16'h16729,4);
TASK_PP(16'h1672A,4);
TASK_PP(16'h1672B,4);
TASK_PP(16'h1672C,4);
TASK_PP(16'h1672D,4);
TASK_PP(16'h1672E,4);
TASK_PP(16'h1672F,4);
TASK_PP(16'h16730,4);
TASK_PP(16'h16731,4);
TASK_PP(16'h16732,4);
TASK_PP(16'h16733,4);
TASK_PP(16'h16734,4);
TASK_PP(16'h16735,4);
TASK_PP(16'h16736,4);
TASK_PP(16'h16737,4);
TASK_PP(16'h16738,4);
TASK_PP(16'h16739,4);
TASK_PP(16'h1673A,4);
TASK_PP(16'h1673B,4);
TASK_PP(16'h1673C,4);
TASK_PP(16'h1673D,4);
TASK_PP(16'h1673E,4);
TASK_PP(16'h1673F,4);
TASK_PP(16'h16740,4);
TASK_PP(16'h16741,4);
TASK_PP(16'h16742,4);
TASK_PP(16'h16743,4);
TASK_PP(16'h16744,4);
TASK_PP(16'h16745,4);
TASK_PP(16'h16746,4);
TASK_PP(16'h16747,4);
TASK_PP(16'h16748,4);
TASK_PP(16'h16749,4);
TASK_PP(16'h1674A,4);
TASK_PP(16'h1674B,4);
TASK_PP(16'h1674C,4);
TASK_PP(16'h1674D,4);
TASK_PP(16'h1674E,4);
TASK_PP(16'h1674F,4);
TASK_PP(16'h16750,4);
TASK_PP(16'h16751,4);
TASK_PP(16'h16752,4);
TASK_PP(16'h16753,4);
TASK_PP(16'h16754,4);
TASK_PP(16'h16755,4);
TASK_PP(16'h16756,4);
TASK_PP(16'h16757,4);
TASK_PP(16'h16758,4);
TASK_PP(16'h16759,4);
TASK_PP(16'h1675A,4);
TASK_PP(16'h1675B,4);
TASK_PP(16'h1675C,4);
TASK_PP(16'h1675D,4);
TASK_PP(16'h1675E,4);
TASK_PP(16'h1675F,4);
TASK_PP(16'h16760,4);
TASK_PP(16'h16761,4);
TASK_PP(16'h16762,4);
TASK_PP(16'h16763,4);
TASK_PP(16'h16764,4);
TASK_PP(16'h16765,4);
TASK_PP(16'h16766,4);
TASK_PP(16'h16767,4);
TASK_PP(16'h16768,4);
TASK_PP(16'h16769,4);
TASK_PP(16'h1676A,4);
TASK_PP(16'h1676B,4);
TASK_PP(16'h1676C,4);
TASK_PP(16'h1676D,4);
TASK_PP(16'h1676E,4);
TASK_PP(16'h1676F,4);
TASK_PP(16'h16770,4);
TASK_PP(16'h16771,4);
TASK_PP(16'h16772,4);
TASK_PP(16'h16773,4);
TASK_PP(16'h16774,4);
TASK_PP(16'h16775,4);
TASK_PP(16'h16776,4);
TASK_PP(16'h16777,4);
TASK_PP(16'h16778,4);
TASK_PP(16'h16779,4);
TASK_PP(16'h1677A,4);
TASK_PP(16'h1677B,4);
TASK_PP(16'h1677C,4);
TASK_PP(16'h1677D,4);
TASK_PP(16'h1677E,4);
TASK_PP(16'h1677F,4);
TASK_PP(16'h16780,4);
TASK_PP(16'h16781,4);
TASK_PP(16'h16782,4);
TASK_PP(16'h16783,4);
TASK_PP(16'h16784,4);
TASK_PP(16'h16785,4);
TASK_PP(16'h16786,4);
TASK_PP(16'h16787,4);
TASK_PP(16'h16788,4);
TASK_PP(16'h16789,4);
TASK_PP(16'h1678A,4);
TASK_PP(16'h1678B,4);
TASK_PP(16'h1678C,4);
TASK_PP(16'h1678D,4);
TASK_PP(16'h1678E,4);
TASK_PP(16'h1678F,4);
TASK_PP(16'h16790,4);
TASK_PP(16'h16791,4);
TASK_PP(16'h16792,4);
TASK_PP(16'h16793,4);
TASK_PP(16'h16794,4);
TASK_PP(16'h16795,4);
TASK_PP(16'h16796,4);
TASK_PP(16'h16797,4);
TASK_PP(16'h16798,4);
TASK_PP(16'h16799,4);
TASK_PP(16'h1679A,4);
TASK_PP(16'h1679B,4);
TASK_PP(16'h1679C,4);
TASK_PP(16'h1679D,4);
TASK_PP(16'h1679E,4);
TASK_PP(16'h1679F,4);
TASK_PP(16'h167A0,4);
TASK_PP(16'h167A1,4);
TASK_PP(16'h167A2,4);
TASK_PP(16'h167A3,4);
TASK_PP(16'h167A4,4);
TASK_PP(16'h167A5,4);
TASK_PP(16'h167A6,4);
TASK_PP(16'h167A7,4);
TASK_PP(16'h167A8,4);
TASK_PP(16'h167A9,4);
TASK_PP(16'h167AA,4);
TASK_PP(16'h167AB,4);
TASK_PP(16'h167AC,4);
TASK_PP(16'h167AD,4);
TASK_PP(16'h167AE,4);
TASK_PP(16'h167AF,4);
TASK_PP(16'h167B0,4);
TASK_PP(16'h167B1,4);
TASK_PP(16'h167B2,4);
TASK_PP(16'h167B3,4);
TASK_PP(16'h167B4,4);
TASK_PP(16'h167B5,4);
TASK_PP(16'h167B6,4);
TASK_PP(16'h167B7,4);
TASK_PP(16'h167B8,4);
TASK_PP(16'h167B9,4);
TASK_PP(16'h167BA,4);
TASK_PP(16'h167BB,4);
TASK_PP(16'h167BC,4);
TASK_PP(16'h167BD,4);
TASK_PP(16'h167BE,4);
TASK_PP(16'h167BF,4);
TASK_PP(16'h167C0,4);
TASK_PP(16'h167C1,4);
TASK_PP(16'h167C2,4);
TASK_PP(16'h167C3,4);
TASK_PP(16'h167C4,4);
TASK_PP(16'h167C5,4);
TASK_PP(16'h167C6,4);
TASK_PP(16'h167C7,4);
TASK_PP(16'h167C8,4);
TASK_PP(16'h167C9,4);
TASK_PP(16'h167CA,4);
TASK_PP(16'h167CB,4);
TASK_PP(16'h167CC,4);
TASK_PP(16'h167CD,4);
TASK_PP(16'h167CE,4);
TASK_PP(16'h167CF,4);
TASK_PP(16'h167D0,4);
TASK_PP(16'h167D1,4);
TASK_PP(16'h167D2,4);
TASK_PP(16'h167D3,4);
TASK_PP(16'h167D4,4);
TASK_PP(16'h167D5,4);
TASK_PP(16'h167D6,4);
TASK_PP(16'h167D7,4);
TASK_PP(16'h167D8,4);
TASK_PP(16'h167D9,4);
TASK_PP(16'h167DA,4);
TASK_PP(16'h167DB,4);
TASK_PP(16'h167DC,4);
TASK_PP(16'h167DD,4);
TASK_PP(16'h167DE,4);
TASK_PP(16'h167DF,4);
TASK_PP(16'h167E0,4);
TASK_PP(16'h167E1,4);
TASK_PP(16'h167E2,4);
TASK_PP(16'h167E3,4);
TASK_PP(16'h167E4,4);
TASK_PP(16'h167E5,4);
TASK_PP(16'h167E6,4);
TASK_PP(16'h167E7,4);
TASK_PP(16'h167E8,4);
TASK_PP(16'h167E9,4);
TASK_PP(16'h167EA,4);
TASK_PP(16'h167EB,4);
TASK_PP(16'h167EC,4);
TASK_PP(16'h167ED,4);
TASK_PP(16'h167EE,4);
TASK_PP(16'h167EF,4);
TASK_PP(16'h167F0,4);
TASK_PP(16'h167F1,4);
TASK_PP(16'h167F2,4);
TASK_PP(16'h167F3,4);
TASK_PP(16'h167F4,4);
TASK_PP(16'h167F5,4);
TASK_PP(16'h167F6,4);
TASK_PP(16'h167F7,4);
TASK_PP(16'h167F8,4);
TASK_PP(16'h167F9,4);
TASK_PP(16'h167FA,4);
TASK_PP(16'h167FB,4);
TASK_PP(16'h167FC,4);
TASK_PP(16'h167FD,4);
TASK_PP(16'h167FE,4);
TASK_PP(16'h167FF,4);
TASK_PP(16'h16800,4);
TASK_PP(16'h16801,4);
TASK_PP(16'h16802,4);
TASK_PP(16'h16803,4);
TASK_PP(16'h16804,4);
TASK_PP(16'h16805,4);
TASK_PP(16'h16806,4);
TASK_PP(16'h16807,4);
TASK_PP(16'h16808,4);
TASK_PP(16'h16809,4);
TASK_PP(16'h1680A,4);
TASK_PP(16'h1680B,4);
TASK_PP(16'h1680C,4);
TASK_PP(16'h1680D,4);
TASK_PP(16'h1680E,4);
TASK_PP(16'h1680F,4);
TASK_PP(16'h16810,4);
TASK_PP(16'h16811,4);
TASK_PP(16'h16812,4);
TASK_PP(16'h16813,4);
TASK_PP(16'h16814,4);
TASK_PP(16'h16815,4);
TASK_PP(16'h16816,4);
TASK_PP(16'h16817,4);
TASK_PP(16'h16818,4);
TASK_PP(16'h16819,4);
TASK_PP(16'h1681A,4);
TASK_PP(16'h1681B,4);
TASK_PP(16'h1681C,4);
TASK_PP(16'h1681D,4);
TASK_PP(16'h1681E,4);
TASK_PP(16'h1681F,4);
TASK_PP(16'h16820,4);
TASK_PP(16'h16821,4);
TASK_PP(16'h16822,4);
TASK_PP(16'h16823,4);
TASK_PP(16'h16824,4);
TASK_PP(16'h16825,4);
TASK_PP(16'h16826,4);
TASK_PP(16'h16827,4);
TASK_PP(16'h16828,4);
TASK_PP(16'h16829,4);
TASK_PP(16'h1682A,4);
TASK_PP(16'h1682B,4);
TASK_PP(16'h1682C,4);
TASK_PP(16'h1682D,4);
TASK_PP(16'h1682E,4);
TASK_PP(16'h1682F,4);
TASK_PP(16'h16830,4);
TASK_PP(16'h16831,4);
TASK_PP(16'h16832,4);
TASK_PP(16'h16833,4);
TASK_PP(16'h16834,4);
TASK_PP(16'h16835,4);
TASK_PP(16'h16836,4);
TASK_PP(16'h16837,4);
TASK_PP(16'h16838,4);
TASK_PP(16'h16839,4);
TASK_PP(16'h1683A,4);
TASK_PP(16'h1683B,4);
TASK_PP(16'h1683C,4);
TASK_PP(16'h1683D,4);
TASK_PP(16'h1683E,4);
TASK_PP(16'h1683F,4);
TASK_PP(16'h16840,4);
TASK_PP(16'h16841,4);
TASK_PP(16'h16842,4);
TASK_PP(16'h16843,4);
TASK_PP(16'h16844,4);
TASK_PP(16'h16845,4);
TASK_PP(16'h16846,4);
TASK_PP(16'h16847,4);
TASK_PP(16'h16848,4);
TASK_PP(16'h16849,4);
TASK_PP(16'h1684A,4);
TASK_PP(16'h1684B,4);
TASK_PP(16'h1684C,4);
TASK_PP(16'h1684D,4);
TASK_PP(16'h1684E,4);
TASK_PP(16'h1684F,4);
TASK_PP(16'h16850,4);
TASK_PP(16'h16851,4);
TASK_PP(16'h16852,4);
TASK_PP(16'h16853,4);
TASK_PP(16'h16854,4);
TASK_PP(16'h16855,4);
TASK_PP(16'h16856,4);
TASK_PP(16'h16857,4);
TASK_PP(16'h16858,4);
TASK_PP(16'h16859,4);
TASK_PP(16'h1685A,4);
TASK_PP(16'h1685B,4);
TASK_PP(16'h1685C,4);
TASK_PP(16'h1685D,4);
TASK_PP(16'h1685E,4);
TASK_PP(16'h1685F,4);
TASK_PP(16'h16860,4);
TASK_PP(16'h16861,4);
TASK_PP(16'h16862,4);
TASK_PP(16'h16863,4);
TASK_PP(16'h16864,4);
TASK_PP(16'h16865,4);
TASK_PP(16'h16866,4);
TASK_PP(16'h16867,4);
TASK_PP(16'h16868,4);
TASK_PP(16'h16869,4);
TASK_PP(16'h1686A,4);
TASK_PP(16'h1686B,4);
TASK_PP(16'h1686C,4);
TASK_PP(16'h1686D,4);
TASK_PP(16'h1686E,4);
TASK_PP(16'h1686F,4);
TASK_PP(16'h16870,4);
TASK_PP(16'h16871,4);
TASK_PP(16'h16872,4);
TASK_PP(16'h16873,4);
TASK_PP(16'h16874,4);
TASK_PP(16'h16875,4);
TASK_PP(16'h16876,4);
TASK_PP(16'h16877,4);
TASK_PP(16'h16878,4);
TASK_PP(16'h16879,4);
TASK_PP(16'h1687A,4);
TASK_PP(16'h1687B,4);
TASK_PP(16'h1687C,4);
TASK_PP(16'h1687D,4);
TASK_PP(16'h1687E,4);
TASK_PP(16'h1687F,4);
TASK_PP(16'h16880,4);
TASK_PP(16'h16881,4);
TASK_PP(16'h16882,4);
TASK_PP(16'h16883,4);
TASK_PP(16'h16884,4);
TASK_PP(16'h16885,4);
TASK_PP(16'h16886,4);
TASK_PP(16'h16887,4);
TASK_PP(16'h16888,4);
TASK_PP(16'h16889,4);
TASK_PP(16'h1688A,4);
TASK_PP(16'h1688B,4);
TASK_PP(16'h1688C,4);
TASK_PP(16'h1688D,4);
TASK_PP(16'h1688E,4);
TASK_PP(16'h1688F,4);
TASK_PP(16'h16890,4);
TASK_PP(16'h16891,4);
TASK_PP(16'h16892,4);
TASK_PP(16'h16893,4);
TASK_PP(16'h16894,4);
TASK_PP(16'h16895,4);
TASK_PP(16'h16896,4);
TASK_PP(16'h16897,4);
TASK_PP(16'h16898,4);
TASK_PP(16'h16899,4);
TASK_PP(16'h1689A,4);
TASK_PP(16'h1689B,4);
TASK_PP(16'h1689C,4);
TASK_PP(16'h1689D,4);
TASK_PP(16'h1689E,4);
TASK_PP(16'h1689F,4);
TASK_PP(16'h168A0,4);
TASK_PP(16'h168A1,4);
TASK_PP(16'h168A2,4);
TASK_PP(16'h168A3,4);
TASK_PP(16'h168A4,4);
TASK_PP(16'h168A5,4);
TASK_PP(16'h168A6,4);
TASK_PP(16'h168A7,4);
TASK_PP(16'h168A8,4);
TASK_PP(16'h168A9,4);
TASK_PP(16'h168AA,4);
TASK_PP(16'h168AB,4);
TASK_PP(16'h168AC,4);
TASK_PP(16'h168AD,4);
TASK_PP(16'h168AE,4);
TASK_PP(16'h168AF,4);
TASK_PP(16'h168B0,4);
TASK_PP(16'h168B1,4);
TASK_PP(16'h168B2,4);
TASK_PP(16'h168B3,4);
TASK_PP(16'h168B4,4);
TASK_PP(16'h168B5,4);
TASK_PP(16'h168B6,4);
TASK_PP(16'h168B7,4);
TASK_PP(16'h168B8,4);
TASK_PP(16'h168B9,4);
TASK_PP(16'h168BA,4);
TASK_PP(16'h168BB,4);
TASK_PP(16'h168BC,4);
TASK_PP(16'h168BD,4);
TASK_PP(16'h168BE,4);
TASK_PP(16'h168BF,4);
TASK_PP(16'h168C0,4);
TASK_PP(16'h168C1,4);
TASK_PP(16'h168C2,4);
TASK_PP(16'h168C3,4);
TASK_PP(16'h168C4,4);
TASK_PP(16'h168C5,4);
TASK_PP(16'h168C6,4);
TASK_PP(16'h168C7,4);
TASK_PP(16'h168C8,4);
TASK_PP(16'h168C9,4);
TASK_PP(16'h168CA,4);
TASK_PP(16'h168CB,4);
TASK_PP(16'h168CC,4);
TASK_PP(16'h168CD,4);
TASK_PP(16'h168CE,4);
TASK_PP(16'h168CF,4);
TASK_PP(16'h168D0,4);
TASK_PP(16'h168D1,4);
TASK_PP(16'h168D2,4);
TASK_PP(16'h168D3,4);
TASK_PP(16'h168D4,4);
TASK_PP(16'h168D5,4);
TASK_PP(16'h168D6,4);
TASK_PP(16'h168D7,4);
TASK_PP(16'h168D8,4);
TASK_PP(16'h168D9,4);
TASK_PP(16'h168DA,4);
TASK_PP(16'h168DB,4);
TASK_PP(16'h168DC,4);
TASK_PP(16'h168DD,4);
TASK_PP(16'h168DE,4);
TASK_PP(16'h168DF,4);
TASK_PP(16'h168E0,4);
TASK_PP(16'h168E1,4);
TASK_PP(16'h168E2,4);
TASK_PP(16'h168E3,4);
TASK_PP(16'h168E4,4);
TASK_PP(16'h168E5,4);
TASK_PP(16'h168E6,4);
TASK_PP(16'h168E7,4);
TASK_PP(16'h168E8,4);
TASK_PP(16'h168E9,4);
TASK_PP(16'h168EA,4);
TASK_PP(16'h168EB,4);
TASK_PP(16'h168EC,4);
TASK_PP(16'h168ED,4);
TASK_PP(16'h168EE,4);
TASK_PP(16'h168EF,4);
TASK_PP(16'h168F0,4);
TASK_PP(16'h168F1,4);
TASK_PP(16'h168F2,4);
TASK_PP(16'h168F3,4);
TASK_PP(16'h168F4,4);
TASK_PP(16'h168F5,4);
TASK_PP(16'h168F6,4);
TASK_PP(16'h168F7,4);
TASK_PP(16'h168F8,4);
TASK_PP(16'h168F9,4);
TASK_PP(16'h168FA,4);
TASK_PP(16'h168FB,4);
TASK_PP(16'h168FC,4);
TASK_PP(16'h168FD,4);
TASK_PP(16'h168FE,4);
TASK_PP(16'h168FF,4);
TASK_PP(16'h16900,4);
TASK_PP(16'h16901,4);
TASK_PP(16'h16902,4);
TASK_PP(16'h16903,4);
TASK_PP(16'h16904,4);
TASK_PP(16'h16905,4);
TASK_PP(16'h16906,4);
TASK_PP(16'h16907,4);
TASK_PP(16'h16908,4);
TASK_PP(16'h16909,4);
TASK_PP(16'h1690A,4);
TASK_PP(16'h1690B,4);
TASK_PP(16'h1690C,4);
TASK_PP(16'h1690D,4);
TASK_PP(16'h1690E,4);
TASK_PP(16'h1690F,4);
TASK_PP(16'h16910,4);
TASK_PP(16'h16911,4);
TASK_PP(16'h16912,4);
TASK_PP(16'h16913,4);
TASK_PP(16'h16914,4);
TASK_PP(16'h16915,4);
TASK_PP(16'h16916,4);
TASK_PP(16'h16917,4);
TASK_PP(16'h16918,4);
TASK_PP(16'h16919,4);
TASK_PP(16'h1691A,4);
TASK_PP(16'h1691B,4);
TASK_PP(16'h1691C,4);
TASK_PP(16'h1691D,4);
TASK_PP(16'h1691E,4);
TASK_PP(16'h1691F,4);
TASK_PP(16'h16920,4);
TASK_PP(16'h16921,4);
TASK_PP(16'h16922,4);
TASK_PP(16'h16923,4);
TASK_PP(16'h16924,4);
TASK_PP(16'h16925,4);
TASK_PP(16'h16926,4);
TASK_PP(16'h16927,4);
TASK_PP(16'h16928,4);
TASK_PP(16'h16929,4);
TASK_PP(16'h1692A,4);
TASK_PP(16'h1692B,4);
TASK_PP(16'h1692C,4);
TASK_PP(16'h1692D,4);
TASK_PP(16'h1692E,4);
TASK_PP(16'h1692F,4);
TASK_PP(16'h16930,4);
TASK_PP(16'h16931,4);
TASK_PP(16'h16932,4);
TASK_PP(16'h16933,4);
TASK_PP(16'h16934,4);
TASK_PP(16'h16935,4);
TASK_PP(16'h16936,4);
TASK_PP(16'h16937,4);
TASK_PP(16'h16938,4);
TASK_PP(16'h16939,4);
TASK_PP(16'h1693A,4);
TASK_PP(16'h1693B,4);
TASK_PP(16'h1693C,4);
TASK_PP(16'h1693D,4);
TASK_PP(16'h1693E,4);
TASK_PP(16'h1693F,4);
TASK_PP(16'h16940,4);
TASK_PP(16'h16941,4);
TASK_PP(16'h16942,4);
TASK_PP(16'h16943,4);
TASK_PP(16'h16944,4);
TASK_PP(16'h16945,4);
TASK_PP(16'h16946,4);
TASK_PP(16'h16947,4);
TASK_PP(16'h16948,4);
TASK_PP(16'h16949,4);
TASK_PP(16'h1694A,4);
TASK_PP(16'h1694B,4);
TASK_PP(16'h1694C,4);
TASK_PP(16'h1694D,4);
TASK_PP(16'h1694E,4);
TASK_PP(16'h1694F,4);
TASK_PP(16'h16950,4);
TASK_PP(16'h16951,4);
TASK_PP(16'h16952,4);
TASK_PP(16'h16953,4);
TASK_PP(16'h16954,4);
TASK_PP(16'h16955,4);
TASK_PP(16'h16956,4);
TASK_PP(16'h16957,4);
TASK_PP(16'h16958,4);
TASK_PP(16'h16959,4);
TASK_PP(16'h1695A,4);
TASK_PP(16'h1695B,4);
TASK_PP(16'h1695C,4);
TASK_PP(16'h1695D,4);
TASK_PP(16'h1695E,4);
TASK_PP(16'h1695F,4);
TASK_PP(16'h16960,4);
TASK_PP(16'h16961,4);
TASK_PP(16'h16962,4);
TASK_PP(16'h16963,4);
TASK_PP(16'h16964,4);
TASK_PP(16'h16965,4);
TASK_PP(16'h16966,4);
TASK_PP(16'h16967,4);
TASK_PP(16'h16968,4);
TASK_PP(16'h16969,4);
TASK_PP(16'h1696A,4);
TASK_PP(16'h1696B,4);
TASK_PP(16'h1696C,4);
TASK_PP(16'h1696D,4);
TASK_PP(16'h1696E,4);
TASK_PP(16'h1696F,4);
TASK_PP(16'h16970,4);
TASK_PP(16'h16971,4);
TASK_PP(16'h16972,4);
TASK_PP(16'h16973,4);
TASK_PP(16'h16974,4);
TASK_PP(16'h16975,4);
TASK_PP(16'h16976,4);
TASK_PP(16'h16977,4);
TASK_PP(16'h16978,4);
TASK_PP(16'h16979,4);
TASK_PP(16'h1697A,4);
TASK_PP(16'h1697B,4);
TASK_PP(16'h1697C,4);
TASK_PP(16'h1697D,4);
TASK_PP(16'h1697E,4);
TASK_PP(16'h1697F,4);
TASK_PP(16'h16980,4);
TASK_PP(16'h16981,4);
TASK_PP(16'h16982,4);
TASK_PP(16'h16983,4);
TASK_PP(16'h16984,4);
TASK_PP(16'h16985,4);
TASK_PP(16'h16986,4);
TASK_PP(16'h16987,4);
TASK_PP(16'h16988,4);
TASK_PP(16'h16989,4);
TASK_PP(16'h1698A,4);
TASK_PP(16'h1698B,4);
TASK_PP(16'h1698C,4);
TASK_PP(16'h1698D,4);
TASK_PP(16'h1698E,4);
TASK_PP(16'h1698F,4);
TASK_PP(16'h16990,4);
TASK_PP(16'h16991,4);
TASK_PP(16'h16992,4);
TASK_PP(16'h16993,4);
TASK_PP(16'h16994,4);
TASK_PP(16'h16995,4);
TASK_PP(16'h16996,4);
TASK_PP(16'h16997,4);
TASK_PP(16'h16998,4);
TASK_PP(16'h16999,4);
TASK_PP(16'h1699A,4);
TASK_PP(16'h1699B,4);
TASK_PP(16'h1699C,4);
TASK_PP(16'h1699D,4);
TASK_PP(16'h1699E,4);
TASK_PP(16'h1699F,4);
TASK_PP(16'h169A0,4);
TASK_PP(16'h169A1,4);
TASK_PP(16'h169A2,4);
TASK_PP(16'h169A3,4);
TASK_PP(16'h169A4,4);
TASK_PP(16'h169A5,4);
TASK_PP(16'h169A6,4);
TASK_PP(16'h169A7,4);
TASK_PP(16'h169A8,4);
TASK_PP(16'h169A9,4);
TASK_PP(16'h169AA,4);
TASK_PP(16'h169AB,4);
TASK_PP(16'h169AC,4);
TASK_PP(16'h169AD,4);
TASK_PP(16'h169AE,4);
TASK_PP(16'h169AF,4);
TASK_PP(16'h169B0,4);
TASK_PP(16'h169B1,4);
TASK_PP(16'h169B2,4);
TASK_PP(16'h169B3,4);
TASK_PP(16'h169B4,4);
TASK_PP(16'h169B5,4);
TASK_PP(16'h169B6,4);
TASK_PP(16'h169B7,4);
TASK_PP(16'h169B8,4);
TASK_PP(16'h169B9,4);
TASK_PP(16'h169BA,4);
TASK_PP(16'h169BB,4);
TASK_PP(16'h169BC,4);
TASK_PP(16'h169BD,4);
TASK_PP(16'h169BE,4);
TASK_PP(16'h169BF,4);
TASK_PP(16'h169C0,4);
TASK_PP(16'h169C1,4);
TASK_PP(16'h169C2,4);
TASK_PP(16'h169C3,4);
TASK_PP(16'h169C4,4);
TASK_PP(16'h169C5,4);
TASK_PP(16'h169C6,4);
TASK_PP(16'h169C7,4);
TASK_PP(16'h169C8,4);
TASK_PP(16'h169C9,4);
TASK_PP(16'h169CA,4);
TASK_PP(16'h169CB,4);
TASK_PP(16'h169CC,4);
TASK_PP(16'h169CD,4);
TASK_PP(16'h169CE,4);
TASK_PP(16'h169CF,4);
TASK_PP(16'h169D0,4);
TASK_PP(16'h169D1,4);
TASK_PP(16'h169D2,4);
TASK_PP(16'h169D3,4);
TASK_PP(16'h169D4,4);
TASK_PP(16'h169D5,4);
TASK_PP(16'h169D6,4);
TASK_PP(16'h169D7,4);
TASK_PP(16'h169D8,4);
TASK_PP(16'h169D9,4);
TASK_PP(16'h169DA,4);
TASK_PP(16'h169DB,4);
TASK_PP(16'h169DC,4);
TASK_PP(16'h169DD,4);
TASK_PP(16'h169DE,4);
TASK_PP(16'h169DF,4);
TASK_PP(16'h169E0,4);
TASK_PP(16'h169E1,4);
TASK_PP(16'h169E2,4);
TASK_PP(16'h169E3,4);
TASK_PP(16'h169E4,4);
TASK_PP(16'h169E5,4);
TASK_PP(16'h169E6,4);
TASK_PP(16'h169E7,4);
TASK_PP(16'h169E8,4);
TASK_PP(16'h169E9,4);
TASK_PP(16'h169EA,4);
TASK_PP(16'h169EB,4);
TASK_PP(16'h169EC,4);
TASK_PP(16'h169ED,4);
TASK_PP(16'h169EE,4);
TASK_PP(16'h169EF,4);
TASK_PP(16'h169F0,4);
TASK_PP(16'h169F1,4);
TASK_PP(16'h169F2,4);
TASK_PP(16'h169F3,4);
TASK_PP(16'h169F4,4);
TASK_PP(16'h169F5,4);
TASK_PP(16'h169F6,4);
TASK_PP(16'h169F7,4);
TASK_PP(16'h169F8,4);
TASK_PP(16'h169F9,4);
TASK_PP(16'h169FA,4);
TASK_PP(16'h169FB,4);
TASK_PP(16'h169FC,4);
TASK_PP(16'h169FD,4);
TASK_PP(16'h169FE,4);
TASK_PP(16'h169FF,4);
TASK_PP(16'h16A00,4);
TASK_PP(16'h16A01,4);
TASK_PP(16'h16A02,4);
TASK_PP(16'h16A03,4);
TASK_PP(16'h16A04,4);
TASK_PP(16'h16A05,4);
TASK_PP(16'h16A06,4);
TASK_PP(16'h16A07,4);
TASK_PP(16'h16A08,4);
TASK_PP(16'h16A09,4);
TASK_PP(16'h16A0A,4);
TASK_PP(16'h16A0B,4);
TASK_PP(16'h16A0C,4);
TASK_PP(16'h16A0D,4);
TASK_PP(16'h16A0E,4);
TASK_PP(16'h16A0F,4);
TASK_PP(16'h16A10,4);
TASK_PP(16'h16A11,4);
TASK_PP(16'h16A12,4);
TASK_PP(16'h16A13,4);
TASK_PP(16'h16A14,4);
TASK_PP(16'h16A15,4);
TASK_PP(16'h16A16,4);
TASK_PP(16'h16A17,4);
TASK_PP(16'h16A18,4);
TASK_PP(16'h16A19,4);
TASK_PP(16'h16A1A,4);
TASK_PP(16'h16A1B,4);
TASK_PP(16'h16A1C,4);
TASK_PP(16'h16A1D,4);
TASK_PP(16'h16A1E,4);
TASK_PP(16'h16A1F,4);
TASK_PP(16'h16A20,4);
TASK_PP(16'h16A21,4);
TASK_PP(16'h16A22,4);
TASK_PP(16'h16A23,4);
TASK_PP(16'h16A24,4);
TASK_PP(16'h16A25,4);
TASK_PP(16'h16A26,4);
TASK_PP(16'h16A27,4);
TASK_PP(16'h16A28,4);
TASK_PP(16'h16A29,4);
TASK_PP(16'h16A2A,4);
TASK_PP(16'h16A2B,4);
TASK_PP(16'h16A2C,4);
TASK_PP(16'h16A2D,4);
TASK_PP(16'h16A2E,4);
TASK_PP(16'h16A2F,4);
TASK_PP(16'h16A30,4);
TASK_PP(16'h16A31,4);
TASK_PP(16'h16A32,4);
TASK_PP(16'h16A33,4);
TASK_PP(16'h16A34,4);
TASK_PP(16'h16A35,4);
TASK_PP(16'h16A36,4);
TASK_PP(16'h16A37,4);
TASK_PP(16'h16A38,4);
TASK_PP(16'h16A39,4);
TASK_PP(16'h16A3A,4);
TASK_PP(16'h16A3B,4);
TASK_PP(16'h16A3C,4);
TASK_PP(16'h16A3D,4);
TASK_PP(16'h16A3E,4);
TASK_PP(16'h16A3F,4);
TASK_PP(16'h16A40,4);
TASK_PP(16'h16A41,4);
TASK_PP(16'h16A42,4);
TASK_PP(16'h16A43,4);
TASK_PP(16'h16A44,4);
TASK_PP(16'h16A45,4);
TASK_PP(16'h16A46,4);
TASK_PP(16'h16A47,4);
TASK_PP(16'h16A48,4);
TASK_PP(16'h16A49,4);
TASK_PP(16'h16A4A,4);
TASK_PP(16'h16A4B,4);
TASK_PP(16'h16A4C,4);
TASK_PP(16'h16A4D,4);
TASK_PP(16'h16A4E,4);
TASK_PP(16'h16A4F,4);
TASK_PP(16'h16A50,4);
TASK_PP(16'h16A51,4);
TASK_PP(16'h16A52,4);
TASK_PP(16'h16A53,4);
TASK_PP(16'h16A54,4);
TASK_PP(16'h16A55,4);
TASK_PP(16'h16A56,4);
TASK_PP(16'h16A57,4);
TASK_PP(16'h16A58,4);
TASK_PP(16'h16A59,4);
TASK_PP(16'h16A5A,4);
TASK_PP(16'h16A5B,4);
TASK_PP(16'h16A5C,4);
TASK_PP(16'h16A5D,4);
TASK_PP(16'h16A5E,4);
TASK_PP(16'h16A5F,4);
TASK_PP(16'h16A60,4);
TASK_PP(16'h16A61,4);
TASK_PP(16'h16A62,4);
TASK_PP(16'h16A63,4);
TASK_PP(16'h16A64,4);
TASK_PP(16'h16A65,4);
TASK_PP(16'h16A66,4);
TASK_PP(16'h16A67,4);
TASK_PP(16'h16A68,4);
TASK_PP(16'h16A69,4);
TASK_PP(16'h16A6A,4);
TASK_PP(16'h16A6B,4);
TASK_PP(16'h16A6C,4);
TASK_PP(16'h16A6D,4);
TASK_PP(16'h16A6E,4);
TASK_PP(16'h16A6F,4);
TASK_PP(16'h16A70,4);
TASK_PP(16'h16A71,4);
TASK_PP(16'h16A72,4);
TASK_PP(16'h16A73,4);
TASK_PP(16'h16A74,4);
TASK_PP(16'h16A75,4);
TASK_PP(16'h16A76,4);
TASK_PP(16'h16A77,4);
TASK_PP(16'h16A78,4);
TASK_PP(16'h16A79,4);
TASK_PP(16'h16A7A,4);
TASK_PP(16'h16A7B,4);
TASK_PP(16'h16A7C,4);
TASK_PP(16'h16A7D,4);
TASK_PP(16'h16A7E,4);
TASK_PP(16'h16A7F,4);
TASK_PP(16'h16A80,4);
TASK_PP(16'h16A81,4);
TASK_PP(16'h16A82,4);
TASK_PP(16'h16A83,4);
TASK_PP(16'h16A84,4);
TASK_PP(16'h16A85,4);
TASK_PP(16'h16A86,4);
TASK_PP(16'h16A87,4);
TASK_PP(16'h16A88,4);
TASK_PP(16'h16A89,4);
TASK_PP(16'h16A8A,4);
TASK_PP(16'h16A8B,4);
TASK_PP(16'h16A8C,4);
TASK_PP(16'h16A8D,4);
TASK_PP(16'h16A8E,4);
TASK_PP(16'h16A8F,4);
TASK_PP(16'h16A90,4);
TASK_PP(16'h16A91,4);
TASK_PP(16'h16A92,4);
TASK_PP(16'h16A93,4);
TASK_PP(16'h16A94,4);
TASK_PP(16'h16A95,4);
TASK_PP(16'h16A96,4);
TASK_PP(16'h16A97,4);
TASK_PP(16'h16A98,4);
TASK_PP(16'h16A99,4);
TASK_PP(16'h16A9A,4);
TASK_PP(16'h16A9B,4);
TASK_PP(16'h16A9C,4);
TASK_PP(16'h16A9D,4);
TASK_PP(16'h16A9E,4);
TASK_PP(16'h16A9F,4);
TASK_PP(16'h16AA0,4);
TASK_PP(16'h16AA1,4);
TASK_PP(16'h16AA2,4);
TASK_PP(16'h16AA3,4);
TASK_PP(16'h16AA4,4);
TASK_PP(16'h16AA5,4);
TASK_PP(16'h16AA6,4);
TASK_PP(16'h16AA7,4);
TASK_PP(16'h16AA8,4);
TASK_PP(16'h16AA9,4);
TASK_PP(16'h16AAA,4);
TASK_PP(16'h16AAB,4);
TASK_PP(16'h16AAC,4);
TASK_PP(16'h16AAD,4);
TASK_PP(16'h16AAE,4);
TASK_PP(16'h16AAF,4);
TASK_PP(16'h16AB0,4);
TASK_PP(16'h16AB1,4);
TASK_PP(16'h16AB2,4);
TASK_PP(16'h16AB3,4);
TASK_PP(16'h16AB4,4);
TASK_PP(16'h16AB5,4);
TASK_PP(16'h16AB6,4);
TASK_PP(16'h16AB7,4);
TASK_PP(16'h16AB8,4);
TASK_PP(16'h16AB9,4);
TASK_PP(16'h16ABA,4);
TASK_PP(16'h16ABB,4);
TASK_PP(16'h16ABC,4);
TASK_PP(16'h16ABD,4);
TASK_PP(16'h16ABE,4);
TASK_PP(16'h16ABF,4);
TASK_PP(16'h16AC0,4);
TASK_PP(16'h16AC1,4);
TASK_PP(16'h16AC2,4);
TASK_PP(16'h16AC3,4);
TASK_PP(16'h16AC4,4);
TASK_PP(16'h16AC5,4);
TASK_PP(16'h16AC6,4);
TASK_PP(16'h16AC7,4);
TASK_PP(16'h16AC8,4);
TASK_PP(16'h16AC9,4);
TASK_PP(16'h16ACA,4);
TASK_PP(16'h16ACB,4);
TASK_PP(16'h16ACC,4);
TASK_PP(16'h16ACD,4);
TASK_PP(16'h16ACE,4);
TASK_PP(16'h16ACF,4);
TASK_PP(16'h16AD0,4);
TASK_PP(16'h16AD1,4);
TASK_PP(16'h16AD2,4);
TASK_PP(16'h16AD3,4);
TASK_PP(16'h16AD4,4);
TASK_PP(16'h16AD5,4);
TASK_PP(16'h16AD6,4);
TASK_PP(16'h16AD7,4);
TASK_PP(16'h16AD8,4);
TASK_PP(16'h16AD9,4);
TASK_PP(16'h16ADA,4);
TASK_PP(16'h16ADB,4);
TASK_PP(16'h16ADC,4);
TASK_PP(16'h16ADD,4);
TASK_PP(16'h16ADE,4);
TASK_PP(16'h16ADF,4);
TASK_PP(16'h16AE0,4);
TASK_PP(16'h16AE1,4);
TASK_PP(16'h16AE2,4);
TASK_PP(16'h16AE3,4);
TASK_PP(16'h16AE4,4);
TASK_PP(16'h16AE5,4);
TASK_PP(16'h16AE6,4);
TASK_PP(16'h16AE7,4);
TASK_PP(16'h16AE8,4);
TASK_PP(16'h16AE9,4);
TASK_PP(16'h16AEA,4);
TASK_PP(16'h16AEB,4);
TASK_PP(16'h16AEC,4);
TASK_PP(16'h16AED,4);
TASK_PP(16'h16AEE,4);
TASK_PP(16'h16AEF,4);
TASK_PP(16'h16AF0,4);
TASK_PP(16'h16AF1,4);
TASK_PP(16'h16AF2,4);
TASK_PP(16'h16AF3,4);
TASK_PP(16'h16AF4,4);
TASK_PP(16'h16AF5,4);
TASK_PP(16'h16AF6,4);
TASK_PP(16'h16AF7,4);
TASK_PP(16'h16AF8,4);
TASK_PP(16'h16AF9,4);
TASK_PP(16'h16AFA,4);
TASK_PP(16'h16AFB,4);
TASK_PP(16'h16AFC,4);
TASK_PP(16'h16AFD,4);
TASK_PP(16'h16AFE,4);
TASK_PP(16'h16AFF,4);
TASK_PP(16'h16B00,4);
TASK_PP(16'h16B01,4);
TASK_PP(16'h16B02,4);
TASK_PP(16'h16B03,4);
TASK_PP(16'h16B04,4);
TASK_PP(16'h16B05,4);
TASK_PP(16'h16B06,4);
TASK_PP(16'h16B07,4);
TASK_PP(16'h16B08,4);
TASK_PP(16'h16B09,4);
TASK_PP(16'h16B0A,4);
TASK_PP(16'h16B0B,4);
TASK_PP(16'h16B0C,4);
TASK_PP(16'h16B0D,4);
TASK_PP(16'h16B0E,4);
TASK_PP(16'h16B0F,4);
TASK_PP(16'h16B10,4);
TASK_PP(16'h16B11,4);
TASK_PP(16'h16B12,4);
TASK_PP(16'h16B13,4);
TASK_PP(16'h16B14,4);
TASK_PP(16'h16B15,4);
TASK_PP(16'h16B16,4);
TASK_PP(16'h16B17,4);
TASK_PP(16'h16B18,4);
TASK_PP(16'h16B19,4);
TASK_PP(16'h16B1A,4);
TASK_PP(16'h16B1B,4);
TASK_PP(16'h16B1C,4);
TASK_PP(16'h16B1D,4);
TASK_PP(16'h16B1E,4);
TASK_PP(16'h16B1F,4);
TASK_PP(16'h16B20,4);
TASK_PP(16'h16B21,4);
TASK_PP(16'h16B22,4);
TASK_PP(16'h16B23,4);
TASK_PP(16'h16B24,4);
TASK_PP(16'h16B25,4);
TASK_PP(16'h16B26,4);
TASK_PP(16'h16B27,4);
TASK_PP(16'h16B28,4);
TASK_PP(16'h16B29,4);
TASK_PP(16'h16B2A,4);
TASK_PP(16'h16B2B,4);
TASK_PP(16'h16B2C,4);
TASK_PP(16'h16B2D,4);
TASK_PP(16'h16B2E,4);
TASK_PP(16'h16B2F,4);
TASK_PP(16'h16B30,4);
TASK_PP(16'h16B31,4);
TASK_PP(16'h16B32,4);
TASK_PP(16'h16B33,4);
TASK_PP(16'h16B34,4);
TASK_PP(16'h16B35,4);
TASK_PP(16'h16B36,4);
TASK_PP(16'h16B37,4);
TASK_PP(16'h16B38,4);
TASK_PP(16'h16B39,4);
TASK_PP(16'h16B3A,4);
TASK_PP(16'h16B3B,4);
TASK_PP(16'h16B3C,4);
TASK_PP(16'h16B3D,4);
TASK_PP(16'h16B3E,4);
TASK_PP(16'h16B3F,4);
TASK_PP(16'h16B40,4);
TASK_PP(16'h16B41,4);
TASK_PP(16'h16B42,4);
TASK_PP(16'h16B43,4);
TASK_PP(16'h16B44,4);
TASK_PP(16'h16B45,4);
TASK_PP(16'h16B46,4);
TASK_PP(16'h16B47,4);
TASK_PP(16'h16B48,4);
TASK_PP(16'h16B49,4);
TASK_PP(16'h16B4A,4);
TASK_PP(16'h16B4B,4);
TASK_PP(16'h16B4C,4);
TASK_PP(16'h16B4D,4);
TASK_PP(16'h16B4E,4);
TASK_PP(16'h16B4F,4);
TASK_PP(16'h16B50,4);
TASK_PP(16'h16B51,4);
TASK_PP(16'h16B52,4);
TASK_PP(16'h16B53,4);
TASK_PP(16'h16B54,4);
TASK_PP(16'h16B55,4);
TASK_PP(16'h16B56,4);
TASK_PP(16'h16B57,4);
TASK_PP(16'h16B58,4);
TASK_PP(16'h16B59,4);
TASK_PP(16'h16B5A,4);
TASK_PP(16'h16B5B,4);
TASK_PP(16'h16B5C,4);
TASK_PP(16'h16B5D,4);
TASK_PP(16'h16B5E,4);
TASK_PP(16'h16B5F,4);
TASK_PP(16'h16B60,4);
TASK_PP(16'h16B61,4);
TASK_PP(16'h16B62,4);
TASK_PP(16'h16B63,4);
TASK_PP(16'h16B64,4);
TASK_PP(16'h16B65,4);
TASK_PP(16'h16B66,4);
TASK_PP(16'h16B67,4);
TASK_PP(16'h16B68,4);
TASK_PP(16'h16B69,4);
TASK_PP(16'h16B6A,4);
TASK_PP(16'h16B6B,4);
TASK_PP(16'h16B6C,4);
TASK_PP(16'h16B6D,4);
TASK_PP(16'h16B6E,4);
TASK_PP(16'h16B6F,4);
TASK_PP(16'h16B70,4);
TASK_PP(16'h16B71,4);
TASK_PP(16'h16B72,4);
TASK_PP(16'h16B73,4);
TASK_PP(16'h16B74,4);
TASK_PP(16'h16B75,4);
TASK_PP(16'h16B76,4);
TASK_PP(16'h16B77,4);
TASK_PP(16'h16B78,4);
TASK_PP(16'h16B79,4);
TASK_PP(16'h16B7A,4);
TASK_PP(16'h16B7B,4);
TASK_PP(16'h16B7C,4);
TASK_PP(16'h16B7D,4);
TASK_PP(16'h16B7E,4);
TASK_PP(16'h16B7F,4);
TASK_PP(16'h16B80,4);
TASK_PP(16'h16B81,4);
TASK_PP(16'h16B82,4);
TASK_PP(16'h16B83,4);
TASK_PP(16'h16B84,4);
TASK_PP(16'h16B85,4);
TASK_PP(16'h16B86,4);
TASK_PP(16'h16B87,4);
TASK_PP(16'h16B88,4);
TASK_PP(16'h16B89,4);
TASK_PP(16'h16B8A,4);
TASK_PP(16'h16B8B,4);
TASK_PP(16'h16B8C,4);
TASK_PP(16'h16B8D,4);
TASK_PP(16'h16B8E,4);
TASK_PP(16'h16B8F,4);
TASK_PP(16'h16B90,4);
TASK_PP(16'h16B91,4);
TASK_PP(16'h16B92,4);
TASK_PP(16'h16B93,4);
TASK_PP(16'h16B94,4);
TASK_PP(16'h16B95,4);
TASK_PP(16'h16B96,4);
TASK_PP(16'h16B97,4);
TASK_PP(16'h16B98,4);
TASK_PP(16'h16B99,4);
TASK_PP(16'h16B9A,4);
TASK_PP(16'h16B9B,4);
TASK_PP(16'h16B9C,4);
TASK_PP(16'h16B9D,4);
TASK_PP(16'h16B9E,4);
TASK_PP(16'h16B9F,4);
TASK_PP(16'h16BA0,4);
TASK_PP(16'h16BA1,4);
TASK_PP(16'h16BA2,4);
TASK_PP(16'h16BA3,4);
TASK_PP(16'h16BA4,4);
TASK_PP(16'h16BA5,4);
TASK_PP(16'h16BA6,4);
TASK_PP(16'h16BA7,4);
TASK_PP(16'h16BA8,4);
TASK_PP(16'h16BA9,4);
TASK_PP(16'h16BAA,4);
TASK_PP(16'h16BAB,4);
TASK_PP(16'h16BAC,4);
TASK_PP(16'h16BAD,4);
TASK_PP(16'h16BAE,4);
TASK_PP(16'h16BAF,4);
TASK_PP(16'h16BB0,4);
TASK_PP(16'h16BB1,4);
TASK_PP(16'h16BB2,4);
TASK_PP(16'h16BB3,4);
TASK_PP(16'h16BB4,4);
TASK_PP(16'h16BB5,4);
TASK_PP(16'h16BB6,4);
TASK_PP(16'h16BB7,4);
TASK_PP(16'h16BB8,4);
TASK_PP(16'h16BB9,4);
TASK_PP(16'h16BBA,4);
TASK_PP(16'h16BBB,4);
TASK_PP(16'h16BBC,4);
TASK_PP(16'h16BBD,4);
TASK_PP(16'h16BBE,4);
TASK_PP(16'h16BBF,4);
TASK_PP(16'h16BC0,4);
TASK_PP(16'h16BC1,4);
TASK_PP(16'h16BC2,4);
TASK_PP(16'h16BC3,4);
TASK_PP(16'h16BC4,4);
TASK_PP(16'h16BC5,4);
TASK_PP(16'h16BC6,4);
TASK_PP(16'h16BC7,4);
TASK_PP(16'h16BC8,4);
TASK_PP(16'h16BC9,4);
TASK_PP(16'h16BCA,4);
TASK_PP(16'h16BCB,4);
TASK_PP(16'h16BCC,4);
TASK_PP(16'h16BCD,4);
TASK_PP(16'h16BCE,4);
TASK_PP(16'h16BCF,4);
TASK_PP(16'h16BD0,4);
TASK_PP(16'h16BD1,4);
TASK_PP(16'h16BD2,4);
TASK_PP(16'h16BD3,4);
TASK_PP(16'h16BD4,4);
TASK_PP(16'h16BD5,4);
TASK_PP(16'h16BD6,4);
TASK_PP(16'h16BD7,4);
TASK_PP(16'h16BD8,4);
TASK_PP(16'h16BD9,4);
TASK_PP(16'h16BDA,4);
TASK_PP(16'h16BDB,4);
TASK_PP(16'h16BDC,4);
TASK_PP(16'h16BDD,4);
TASK_PP(16'h16BDE,4);
TASK_PP(16'h16BDF,4);
TASK_PP(16'h16BE0,4);
TASK_PP(16'h16BE1,4);
TASK_PP(16'h16BE2,4);
TASK_PP(16'h16BE3,4);
TASK_PP(16'h16BE4,4);
TASK_PP(16'h16BE5,4);
TASK_PP(16'h16BE6,4);
TASK_PP(16'h16BE7,4);
TASK_PP(16'h16BE8,4);
TASK_PP(16'h16BE9,4);
TASK_PP(16'h16BEA,4);
TASK_PP(16'h16BEB,4);
TASK_PP(16'h16BEC,4);
TASK_PP(16'h16BED,4);
TASK_PP(16'h16BEE,4);
TASK_PP(16'h16BEF,4);
TASK_PP(16'h16BF0,4);
TASK_PP(16'h16BF1,4);
TASK_PP(16'h16BF2,4);
TASK_PP(16'h16BF3,4);
TASK_PP(16'h16BF4,4);
TASK_PP(16'h16BF5,4);
TASK_PP(16'h16BF6,4);
TASK_PP(16'h16BF7,4);
TASK_PP(16'h16BF8,4);
TASK_PP(16'h16BF9,4);
TASK_PP(16'h16BFA,4);
TASK_PP(16'h16BFB,4);
TASK_PP(16'h16BFC,4);
TASK_PP(16'h16BFD,4);
TASK_PP(16'h16BFE,4);
TASK_PP(16'h16BFF,4);
TASK_PP(16'h16C00,4);
TASK_PP(16'h16C01,4);
TASK_PP(16'h16C02,4);
TASK_PP(16'h16C03,4);
TASK_PP(16'h16C04,4);
TASK_PP(16'h16C05,4);
TASK_PP(16'h16C06,4);
TASK_PP(16'h16C07,4);
TASK_PP(16'h16C08,4);
TASK_PP(16'h16C09,4);
TASK_PP(16'h16C0A,4);
TASK_PP(16'h16C0B,4);
TASK_PP(16'h16C0C,4);
TASK_PP(16'h16C0D,4);
TASK_PP(16'h16C0E,4);
TASK_PP(16'h16C0F,4);
TASK_PP(16'h16C10,4);
TASK_PP(16'h16C11,4);
TASK_PP(16'h16C12,4);
TASK_PP(16'h16C13,4);
TASK_PP(16'h16C14,4);
TASK_PP(16'h16C15,4);
TASK_PP(16'h16C16,4);
TASK_PP(16'h16C17,4);
TASK_PP(16'h16C18,4);
TASK_PP(16'h16C19,4);
TASK_PP(16'h16C1A,4);
TASK_PP(16'h16C1B,4);
TASK_PP(16'h16C1C,4);
TASK_PP(16'h16C1D,4);
TASK_PP(16'h16C1E,4);
TASK_PP(16'h16C1F,4);
TASK_PP(16'h16C20,4);
TASK_PP(16'h16C21,4);
TASK_PP(16'h16C22,4);
TASK_PP(16'h16C23,4);
TASK_PP(16'h16C24,4);
TASK_PP(16'h16C25,4);
TASK_PP(16'h16C26,4);
TASK_PP(16'h16C27,4);
TASK_PP(16'h16C28,4);
TASK_PP(16'h16C29,4);
TASK_PP(16'h16C2A,4);
TASK_PP(16'h16C2B,4);
TASK_PP(16'h16C2C,4);
TASK_PP(16'h16C2D,4);
TASK_PP(16'h16C2E,4);
TASK_PP(16'h16C2F,4);
TASK_PP(16'h16C30,4);
TASK_PP(16'h16C31,4);
TASK_PP(16'h16C32,4);
TASK_PP(16'h16C33,4);
TASK_PP(16'h16C34,4);
TASK_PP(16'h16C35,4);
TASK_PP(16'h16C36,4);
TASK_PP(16'h16C37,4);
TASK_PP(16'h16C38,4);
TASK_PP(16'h16C39,4);
TASK_PP(16'h16C3A,4);
TASK_PP(16'h16C3B,4);
TASK_PP(16'h16C3C,4);
TASK_PP(16'h16C3D,4);
TASK_PP(16'h16C3E,4);
TASK_PP(16'h16C3F,4);
TASK_PP(16'h16C40,4);
TASK_PP(16'h16C41,4);
TASK_PP(16'h16C42,4);
TASK_PP(16'h16C43,4);
TASK_PP(16'h16C44,4);
TASK_PP(16'h16C45,4);
TASK_PP(16'h16C46,4);
TASK_PP(16'h16C47,4);
TASK_PP(16'h16C48,4);
TASK_PP(16'h16C49,4);
TASK_PP(16'h16C4A,4);
TASK_PP(16'h16C4B,4);
TASK_PP(16'h16C4C,4);
TASK_PP(16'h16C4D,4);
TASK_PP(16'h16C4E,4);
TASK_PP(16'h16C4F,4);
TASK_PP(16'h16C50,4);
TASK_PP(16'h16C51,4);
TASK_PP(16'h16C52,4);
TASK_PP(16'h16C53,4);
TASK_PP(16'h16C54,4);
TASK_PP(16'h16C55,4);
TASK_PP(16'h16C56,4);
TASK_PP(16'h16C57,4);
TASK_PP(16'h16C58,4);
TASK_PP(16'h16C59,4);
TASK_PP(16'h16C5A,4);
TASK_PP(16'h16C5B,4);
TASK_PP(16'h16C5C,4);
TASK_PP(16'h16C5D,4);
TASK_PP(16'h16C5E,4);
TASK_PP(16'h16C5F,4);
TASK_PP(16'h16C60,4);
TASK_PP(16'h16C61,4);
TASK_PP(16'h16C62,4);
TASK_PP(16'h16C63,4);
TASK_PP(16'h16C64,4);
TASK_PP(16'h16C65,4);
TASK_PP(16'h16C66,4);
TASK_PP(16'h16C67,4);
TASK_PP(16'h16C68,4);
TASK_PP(16'h16C69,4);
TASK_PP(16'h16C6A,4);
TASK_PP(16'h16C6B,4);
TASK_PP(16'h16C6C,4);
TASK_PP(16'h16C6D,4);
TASK_PP(16'h16C6E,4);
TASK_PP(16'h16C6F,4);
TASK_PP(16'h16C70,4);
TASK_PP(16'h16C71,4);
TASK_PP(16'h16C72,4);
TASK_PP(16'h16C73,4);
TASK_PP(16'h16C74,4);
TASK_PP(16'h16C75,4);
TASK_PP(16'h16C76,4);
TASK_PP(16'h16C77,4);
TASK_PP(16'h16C78,4);
TASK_PP(16'h16C79,4);
TASK_PP(16'h16C7A,4);
TASK_PP(16'h16C7B,4);
TASK_PP(16'h16C7C,4);
TASK_PP(16'h16C7D,4);
TASK_PP(16'h16C7E,4);
TASK_PP(16'h16C7F,4);
TASK_PP(16'h16C80,4);
TASK_PP(16'h16C81,4);
TASK_PP(16'h16C82,4);
TASK_PP(16'h16C83,4);
TASK_PP(16'h16C84,4);
TASK_PP(16'h16C85,4);
TASK_PP(16'h16C86,4);
TASK_PP(16'h16C87,4);
TASK_PP(16'h16C88,4);
TASK_PP(16'h16C89,4);
TASK_PP(16'h16C8A,4);
TASK_PP(16'h16C8B,4);
TASK_PP(16'h16C8C,4);
TASK_PP(16'h16C8D,4);
TASK_PP(16'h16C8E,4);
TASK_PP(16'h16C8F,4);
TASK_PP(16'h16C90,4);
TASK_PP(16'h16C91,4);
TASK_PP(16'h16C92,4);
TASK_PP(16'h16C93,4);
TASK_PP(16'h16C94,4);
TASK_PP(16'h16C95,4);
TASK_PP(16'h16C96,4);
TASK_PP(16'h16C97,4);
TASK_PP(16'h16C98,4);
TASK_PP(16'h16C99,4);
TASK_PP(16'h16C9A,4);
TASK_PP(16'h16C9B,4);
TASK_PP(16'h16C9C,4);
TASK_PP(16'h16C9D,4);
TASK_PP(16'h16C9E,4);
TASK_PP(16'h16C9F,4);
TASK_PP(16'h16CA0,4);
TASK_PP(16'h16CA1,4);
TASK_PP(16'h16CA2,4);
TASK_PP(16'h16CA3,4);
TASK_PP(16'h16CA4,4);
TASK_PP(16'h16CA5,4);
TASK_PP(16'h16CA6,4);
TASK_PP(16'h16CA7,4);
TASK_PP(16'h16CA8,4);
TASK_PP(16'h16CA9,4);
TASK_PP(16'h16CAA,4);
TASK_PP(16'h16CAB,4);
TASK_PP(16'h16CAC,4);
TASK_PP(16'h16CAD,4);
TASK_PP(16'h16CAE,4);
TASK_PP(16'h16CAF,4);
TASK_PP(16'h16CB0,4);
TASK_PP(16'h16CB1,4);
TASK_PP(16'h16CB2,4);
TASK_PP(16'h16CB3,4);
TASK_PP(16'h16CB4,4);
TASK_PP(16'h16CB5,4);
TASK_PP(16'h16CB6,4);
TASK_PP(16'h16CB7,4);
TASK_PP(16'h16CB8,4);
TASK_PP(16'h16CB9,4);
TASK_PP(16'h16CBA,4);
TASK_PP(16'h16CBB,4);
TASK_PP(16'h16CBC,4);
TASK_PP(16'h16CBD,4);
TASK_PP(16'h16CBE,4);
TASK_PP(16'h16CBF,4);
TASK_PP(16'h16CC0,4);
TASK_PP(16'h16CC1,4);
TASK_PP(16'h16CC2,4);
TASK_PP(16'h16CC3,4);
TASK_PP(16'h16CC4,4);
TASK_PP(16'h16CC5,4);
TASK_PP(16'h16CC6,4);
TASK_PP(16'h16CC7,4);
TASK_PP(16'h16CC8,4);
TASK_PP(16'h16CC9,4);
TASK_PP(16'h16CCA,4);
TASK_PP(16'h16CCB,4);
TASK_PP(16'h16CCC,4);
TASK_PP(16'h16CCD,4);
TASK_PP(16'h16CCE,4);
TASK_PP(16'h16CCF,4);
TASK_PP(16'h16CD0,4);
TASK_PP(16'h16CD1,4);
TASK_PP(16'h16CD2,4);
TASK_PP(16'h16CD3,4);
TASK_PP(16'h16CD4,4);
TASK_PP(16'h16CD5,4);
TASK_PP(16'h16CD6,4);
TASK_PP(16'h16CD7,4);
TASK_PP(16'h16CD8,4);
TASK_PP(16'h16CD9,4);
TASK_PP(16'h16CDA,4);
TASK_PP(16'h16CDB,4);
TASK_PP(16'h16CDC,4);
TASK_PP(16'h16CDD,4);
TASK_PP(16'h16CDE,4);
TASK_PP(16'h16CDF,4);
TASK_PP(16'h16CE0,4);
TASK_PP(16'h16CE1,4);
TASK_PP(16'h16CE2,4);
TASK_PP(16'h16CE3,4);
TASK_PP(16'h16CE4,4);
TASK_PP(16'h16CE5,4);
TASK_PP(16'h16CE6,4);
TASK_PP(16'h16CE7,4);
TASK_PP(16'h16CE8,4);
TASK_PP(16'h16CE9,4);
TASK_PP(16'h16CEA,4);
TASK_PP(16'h16CEB,4);
TASK_PP(16'h16CEC,4);
TASK_PP(16'h16CED,4);
TASK_PP(16'h16CEE,4);
TASK_PP(16'h16CEF,4);
TASK_PP(16'h16CF0,4);
TASK_PP(16'h16CF1,4);
TASK_PP(16'h16CF2,4);
TASK_PP(16'h16CF3,4);
TASK_PP(16'h16CF4,4);
TASK_PP(16'h16CF5,4);
TASK_PP(16'h16CF6,4);
TASK_PP(16'h16CF7,4);
TASK_PP(16'h16CF8,4);
TASK_PP(16'h16CF9,4);
TASK_PP(16'h16CFA,4);
TASK_PP(16'h16CFB,4);
TASK_PP(16'h16CFC,4);
TASK_PP(16'h16CFD,4);
TASK_PP(16'h16CFE,4);
TASK_PP(16'h16CFF,4);
TASK_PP(16'h16D00,4);
TASK_PP(16'h16D01,4);
TASK_PP(16'h16D02,4);
TASK_PP(16'h16D03,4);
TASK_PP(16'h16D04,4);
TASK_PP(16'h16D05,4);
TASK_PP(16'h16D06,4);
TASK_PP(16'h16D07,4);
TASK_PP(16'h16D08,4);
TASK_PP(16'h16D09,4);
TASK_PP(16'h16D0A,4);
TASK_PP(16'h16D0B,4);
TASK_PP(16'h16D0C,4);
TASK_PP(16'h16D0D,4);
TASK_PP(16'h16D0E,4);
TASK_PP(16'h16D0F,4);
TASK_PP(16'h16D10,4);
TASK_PP(16'h16D11,4);
TASK_PP(16'h16D12,4);
TASK_PP(16'h16D13,4);
TASK_PP(16'h16D14,4);
TASK_PP(16'h16D15,4);
TASK_PP(16'h16D16,4);
TASK_PP(16'h16D17,4);
TASK_PP(16'h16D18,4);
TASK_PP(16'h16D19,4);
TASK_PP(16'h16D1A,4);
TASK_PP(16'h16D1B,4);
TASK_PP(16'h16D1C,4);
TASK_PP(16'h16D1D,4);
TASK_PP(16'h16D1E,4);
TASK_PP(16'h16D1F,4);
TASK_PP(16'h16D20,4);
TASK_PP(16'h16D21,4);
TASK_PP(16'h16D22,4);
TASK_PP(16'h16D23,4);
TASK_PP(16'h16D24,4);
TASK_PP(16'h16D25,4);
TASK_PP(16'h16D26,4);
TASK_PP(16'h16D27,4);
TASK_PP(16'h16D28,4);
TASK_PP(16'h16D29,4);
TASK_PP(16'h16D2A,4);
TASK_PP(16'h16D2B,4);
TASK_PP(16'h16D2C,4);
TASK_PP(16'h16D2D,4);
TASK_PP(16'h16D2E,4);
TASK_PP(16'h16D2F,4);
TASK_PP(16'h16D30,4);
TASK_PP(16'h16D31,4);
TASK_PP(16'h16D32,4);
TASK_PP(16'h16D33,4);
TASK_PP(16'h16D34,4);
TASK_PP(16'h16D35,4);
TASK_PP(16'h16D36,4);
TASK_PP(16'h16D37,4);
TASK_PP(16'h16D38,4);
TASK_PP(16'h16D39,4);
TASK_PP(16'h16D3A,4);
TASK_PP(16'h16D3B,4);
TASK_PP(16'h16D3C,4);
TASK_PP(16'h16D3D,4);
TASK_PP(16'h16D3E,4);
TASK_PP(16'h16D3F,4);
TASK_PP(16'h16D40,4);
TASK_PP(16'h16D41,4);
TASK_PP(16'h16D42,4);
TASK_PP(16'h16D43,4);
TASK_PP(16'h16D44,4);
TASK_PP(16'h16D45,4);
TASK_PP(16'h16D46,4);
TASK_PP(16'h16D47,4);
TASK_PP(16'h16D48,4);
TASK_PP(16'h16D49,4);
TASK_PP(16'h16D4A,4);
TASK_PP(16'h16D4B,4);
TASK_PP(16'h16D4C,4);
TASK_PP(16'h16D4D,4);
TASK_PP(16'h16D4E,4);
TASK_PP(16'h16D4F,4);
TASK_PP(16'h16D50,4);
TASK_PP(16'h16D51,4);
TASK_PP(16'h16D52,4);
TASK_PP(16'h16D53,4);
TASK_PP(16'h16D54,4);
TASK_PP(16'h16D55,4);
TASK_PP(16'h16D56,4);
TASK_PP(16'h16D57,4);
TASK_PP(16'h16D58,4);
TASK_PP(16'h16D59,4);
TASK_PP(16'h16D5A,4);
TASK_PP(16'h16D5B,4);
TASK_PP(16'h16D5C,4);
TASK_PP(16'h16D5D,4);
TASK_PP(16'h16D5E,4);
TASK_PP(16'h16D5F,4);
TASK_PP(16'h16D60,4);
TASK_PP(16'h16D61,4);
TASK_PP(16'h16D62,4);
TASK_PP(16'h16D63,4);
TASK_PP(16'h16D64,4);
TASK_PP(16'h16D65,4);
TASK_PP(16'h16D66,4);
TASK_PP(16'h16D67,4);
TASK_PP(16'h16D68,4);
TASK_PP(16'h16D69,4);
TASK_PP(16'h16D6A,4);
TASK_PP(16'h16D6B,4);
TASK_PP(16'h16D6C,4);
TASK_PP(16'h16D6D,4);
TASK_PP(16'h16D6E,4);
TASK_PP(16'h16D6F,4);
TASK_PP(16'h16D70,4);
TASK_PP(16'h16D71,4);
TASK_PP(16'h16D72,4);
TASK_PP(16'h16D73,4);
TASK_PP(16'h16D74,4);
TASK_PP(16'h16D75,4);
TASK_PP(16'h16D76,4);
TASK_PP(16'h16D77,4);
TASK_PP(16'h16D78,4);
TASK_PP(16'h16D79,4);
TASK_PP(16'h16D7A,4);
TASK_PP(16'h16D7B,4);
TASK_PP(16'h16D7C,4);
TASK_PP(16'h16D7D,4);
TASK_PP(16'h16D7E,4);
TASK_PP(16'h16D7F,4);
TASK_PP(16'h16D80,4);
TASK_PP(16'h16D81,4);
TASK_PP(16'h16D82,4);
TASK_PP(16'h16D83,4);
TASK_PP(16'h16D84,4);
TASK_PP(16'h16D85,4);
TASK_PP(16'h16D86,4);
TASK_PP(16'h16D87,4);
TASK_PP(16'h16D88,4);
TASK_PP(16'h16D89,4);
TASK_PP(16'h16D8A,4);
TASK_PP(16'h16D8B,4);
TASK_PP(16'h16D8C,4);
TASK_PP(16'h16D8D,4);
TASK_PP(16'h16D8E,4);
TASK_PP(16'h16D8F,4);
TASK_PP(16'h16D90,4);
TASK_PP(16'h16D91,4);
TASK_PP(16'h16D92,4);
TASK_PP(16'h16D93,4);
TASK_PP(16'h16D94,4);
TASK_PP(16'h16D95,4);
TASK_PP(16'h16D96,4);
TASK_PP(16'h16D97,4);
TASK_PP(16'h16D98,4);
TASK_PP(16'h16D99,4);
TASK_PP(16'h16D9A,4);
TASK_PP(16'h16D9B,4);
TASK_PP(16'h16D9C,4);
TASK_PP(16'h16D9D,4);
TASK_PP(16'h16D9E,4);
TASK_PP(16'h16D9F,4);
TASK_PP(16'h16DA0,4);
TASK_PP(16'h16DA1,4);
TASK_PP(16'h16DA2,4);
TASK_PP(16'h16DA3,4);
TASK_PP(16'h16DA4,4);
TASK_PP(16'h16DA5,4);
TASK_PP(16'h16DA6,4);
TASK_PP(16'h16DA7,4);
TASK_PP(16'h16DA8,4);
TASK_PP(16'h16DA9,4);
TASK_PP(16'h16DAA,4);
TASK_PP(16'h16DAB,4);
TASK_PP(16'h16DAC,4);
TASK_PP(16'h16DAD,4);
TASK_PP(16'h16DAE,4);
TASK_PP(16'h16DAF,4);
TASK_PP(16'h16DB0,4);
TASK_PP(16'h16DB1,4);
TASK_PP(16'h16DB2,4);
TASK_PP(16'h16DB3,4);
TASK_PP(16'h16DB4,4);
TASK_PP(16'h16DB5,4);
TASK_PP(16'h16DB6,4);
TASK_PP(16'h16DB7,4);
TASK_PP(16'h16DB8,4);
TASK_PP(16'h16DB9,4);
TASK_PP(16'h16DBA,4);
TASK_PP(16'h16DBB,4);
TASK_PP(16'h16DBC,4);
TASK_PP(16'h16DBD,4);
TASK_PP(16'h16DBE,4);
TASK_PP(16'h16DBF,4);
TASK_PP(16'h16DC0,4);
TASK_PP(16'h16DC1,4);
TASK_PP(16'h16DC2,4);
TASK_PP(16'h16DC3,4);
TASK_PP(16'h16DC4,4);
TASK_PP(16'h16DC5,4);
TASK_PP(16'h16DC6,4);
TASK_PP(16'h16DC7,4);
TASK_PP(16'h16DC8,4);
TASK_PP(16'h16DC9,4);
TASK_PP(16'h16DCA,4);
TASK_PP(16'h16DCB,4);
TASK_PP(16'h16DCC,4);
TASK_PP(16'h16DCD,4);
TASK_PP(16'h16DCE,4);
TASK_PP(16'h16DCF,4);
TASK_PP(16'h16DD0,4);
TASK_PP(16'h16DD1,4);
TASK_PP(16'h16DD2,4);
TASK_PP(16'h16DD3,4);
TASK_PP(16'h16DD4,4);
TASK_PP(16'h16DD5,4);
TASK_PP(16'h16DD6,4);
TASK_PP(16'h16DD7,4);
TASK_PP(16'h16DD8,4);
TASK_PP(16'h16DD9,4);
TASK_PP(16'h16DDA,4);
TASK_PP(16'h16DDB,4);
TASK_PP(16'h16DDC,4);
TASK_PP(16'h16DDD,4);
TASK_PP(16'h16DDE,4);
TASK_PP(16'h16DDF,4);
TASK_PP(16'h16DE0,4);
TASK_PP(16'h16DE1,4);
TASK_PP(16'h16DE2,4);
TASK_PP(16'h16DE3,4);
TASK_PP(16'h16DE4,4);
TASK_PP(16'h16DE5,4);
TASK_PP(16'h16DE6,4);
TASK_PP(16'h16DE7,4);
TASK_PP(16'h16DE8,4);
TASK_PP(16'h16DE9,4);
TASK_PP(16'h16DEA,4);
TASK_PP(16'h16DEB,4);
TASK_PP(16'h16DEC,4);
TASK_PP(16'h16DED,4);
TASK_PP(16'h16DEE,4);
TASK_PP(16'h16DEF,4);
TASK_PP(16'h16DF0,4);
TASK_PP(16'h16DF1,4);
TASK_PP(16'h16DF2,4);
TASK_PP(16'h16DF3,4);
TASK_PP(16'h16DF4,4);
TASK_PP(16'h16DF5,4);
TASK_PP(16'h16DF6,4);
TASK_PP(16'h16DF7,4);
TASK_PP(16'h16DF8,4);
TASK_PP(16'h16DF9,4);
TASK_PP(16'h16DFA,4);
TASK_PP(16'h16DFB,4);
TASK_PP(16'h16DFC,4);
TASK_PP(16'h16DFD,4);
TASK_PP(16'h16DFE,4);
TASK_PP(16'h16DFF,4);
TASK_PP(16'h16E00,4);
TASK_PP(16'h16E01,4);
TASK_PP(16'h16E02,4);
TASK_PP(16'h16E03,4);
TASK_PP(16'h16E04,4);
TASK_PP(16'h16E05,4);
TASK_PP(16'h16E06,4);
TASK_PP(16'h16E07,4);
TASK_PP(16'h16E08,4);
TASK_PP(16'h16E09,4);
TASK_PP(16'h16E0A,4);
TASK_PP(16'h16E0B,4);
TASK_PP(16'h16E0C,4);
TASK_PP(16'h16E0D,4);
TASK_PP(16'h16E0E,4);
TASK_PP(16'h16E0F,4);
TASK_PP(16'h16E10,4);
TASK_PP(16'h16E11,4);
TASK_PP(16'h16E12,4);
TASK_PP(16'h16E13,4);
TASK_PP(16'h16E14,4);
TASK_PP(16'h16E15,4);
TASK_PP(16'h16E16,4);
TASK_PP(16'h16E17,4);
TASK_PP(16'h16E18,4);
TASK_PP(16'h16E19,4);
TASK_PP(16'h16E1A,4);
TASK_PP(16'h16E1B,4);
TASK_PP(16'h16E1C,4);
TASK_PP(16'h16E1D,4);
TASK_PP(16'h16E1E,4);
TASK_PP(16'h16E1F,4);
TASK_PP(16'h16E20,4);
TASK_PP(16'h16E21,4);
TASK_PP(16'h16E22,4);
TASK_PP(16'h16E23,4);
TASK_PP(16'h16E24,4);
TASK_PP(16'h16E25,4);
TASK_PP(16'h16E26,4);
TASK_PP(16'h16E27,4);
TASK_PP(16'h16E28,4);
TASK_PP(16'h16E29,4);
TASK_PP(16'h16E2A,4);
TASK_PP(16'h16E2B,4);
TASK_PP(16'h16E2C,4);
TASK_PP(16'h16E2D,4);
TASK_PP(16'h16E2E,4);
TASK_PP(16'h16E2F,4);
TASK_PP(16'h16E30,4);
TASK_PP(16'h16E31,4);
TASK_PP(16'h16E32,4);
TASK_PP(16'h16E33,4);
TASK_PP(16'h16E34,4);
TASK_PP(16'h16E35,4);
TASK_PP(16'h16E36,4);
TASK_PP(16'h16E37,4);
TASK_PP(16'h16E38,4);
TASK_PP(16'h16E39,4);
TASK_PP(16'h16E3A,4);
TASK_PP(16'h16E3B,4);
TASK_PP(16'h16E3C,4);
TASK_PP(16'h16E3D,4);
TASK_PP(16'h16E3E,4);
TASK_PP(16'h16E3F,4);
TASK_PP(16'h16E40,4);
TASK_PP(16'h16E41,4);
TASK_PP(16'h16E42,4);
TASK_PP(16'h16E43,4);
TASK_PP(16'h16E44,4);
TASK_PP(16'h16E45,4);
TASK_PP(16'h16E46,4);
TASK_PP(16'h16E47,4);
TASK_PP(16'h16E48,4);
TASK_PP(16'h16E49,4);
TASK_PP(16'h16E4A,4);
TASK_PP(16'h16E4B,4);
TASK_PP(16'h16E4C,4);
TASK_PP(16'h16E4D,4);
TASK_PP(16'h16E4E,4);
TASK_PP(16'h16E4F,4);
TASK_PP(16'h16E50,4);
TASK_PP(16'h16E51,4);
TASK_PP(16'h16E52,4);
TASK_PP(16'h16E53,4);
TASK_PP(16'h16E54,4);
TASK_PP(16'h16E55,4);
TASK_PP(16'h16E56,4);
TASK_PP(16'h16E57,4);
TASK_PP(16'h16E58,4);
TASK_PP(16'h16E59,4);
TASK_PP(16'h16E5A,4);
TASK_PP(16'h16E5B,4);
TASK_PP(16'h16E5C,4);
TASK_PP(16'h16E5D,4);
TASK_PP(16'h16E5E,4);
TASK_PP(16'h16E5F,4);
TASK_PP(16'h16E60,4);
TASK_PP(16'h16E61,4);
TASK_PP(16'h16E62,4);
TASK_PP(16'h16E63,4);
TASK_PP(16'h16E64,4);
TASK_PP(16'h16E65,4);
TASK_PP(16'h16E66,4);
TASK_PP(16'h16E67,4);
TASK_PP(16'h16E68,4);
TASK_PP(16'h16E69,4);
TASK_PP(16'h16E6A,4);
TASK_PP(16'h16E6B,4);
TASK_PP(16'h16E6C,4);
TASK_PP(16'h16E6D,4);
TASK_PP(16'h16E6E,4);
TASK_PP(16'h16E6F,4);
TASK_PP(16'h16E70,4);
TASK_PP(16'h16E71,4);
TASK_PP(16'h16E72,4);
TASK_PP(16'h16E73,4);
TASK_PP(16'h16E74,4);
TASK_PP(16'h16E75,4);
TASK_PP(16'h16E76,4);
TASK_PP(16'h16E77,4);
TASK_PP(16'h16E78,4);
TASK_PP(16'h16E79,4);
TASK_PP(16'h16E7A,4);
TASK_PP(16'h16E7B,4);
TASK_PP(16'h16E7C,4);
TASK_PP(16'h16E7D,4);
TASK_PP(16'h16E7E,4);
TASK_PP(16'h16E7F,4);
TASK_PP(16'h16E80,4);
TASK_PP(16'h16E81,4);
TASK_PP(16'h16E82,4);
TASK_PP(16'h16E83,4);
TASK_PP(16'h16E84,4);
TASK_PP(16'h16E85,4);
TASK_PP(16'h16E86,4);
TASK_PP(16'h16E87,4);
TASK_PP(16'h16E88,4);
TASK_PP(16'h16E89,4);
TASK_PP(16'h16E8A,4);
TASK_PP(16'h16E8B,4);
TASK_PP(16'h16E8C,4);
TASK_PP(16'h16E8D,4);
TASK_PP(16'h16E8E,4);
TASK_PP(16'h16E8F,4);
TASK_PP(16'h16E90,4);
TASK_PP(16'h16E91,4);
TASK_PP(16'h16E92,4);
TASK_PP(16'h16E93,4);
TASK_PP(16'h16E94,4);
TASK_PP(16'h16E95,4);
TASK_PP(16'h16E96,4);
TASK_PP(16'h16E97,4);
TASK_PP(16'h16E98,4);
TASK_PP(16'h16E99,4);
TASK_PP(16'h16E9A,4);
TASK_PP(16'h16E9B,4);
TASK_PP(16'h16E9C,4);
TASK_PP(16'h16E9D,4);
TASK_PP(16'h16E9E,4);
TASK_PP(16'h16E9F,4);
TASK_PP(16'h16EA0,4);
TASK_PP(16'h16EA1,4);
TASK_PP(16'h16EA2,4);
TASK_PP(16'h16EA3,4);
TASK_PP(16'h16EA4,4);
TASK_PP(16'h16EA5,4);
TASK_PP(16'h16EA6,4);
TASK_PP(16'h16EA7,4);
TASK_PP(16'h16EA8,4);
TASK_PP(16'h16EA9,4);
TASK_PP(16'h16EAA,4);
TASK_PP(16'h16EAB,4);
TASK_PP(16'h16EAC,4);
TASK_PP(16'h16EAD,4);
TASK_PP(16'h16EAE,4);
TASK_PP(16'h16EAF,4);
TASK_PP(16'h16EB0,4);
TASK_PP(16'h16EB1,4);
TASK_PP(16'h16EB2,4);
TASK_PP(16'h16EB3,4);
TASK_PP(16'h16EB4,4);
TASK_PP(16'h16EB5,4);
TASK_PP(16'h16EB6,4);
TASK_PP(16'h16EB7,4);
TASK_PP(16'h16EB8,4);
TASK_PP(16'h16EB9,4);
TASK_PP(16'h16EBA,4);
TASK_PP(16'h16EBB,4);
TASK_PP(16'h16EBC,4);
TASK_PP(16'h16EBD,4);
TASK_PP(16'h16EBE,4);
TASK_PP(16'h16EBF,4);
TASK_PP(16'h16EC0,4);
TASK_PP(16'h16EC1,4);
TASK_PP(16'h16EC2,4);
TASK_PP(16'h16EC3,4);
TASK_PP(16'h16EC4,4);
TASK_PP(16'h16EC5,4);
TASK_PP(16'h16EC6,4);
TASK_PP(16'h16EC7,4);
TASK_PP(16'h16EC8,4);
TASK_PP(16'h16EC9,4);
TASK_PP(16'h16ECA,4);
TASK_PP(16'h16ECB,4);
TASK_PP(16'h16ECC,4);
TASK_PP(16'h16ECD,4);
TASK_PP(16'h16ECE,4);
TASK_PP(16'h16ECF,4);
TASK_PP(16'h16ED0,4);
TASK_PP(16'h16ED1,4);
TASK_PP(16'h16ED2,4);
TASK_PP(16'h16ED3,4);
TASK_PP(16'h16ED4,4);
TASK_PP(16'h16ED5,4);
TASK_PP(16'h16ED6,4);
TASK_PP(16'h16ED7,4);
TASK_PP(16'h16ED8,4);
TASK_PP(16'h16ED9,4);
TASK_PP(16'h16EDA,4);
TASK_PP(16'h16EDB,4);
TASK_PP(16'h16EDC,4);
TASK_PP(16'h16EDD,4);
TASK_PP(16'h16EDE,4);
TASK_PP(16'h16EDF,4);
TASK_PP(16'h16EE0,4);
TASK_PP(16'h16EE1,4);
TASK_PP(16'h16EE2,4);
TASK_PP(16'h16EE3,4);
TASK_PP(16'h16EE4,4);
TASK_PP(16'h16EE5,4);
TASK_PP(16'h16EE6,4);
TASK_PP(16'h16EE7,4);
TASK_PP(16'h16EE8,4);
TASK_PP(16'h16EE9,4);
TASK_PP(16'h16EEA,4);
TASK_PP(16'h16EEB,4);
TASK_PP(16'h16EEC,4);
TASK_PP(16'h16EED,4);
TASK_PP(16'h16EEE,4);
TASK_PP(16'h16EEF,4);
TASK_PP(16'h16EF0,4);
TASK_PP(16'h16EF1,4);
TASK_PP(16'h16EF2,4);
TASK_PP(16'h16EF3,4);
TASK_PP(16'h16EF4,4);
TASK_PP(16'h16EF5,4);
TASK_PP(16'h16EF6,4);
TASK_PP(16'h16EF7,4);
TASK_PP(16'h16EF8,4);
TASK_PP(16'h16EF9,4);
TASK_PP(16'h16EFA,4);
TASK_PP(16'h16EFB,4);
TASK_PP(16'h16EFC,4);
TASK_PP(16'h16EFD,4);
TASK_PP(16'h16EFE,4);
TASK_PP(16'h16EFF,4);
TASK_PP(16'h16F00,4);
TASK_PP(16'h16F01,4);
TASK_PP(16'h16F02,4);
TASK_PP(16'h16F03,4);
TASK_PP(16'h16F04,4);
TASK_PP(16'h16F05,4);
TASK_PP(16'h16F06,4);
TASK_PP(16'h16F07,4);
TASK_PP(16'h16F08,4);
TASK_PP(16'h16F09,4);
TASK_PP(16'h16F0A,4);
TASK_PP(16'h16F0B,4);
TASK_PP(16'h16F0C,4);
TASK_PP(16'h16F0D,4);
TASK_PP(16'h16F0E,4);
TASK_PP(16'h16F0F,4);
TASK_PP(16'h16F10,4);
TASK_PP(16'h16F11,4);
TASK_PP(16'h16F12,4);
TASK_PP(16'h16F13,4);
TASK_PP(16'h16F14,4);
TASK_PP(16'h16F15,4);
TASK_PP(16'h16F16,4);
TASK_PP(16'h16F17,4);
TASK_PP(16'h16F18,4);
TASK_PP(16'h16F19,4);
TASK_PP(16'h16F1A,4);
TASK_PP(16'h16F1B,4);
TASK_PP(16'h16F1C,4);
TASK_PP(16'h16F1D,4);
TASK_PP(16'h16F1E,4);
TASK_PP(16'h16F1F,4);
TASK_PP(16'h16F20,4);
TASK_PP(16'h16F21,4);
TASK_PP(16'h16F22,4);
TASK_PP(16'h16F23,4);
TASK_PP(16'h16F24,4);
TASK_PP(16'h16F25,4);
TASK_PP(16'h16F26,4);
TASK_PP(16'h16F27,4);
TASK_PP(16'h16F28,4);
TASK_PP(16'h16F29,4);
TASK_PP(16'h16F2A,4);
TASK_PP(16'h16F2B,4);
TASK_PP(16'h16F2C,4);
TASK_PP(16'h16F2D,4);
TASK_PP(16'h16F2E,4);
TASK_PP(16'h16F2F,4);
TASK_PP(16'h16F30,4);
TASK_PP(16'h16F31,4);
TASK_PP(16'h16F32,4);
TASK_PP(16'h16F33,4);
TASK_PP(16'h16F34,4);
TASK_PP(16'h16F35,4);
TASK_PP(16'h16F36,4);
TASK_PP(16'h16F37,4);
TASK_PP(16'h16F38,4);
TASK_PP(16'h16F39,4);
TASK_PP(16'h16F3A,4);
TASK_PP(16'h16F3B,4);
TASK_PP(16'h16F3C,4);
TASK_PP(16'h16F3D,4);
TASK_PP(16'h16F3E,4);
TASK_PP(16'h16F3F,4);
TASK_PP(16'h16F40,4);
TASK_PP(16'h16F41,4);
TASK_PP(16'h16F42,4);
TASK_PP(16'h16F43,4);
TASK_PP(16'h16F44,4);
TASK_PP(16'h16F45,4);
TASK_PP(16'h16F46,4);
TASK_PP(16'h16F47,4);
TASK_PP(16'h16F48,4);
TASK_PP(16'h16F49,4);
TASK_PP(16'h16F4A,4);
TASK_PP(16'h16F4B,4);
TASK_PP(16'h16F4C,4);
TASK_PP(16'h16F4D,4);
TASK_PP(16'h16F4E,4);
TASK_PP(16'h16F4F,4);
TASK_PP(16'h16F50,4);
TASK_PP(16'h16F51,4);
TASK_PP(16'h16F52,4);
TASK_PP(16'h16F53,4);
TASK_PP(16'h16F54,4);
TASK_PP(16'h16F55,4);
TASK_PP(16'h16F56,4);
TASK_PP(16'h16F57,4);
TASK_PP(16'h16F58,4);
TASK_PP(16'h16F59,4);
TASK_PP(16'h16F5A,4);
TASK_PP(16'h16F5B,4);
TASK_PP(16'h16F5C,4);
TASK_PP(16'h16F5D,4);
TASK_PP(16'h16F5E,4);
TASK_PP(16'h16F5F,4);
TASK_PP(16'h16F60,4);
TASK_PP(16'h16F61,4);
TASK_PP(16'h16F62,4);
TASK_PP(16'h16F63,4);
TASK_PP(16'h16F64,4);
TASK_PP(16'h16F65,4);
TASK_PP(16'h16F66,4);
TASK_PP(16'h16F67,4);
TASK_PP(16'h16F68,4);
TASK_PP(16'h16F69,4);
TASK_PP(16'h16F6A,4);
TASK_PP(16'h16F6B,4);
TASK_PP(16'h16F6C,4);
TASK_PP(16'h16F6D,4);
TASK_PP(16'h16F6E,4);
TASK_PP(16'h16F6F,4);
TASK_PP(16'h16F70,4);
TASK_PP(16'h16F71,4);
TASK_PP(16'h16F72,4);
TASK_PP(16'h16F73,4);
TASK_PP(16'h16F74,4);
TASK_PP(16'h16F75,4);
TASK_PP(16'h16F76,4);
TASK_PP(16'h16F77,4);
TASK_PP(16'h16F78,4);
TASK_PP(16'h16F79,4);
TASK_PP(16'h16F7A,4);
TASK_PP(16'h16F7B,4);
TASK_PP(16'h16F7C,4);
TASK_PP(16'h16F7D,4);
TASK_PP(16'h16F7E,4);
TASK_PP(16'h16F7F,4);
TASK_PP(16'h16F80,4);
TASK_PP(16'h16F81,4);
TASK_PP(16'h16F82,4);
TASK_PP(16'h16F83,4);
TASK_PP(16'h16F84,4);
TASK_PP(16'h16F85,4);
TASK_PP(16'h16F86,4);
TASK_PP(16'h16F87,4);
TASK_PP(16'h16F88,4);
TASK_PP(16'h16F89,4);
TASK_PP(16'h16F8A,4);
TASK_PP(16'h16F8B,4);
TASK_PP(16'h16F8C,4);
TASK_PP(16'h16F8D,4);
TASK_PP(16'h16F8E,4);
TASK_PP(16'h16F8F,4);
TASK_PP(16'h16F90,4);
TASK_PP(16'h16F91,4);
TASK_PP(16'h16F92,4);
TASK_PP(16'h16F93,4);
TASK_PP(16'h16F94,4);
TASK_PP(16'h16F95,4);
TASK_PP(16'h16F96,4);
TASK_PP(16'h16F97,4);
TASK_PP(16'h16F98,4);
TASK_PP(16'h16F99,4);
TASK_PP(16'h16F9A,4);
TASK_PP(16'h16F9B,4);
TASK_PP(16'h16F9C,4);
TASK_PP(16'h16F9D,4);
TASK_PP(16'h16F9E,4);
TASK_PP(16'h16F9F,4);
TASK_PP(16'h16FA0,4);
TASK_PP(16'h16FA1,4);
TASK_PP(16'h16FA2,4);
TASK_PP(16'h16FA3,4);
TASK_PP(16'h16FA4,4);
TASK_PP(16'h16FA5,4);
TASK_PP(16'h16FA6,4);
TASK_PP(16'h16FA7,4);
TASK_PP(16'h16FA8,4);
TASK_PP(16'h16FA9,4);
TASK_PP(16'h16FAA,4);
TASK_PP(16'h16FAB,4);
TASK_PP(16'h16FAC,4);
TASK_PP(16'h16FAD,4);
TASK_PP(16'h16FAE,4);
TASK_PP(16'h16FAF,4);
TASK_PP(16'h16FB0,4);
TASK_PP(16'h16FB1,4);
TASK_PP(16'h16FB2,4);
TASK_PP(16'h16FB3,4);
TASK_PP(16'h16FB4,4);
TASK_PP(16'h16FB5,4);
TASK_PP(16'h16FB6,4);
TASK_PP(16'h16FB7,4);
TASK_PP(16'h16FB8,4);
TASK_PP(16'h16FB9,4);
TASK_PP(16'h16FBA,4);
TASK_PP(16'h16FBB,4);
TASK_PP(16'h16FBC,4);
TASK_PP(16'h16FBD,4);
TASK_PP(16'h16FBE,4);
TASK_PP(16'h16FBF,4);
TASK_PP(16'h16FC0,4);
TASK_PP(16'h16FC1,4);
TASK_PP(16'h16FC2,4);
TASK_PP(16'h16FC3,4);
TASK_PP(16'h16FC4,4);
TASK_PP(16'h16FC5,4);
TASK_PP(16'h16FC6,4);
TASK_PP(16'h16FC7,4);
TASK_PP(16'h16FC8,4);
TASK_PP(16'h16FC9,4);
TASK_PP(16'h16FCA,4);
TASK_PP(16'h16FCB,4);
TASK_PP(16'h16FCC,4);
TASK_PP(16'h16FCD,4);
TASK_PP(16'h16FCE,4);
TASK_PP(16'h16FCF,4);
TASK_PP(16'h16FD0,4);
TASK_PP(16'h16FD1,4);
TASK_PP(16'h16FD2,4);
TASK_PP(16'h16FD3,4);
TASK_PP(16'h16FD4,4);
TASK_PP(16'h16FD5,4);
TASK_PP(16'h16FD6,4);
TASK_PP(16'h16FD7,4);
TASK_PP(16'h16FD8,4);
TASK_PP(16'h16FD9,4);
TASK_PP(16'h16FDA,4);
TASK_PP(16'h16FDB,4);
TASK_PP(16'h16FDC,4);
TASK_PP(16'h16FDD,4);
TASK_PP(16'h16FDE,4);
TASK_PP(16'h16FDF,4);
TASK_PP(16'h16FE0,4);
TASK_PP(16'h16FE1,4);
TASK_PP(16'h16FE2,4);
TASK_PP(16'h16FE3,4);
TASK_PP(16'h16FE4,4);
TASK_PP(16'h16FE5,4);
TASK_PP(16'h16FE6,4);
TASK_PP(16'h16FE7,4);
TASK_PP(16'h16FE8,4);
TASK_PP(16'h16FE9,4);
TASK_PP(16'h16FEA,4);
TASK_PP(16'h16FEB,4);
TASK_PP(16'h16FEC,4);
TASK_PP(16'h16FED,4);
TASK_PP(16'h16FEE,4);
TASK_PP(16'h16FEF,4);
TASK_PP(16'h16FF0,4);
TASK_PP(16'h16FF1,4);
TASK_PP(16'h16FF2,4);
TASK_PP(16'h16FF3,4);
TASK_PP(16'h16FF4,4);
TASK_PP(16'h16FF5,4);
TASK_PP(16'h16FF6,4);
TASK_PP(16'h16FF7,4);
TASK_PP(16'h16FF8,4);
TASK_PP(16'h16FF9,4);
TASK_PP(16'h16FFA,4);
TASK_PP(16'h16FFB,4);
TASK_PP(16'h16FFC,4);
TASK_PP(16'h16FFD,4);
TASK_PP(16'h16FFE,4);
TASK_PP(16'h16FFF,4);
TASK_PP(16'h17000,4);
TASK_PP(16'h17001,4);
TASK_PP(16'h17002,4);
TASK_PP(16'h17003,4);
TASK_PP(16'h17004,4);
TASK_PP(16'h17005,4);
TASK_PP(16'h17006,4);
TASK_PP(16'h17007,4);
TASK_PP(16'h17008,4);
TASK_PP(16'h17009,4);
TASK_PP(16'h1700A,4);
TASK_PP(16'h1700B,4);
TASK_PP(16'h1700C,4);
TASK_PP(16'h1700D,4);
TASK_PP(16'h1700E,4);
TASK_PP(16'h1700F,4);
TASK_PP(16'h17010,4);
TASK_PP(16'h17011,4);
TASK_PP(16'h17012,4);
TASK_PP(16'h17013,4);
TASK_PP(16'h17014,4);
TASK_PP(16'h17015,4);
TASK_PP(16'h17016,4);
TASK_PP(16'h17017,4);
TASK_PP(16'h17018,4);
TASK_PP(16'h17019,4);
TASK_PP(16'h1701A,4);
TASK_PP(16'h1701B,4);
TASK_PP(16'h1701C,4);
TASK_PP(16'h1701D,4);
TASK_PP(16'h1701E,4);
TASK_PP(16'h1701F,4);
TASK_PP(16'h17020,4);
TASK_PP(16'h17021,4);
TASK_PP(16'h17022,4);
TASK_PP(16'h17023,4);
TASK_PP(16'h17024,4);
TASK_PP(16'h17025,4);
TASK_PP(16'h17026,4);
TASK_PP(16'h17027,4);
TASK_PP(16'h17028,4);
TASK_PP(16'h17029,4);
TASK_PP(16'h1702A,4);
TASK_PP(16'h1702B,4);
TASK_PP(16'h1702C,4);
TASK_PP(16'h1702D,4);
TASK_PP(16'h1702E,4);
TASK_PP(16'h1702F,4);
TASK_PP(16'h17030,4);
TASK_PP(16'h17031,4);
TASK_PP(16'h17032,4);
TASK_PP(16'h17033,4);
TASK_PP(16'h17034,4);
TASK_PP(16'h17035,4);
TASK_PP(16'h17036,4);
TASK_PP(16'h17037,4);
TASK_PP(16'h17038,4);
TASK_PP(16'h17039,4);
TASK_PP(16'h1703A,4);
TASK_PP(16'h1703B,4);
TASK_PP(16'h1703C,4);
TASK_PP(16'h1703D,4);
TASK_PP(16'h1703E,4);
TASK_PP(16'h1703F,4);
TASK_PP(16'h17040,4);
TASK_PP(16'h17041,4);
TASK_PP(16'h17042,4);
TASK_PP(16'h17043,4);
TASK_PP(16'h17044,4);
TASK_PP(16'h17045,4);
TASK_PP(16'h17046,4);
TASK_PP(16'h17047,4);
TASK_PP(16'h17048,4);
TASK_PP(16'h17049,4);
TASK_PP(16'h1704A,4);
TASK_PP(16'h1704B,4);
TASK_PP(16'h1704C,4);
TASK_PP(16'h1704D,4);
TASK_PP(16'h1704E,4);
TASK_PP(16'h1704F,4);
TASK_PP(16'h17050,4);
TASK_PP(16'h17051,4);
TASK_PP(16'h17052,4);
TASK_PP(16'h17053,4);
TASK_PP(16'h17054,4);
TASK_PP(16'h17055,4);
TASK_PP(16'h17056,4);
TASK_PP(16'h17057,4);
TASK_PP(16'h17058,4);
TASK_PP(16'h17059,4);
TASK_PP(16'h1705A,4);
TASK_PP(16'h1705B,4);
TASK_PP(16'h1705C,4);
TASK_PP(16'h1705D,4);
TASK_PP(16'h1705E,4);
TASK_PP(16'h1705F,4);
TASK_PP(16'h17060,4);
TASK_PP(16'h17061,4);
TASK_PP(16'h17062,4);
TASK_PP(16'h17063,4);
TASK_PP(16'h17064,4);
TASK_PP(16'h17065,4);
TASK_PP(16'h17066,4);
TASK_PP(16'h17067,4);
TASK_PP(16'h17068,4);
TASK_PP(16'h17069,4);
TASK_PP(16'h1706A,4);
TASK_PP(16'h1706B,4);
TASK_PP(16'h1706C,4);
TASK_PP(16'h1706D,4);
TASK_PP(16'h1706E,4);
TASK_PP(16'h1706F,4);
TASK_PP(16'h17070,4);
TASK_PP(16'h17071,4);
TASK_PP(16'h17072,4);
TASK_PP(16'h17073,4);
TASK_PP(16'h17074,4);
TASK_PP(16'h17075,4);
TASK_PP(16'h17076,4);
TASK_PP(16'h17077,4);
TASK_PP(16'h17078,4);
TASK_PP(16'h17079,4);
TASK_PP(16'h1707A,4);
TASK_PP(16'h1707B,4);
TASK_PP(16'h1707C,4);
TASK_PP(16'h1707D,4);
TASK_PP(16'h1707E,4);
TASK_PP(16'h1707F,4);
TASK_PP(16'h17080,4);
TASK_PP(16'h17081,4);
TASK_PP(16'h17082,4);
TASK_PP(16'h17083,4);
TASK_PP(16'h17084,4);
TASK_PP(16'h17085,4);
TASK_PP(16'h17086,4);
TASK_PP(16'h17087,4);
TASK_PP(16'h17088,4);
TASK_PP(16'h17089,4);
TASK_PP(16'h1708A,4);
TASK_PP(16'h1708B,4);
TASK_PP(16'h1708C,4);
TASK_PP(16'h1708D,4);
TASK_PP(16'h1708E,4);
TASK_PP(16'h1708F,4);
TASK_PP(16'h17090,4);
TASK_PP(16'h17091,4);
TASK_PP(16'h17092,4);
TASK_PP(16'h17093,4);
TASK_PP(16'h17094,4);
TASK_PP(16'h17095,4);
TASK_PP(16'h17096,4);
TASK_PP(16'h17097,4);
TASK_PP(16'h17098,4);
TASK_PP(16'h17099,4);
TASK_PP(16'h1709A,4);
TASK_PP(16'h1709B,4);
TASK_PP(16'h1709C,4);
TASK_PP(16'h1709D,4);
TASK_PP(16'h1709E,4);
TASK_PP(16'h1709F,4);
TASK_PP(16'h170A0,4);
TASK_PP(16'h170A1,4);
TASK_PP(16'h170A2,4);
TASK_PP(16'h170A3,4);
TASK_PP(16'h170A4,4);
TASK_PP(16'h170A5,4);
TASK_PP(16'h170A6,4);
TASK_PP(16'h170A7,4);
TASK_PP(16'h170A8,4);
TASK_PP(16'h170A9,4);
TASK_PP(16'h170AA,4);
TASK_PP(16'h170AB,4);
TASK_PP(16'h170AC,4);
TASK_PP(16'h170AD,4);
TASK_PP(16'h170AE,4);
TASK_PP(16'h170AF,4);
TASK_PP(16'h170B0,4);
TASK_PP(16'h170B1,4);
TASK_PP(16'h170B2,4);
TASK_PP(16'h170B3,4);
TASK_PP(16'h170B4,4);
TASK_PP(16'h170B5,4);
TASK_PP(16'h170B6,4);
TASK_PP(16'h170B7,4);
TASK_PP(16'h170B8,4);
TASK_PP(16'h170B9,4);
TASK_PP(16'h170BA,4);
TASK_PP(16'h170BB,4);
TASK_PP(16'h170BC,4);
TASK_PP(16'h170BD,4);
TASK_PP(16'h170BE,4);
TASK_PP(16'h170BF,4);
TASK_PP(16'h170C0,4);
TASK_PP(16'h170C1,4);
TASK_PP(16'h170C2,4);
TASK_PP(16'h170C3,4);
TASK_PP(16'h170C4,4);
TASK_PP(16'h170C5,4);
TASK_PP(16'h170C6,4);
TASK_PP(16'h170C7,4);
TASK_PP(16'h170C8,4);
TASK_PP(16'h170C9,4);
TASK_PP(16'h170CA,4);
TASK_PP(16'h170CB,4);
TASK_PP(16'h170CC,4);
TASK_PP(16'h170CD,4);
TASK_PP(16'h170CE,4);
TASK_PP(16'h170CF,4);
TASK_PP(16'h170D0,4);
TASK_PP(16'h170D1,4);
TASK_PP(16'h170D2,4);
TASK_PP(16'h170D3,4);
TASK_PP(16'h170D4,4);
TASK_PP(16'h170D5,4);
TASK_PP(16'h170D6,4);
TASK_PP(16'h170D7,4);
TASK_PP(16'h170D8,4);
TASK_PP(16'h170D9,4);
TASK_PP(16'h170DA,4);
TASK_PP(16'h170DB,4);
TASK_PP(16'h170DC,4);
TASK_PP(16'h170DD,4);
TASK_PP(16'h170DE,4);
TASK_PP(16'h170DF,4);
TASK_PP(16'h170E0,4);
TASK_PP(16'h170E1,4);
TASK_PP(16'h170E2,4);
TASK_PP(16'h170E3,4);
TASK_PP(16'h170E4,4);
TASK_PP(16'h170E5,4);
TASK_PP(16'h170E6,4);
TASK_PP(16'h170E7,4);
TASK_PP(16'h170E8,4);
TASK_PP(16'h170E9,4);
TASK_PP(16'h170EA,4);
TASK_PP(16'h170EB,4);
TASK_PP(16'h170EC,4);
TASK_PP(16'h170ED,4);
TASK_PP(16'h170EE,4);
TASK_PP(16'h170EF,4);
TASK_PP(16'h170F0,4);
TASK_PP(16'h170F1,4);
TASK_PP(16'h170F2,4);
TASK_PP(16'h170F3,4);
TASK_PP(16'h170F4,4);
TASK_PP(16'h170F5,4);
TASK_PP(16'h170F6,4);
TASK_PP(16'h170F7,4);
TASK_PP(16'h170F8,4);
TASK_PP(16'h170F9,4);
TASK_PP(16'h170FA,4);
TASK_PP(16'h170FB,4);
TASK_PP(16'h170FC,4);
TASK_PP(16'h170FD,4);
TASK_PP(16'h170FE,4);
TASK_PP(16'h170FF,4);
TASK_PP(16'h17100,4);
TASK_PP(16'h17101,4);
TASK_PP(16'h17102,4);
TASK_PP(16'h17103,4);
TASK_PP(16'h17104,4);
TASK_PP(16'h17105,4);
TASK_PP(16'h17106,4);
TASK_PP(16'h17107,4);
TASK_PP(16'h17108,4);
TASK_PP(16'h17109,4);
TASK_PP(16'h1710A,4);
TASK_PP(16'h1710B,4);
TASK_PP(16'h1710C,4);
TASK_PP(16'h1710D,4);
TASK_PP(16'h1710E,4);
TASK_PP(16'h1710F,4);
TASK_PP(16'h17110,4);
TASK_PP(16'h17111,4);
TASK_PP(16'h17112,4);
TASK_PP(16'h17113,4);
TASK_PP(16'h17114,4);
TASK_PP(16'h17115,4);
TASK_PP(16'h17116,4);
TASK_PP(16'h17117,4);
TASK_PP(16'h17118,4);
TASK_PP(16'h17119,4);
TASK_PP(16'h1711A,4);
TASK_PP(16'h1711B,4);
TASK_PP(16'h1711C,4);
TASK_PP(16'h1711D,4);
TASK_PP(16'h1711E,4);
TASK_PP(16'h1711F,4);
TASK_PP(16'h17120,4);
TASK_PP(16'h17121,4);
TASK_PP(16'h17122,4);
TASK_PP(16'h17123,4);
TASK_PP(16'h17124,4);
TASK_PP(16'h17125,4);
TASK_PP(16'h17126,4);
TASK_PP(16'h17127,4);
TASK_PP(16'h17128,4);
TASK_PP(16'h17129,4);
TASK_PP(16'h1712A,4);
TASK_PP(16'h1712B,4);
TASK_PP(16'h1712C,4);
TASK_PP(16'h1712D,4);
TASK_PP(16'h1712E,4);
TASK_PP(16'h1712F,4);
TASK_PP(16'h17130,4);
TASK_PP(16'h17131,4);
TASK_PP(16'h17132,4);
TASK_PP(16'h17133,4);
TASK_PP(16'h17134,4);
TASK_PP(16'h17135,4);
TASK_PP(16'h17136,4);
TASK_PP(16'h17137,4);
TASK_PP(16'h17138,4);
TASK_PP(16'h17139,4);
TASK_PP(16'h1713A,4);
TASK_PP(16'h1713B,4);
TASK_PP(16'h1713C,4);
TASK_PP(16'h1713D,4);
TASK_PP(16'h1713E,4);
TASK_PP(16'h1713F,4);
TASK_PP(16'h17140,4);
TASK_PP(16'h17141,4);
TASK_PP(16'h17142,4);
TASK_PP(16'h17143,4);
TASK_PP(16'h17144,4);
TASK_PP(16'h17145,4);
TASK_PP(16'h17146,4);
TASK_PP(16'h17147,4);
TASK_PP(16'h17148,4);
TASK_PP(16'h17149,4);
TASK_PP(16'h1714A,4);
TASK_PP(16'h1714B,4);
TASK_PP(16'h1714C,4);
TASK_PP(16'h1714D,4);
TASK_PP(16'h1714E,4);
TASK_PP(16'h1714F,4);
TASK_PP(16'h17150,4);
TASK_PP(16'h17151,4);
TASK_PP(16'h17152,4);
TASK_PP(16'h17153,4);
TASK_PP(16'h17154,4);
TASK_PP(16'h17155,4);
TASK_PP(16'h17156,4);
TASK_PP(16'h17157,4);
TASK_PP(16'h17158,4);
TASK_PP(16'h17159,4);
TASK_PP(16'h1715A,4);
TASK_PP(16'h1715B,4);
TASK_PP(16'h1715C,4);
TASK_PP(16'h1715D,4);
TASK_PP(16'h1715E,4);
TASK_PP(16'h1715F,4);
TASK_PP(16'h17160,4);
TASK_PP(16'h17161,4);
TASK_PP(16'h17162,4);
TASK_PP(16'h17163,4);
TASK_PP(16'h17164,4);
TASK_PP(16'h17165,4);
TASK_PP(16'h17166,4);
TASK_PP(16'h17167,4);
TASK_PP(16'h17168,4);
TASK_PP(16'h17169,4);
TASK_PP(16'h1716A,4);
TASK_PP(16'h1716B,4);
TASK_PP(16'h1716C,4);
TASK_PP(16'h1716D,4);
TASK_PP(16'h1716E,4);
TASK_PP(16'h1716F,4);
TASK_PP(16'h17170,4);
TASK_PP(16'h17171,4);
TASK_PP(16'h17172,4);
TASK_PP(16'h17173,4);
TASK_PP(16'h17174,4);
TASK_PP(16'h17175,4);
TASK_PP(16'h17176,4);
TASK_PP(16'h17177,4);
TASK_PP(16'h17178,4);
TASK_PP(16'h17179,4);
TASK_PP(16'h1717A,4);
TASK_PP(16'h1717B,4);
TASK_PP(16'h1717C,4);
TASK_PP(16'h1717D,4);
TASK_PP(16'h1717E,4);
TASK_PP(16'h1717F,4);
TASK_PP(16'h17180,4);
TASK_PP(16'h17181,4);
TASK_PP(16'h17182,4);
TASK_PP(16'h17183,4);
TASK_PP(16'h17184,4);
TASK_PP(16'h17185,4);
TASK_PP(16'h17186,4);
TASK_PP(16'h17187,4);
TASK_PP(16'h17188,4);
TASK_PP(16'h17189,4);
TASK_PP(16'h1718A,4);
TASK_PP(16'h1718B,4);
TASK_PP(16'h1718C,4);
TASK_PP(16'h1718D,4);
TASK_PP(16'h1718E,4);
TASK_PP(16'h1718F,4);
TASK_PP(16'h17190,4);
TASK_PP(16'h17191,4);
TASK_PP(16'h17192,4);
TASK_PP(16'h17193,4);
TASK_PP(16'h17194,4);
TASK_PP(16'h17195,4);
TASK_PP(16'h17196,4);
TASK_PP(16'h17197,4);
TASK_PP(16'h17198,4);
TASK_PP(16'h17199,4);
TASK_PP(16'h1719A,4);
TASK_PP(16'h1719B,4);
TASK_PP(16'h1719C,4);
TASK_PP(16'h1719D,4);
TASK_PP(16'h1719E,4);
TASK_PP(16'h1719F,4);
TASK_PP(16'h171A0,4);
TASK_PP(16'h171A1,4);
TASK_PP(16'h171A2,4);
TASK_PP(16'h171A3,4);
TASK_PP(16'h171A4,4);
TASK_PP(16'h171A5,4);
TASK_PP(16'h171A6,4);
TASK_PP(16'h171A7,4);
TASK_PP(16'h171A8,4);
TASK_PP(16'h171A9,4);
TASK_PP(16'h171AA,4);
TASK_PP(16'h171AB,4);
TASK_PP(16'h171AC,4);
TASK_PP(16'h171AD,4);
TASK_PP(16'h171AE,4);
TASK_PP(16'h171AF,4);
TASK_PP(16'h171B0,4);
TASK_PP(16'h171B1,4);
TASK_PP(16'h171B2,4);
TASK_PP(16'h171B3,4);
TASK_PP(16'h171B4,4);
TASK_PP(16'h171B5,4);
TASK_PP(16'h171B6,4);
TASK_PP(16'h171B7,4);
TASK_PP(16'h171B8,4);
TASK_PP(16'h171B9,4);
TASK_PP(16'h171BA,4);
TASK_PP(16'h171BB,4);
TASK_PP(16'h171BC,4);
TASK_PP(16'h171BD,4);
TASK_PP(16'h171BE,4);
TASK_PP(16'h171BF,4);
TASK_PP(16'h171C0,4);
TASK_PP(16'h171C1,4);
TASK_PP(16'h171C2,4);
TASK_PP(16'h171C3,4);
TASK_PP(16'h171C4,4);
TASK_PP(16'h171C5,4);
TASK_PP(16'h171C6,4);
TASK_PP(16'h171C7,4);
TASK_PP(16'h171C8,4);
TASK_PP(16'h171C9,4);
TASK_PP(16'h171CA,4);
TASK_PP(16'h171CB,4);
TASK_PP(16'h171CC,4);
TASK_PP(16'h171CD,4);
TASK_PP(16'h171CE,4);
TASK_PP(16'h171CF,4);
TASK_PP(16'h171D0,4);
TASK_PP(16'h171D1,4);
TASK_PP(16'h171D2,4);
TASK_PP(16'h171D3,4);
TASK_PP(16'h171D4,4);
TASK_PP(16'h171D5,4);
TASK_PP(16'h171D6,4);
TASK_PP(16'h171D7,4);
TASK_PP(16'h171D8,4);
TASK_PP(16'h171D9,4);
TASK_PP(16'h171DA,4);
TASK_PP(16'h171DB,4);
TASK_PP(16'h171DC,4);
TASK_PP(16'h171DD,4);
TASK_PP(16'h171DE,4);
TASK_PP(16'h171DF,4);
TASK_PP(16'h171E0,4);
TASK_PP(16'h171E1,4);
TASK_PP(16'h171E2,4);
TASK_PP(16'h171E3,4);
TASK_PP(16'h171E4,4);
TASK_PP(16'h171E5,4);
TASK_PP(16'h171E6,4);
TASK_PP(16'h171E7,4);
TASK_PP(16'h171E8,4);
TASK_PP(16'h171E9,4);
TASK_PP(16'h171EA,4);
TASK_PP(16'h171EB,4);
TASK_PP(16'h171EC,4);
TASK_PP(16'h171ED,4);
TASK_PP(16'h171EE,4);
TASK_PP(16'h171EF,4);
TASK_PP(16'h171F0,4);
TASK_PP(16'h171F1,4);
TASK_PP(16'h171F2,4);
TASK_PP(16'h171F3,4);
TASK_PP(16'h171F4,4);
TASK_PP(16'h171F5,4);
TASK_PP(16'h171F6,4);
TASK_PP(16'h171F7,4);
TASK_PP(16'h171F8,4);
TASK_PP(16'h171F9,4);
TASK_PP(16'h171FA,4);
TASK_PP(16'h171FB,4);
TASK_PP(16'h171FC,4);
TASK_PP(16'h171FD,4);
TASK_PP(16'h171FE,4);
TASK_PP(16'h171FF,4);
TASK_PP(16'h17200,4);
TASK_PP(16'h17201,4);
TASK_PP(16'h17202,4);
TASK_PP(16'h17203,4);
TASK_PP(16'h17204,4);
TASK_PP(16'h17205,4);
TASK_PP(16'h17206,4);
TASK_PP(16'h17207,4);
TASK_PP(16'h17208,4);
TASK_PP(16'h17209,4);
TASK_PP(16'h1720A,4);
TASK_PP(16'h1720B,4);
TASK_PP(16'h1720C,4);
TASK_PP(16'h1720D,4);
TASK_PP(16'h1720E,4);
TASK_PP(16'h1720F,4);
TASK_PP(16'h17210,4);
TASK_PP(16'h17211,4);
TASK_PP(16'h17212,4);
TASK_PP(16'h17213,4);
TASK_PP(16'h17214,4);
TASK_PP(16'h17215,4);
TASK_PP(16'h17216,4);
TASK_PP(16'h17217,4);
TASK_PP(16'h17218,4);
TASK_PP(16'h17219,4);
TASK_PP(16'h1721A,4);
TASK_PP(16'h1721B,4);
TASK_PP(16'h1721C,4);
TASK_PP(16'h1721D,4);
TASK_PP(16'h1721E,4);
TASK_PP(16'h1721F,4);
TASK_PP(16'h17220,4);
TASK_PP(16'h17221,4);
TASK_PP(16'h17222,4);
TASK_PP(16'h17223,4);
TASK_PP(16'h17224,4);
TASK_PP(16'h17225,4);
TASK_PP(16'h17226,4);
TASK_PP(16'h17227,4);
TASK_PP(16'h17228,4);
TASK_PP(16'h17229,4);
TASK_PP(16'h1722A,4);
TASK_PP(16'h1722B,4);
TASK_PP(16'h1722C,4);
TASK_PP(16'h1722D,4);
TASK_PP(16'h1722E,4);
TASK_PP(16'h1722F,4);
TASK_PP(16'h17230,4);
TASK_PP(16'h17231,4);
TASK_PP(16'h17232,4);
TASK_PP(16'h17233,4);
TASK_PP(16'h17234,4);
TASK_PP(16'h17235,4);
TASK_PP(16'h17236,4);
TASK_PP(16'h17237,4);
TASK_PP(16'h17238,4);
TASK_PP(16'h17239,4);
TASK_PP(16'h1723A,4);
TASK_PP(16'h1723B,4);
TASK_PP(16'h1723C,4);
TASK_PP(16'h1723D,4);
TASK_PP(16'h1723E,4);
TASK_PP(16'h1723F,4);
TASK_PP(16'h17240,4);
TASK_PP(16'h17241,4);
TASK_PP(16'h17242,4);
TASK_PP(16'h17243,4);
TASK_PP(16'h17244,4);
TASK_PP(16'h17245,4);
TASK_PP(16'h17246,4);
TASK_PP(16'h17247,4);
TASK_PP(16'h17248,4);
TASK_PP(16'h17249,4);
TASK_PP(16'h1724A,4);
TASK_PP(16'h1724B,4);
TASK_PP(16'h1724C,4);
TASK_PP(16'h1724D,4);
TASK_PP(16'h1724E,4);
TASK_PP(16'h1724F,4);
TASK_PP(16'h17250,4);
TASK_PP(16'h17251,4);
TASK_PP(16'h17252,4);
TASK_PP(16'h17253,4);
TASK_PP(16'h17254,4);
TASK_PP(16'h17255,4);
TASK_PP(16'h17256,4);
TASK_PP(16'h17257,4);
TASK_PP(16'h17258,4);
TASK_PP(16'h17259,4);
TASK_PP(16'h1725A,4);
TASK_PP(16'h1725B,4);
TASK_PP(16'h1725C,4);
TASK_PP(16'h1725D,4);
TASK_PP(16'h1725E,4);
TASK_PP(16'h1725F,4);
TASK_PP(16'h17260,4);
TASK_PP(16'h17261,4);
TASK_PP(16'h17262,4);
TASK_PP(16'h17263,4);
TASK_PP(16'h17264,4);
TASK_PP(16'h17265,4);
TASK_PP(16'h17266,4);
TASK_PP(16'h17267,4);
TASK_PP(16'h17268,4);
TASK_PP(16'h17269,4);
TASK_PP(16'h1726A,4);
TASK_PP(16'h1726B,4);
TASK_PP(16'h1726C,4);
TASK_PP(16'h1726D,4);
TASK_PP(16'h1726E,4);
TASK_PP(16'h1726F,4);
TASK_PP(16'h17270,4);
TASK_PP(16'h17271,4);
TASK_PP(16'h17272,4);
TASK_PP(16'h17273,4);
TASK_PP(16'h17274,4);
TASK_PP(16'h17275,4);
TASK_PP(16'h17276,4);
TASK_PP(16'h17277,4);
TASK_PP(16'h17278,4);
TASK_PP(16'h17279,4);
TASK_PP(16'h1727A,4);
TASK_PP(16'h1727B,4);
TASK_PP(16'h1727C,4);
TASK_PP(16'h1727D,4);
TASK_PP(16'h1727E,4);
TASK_PP(16'h1727F,4);
TASK_PP(16'h17280,4);
TASK_PP(16'h17281,4);
TASK_PP(16'h17282,4);
TASK_PP(16'h17283,4);
TASK_PP(16'h17284,4);
TASK_PP(16'h17285,4);
TASK_PP(16'h17286,4);
TASK_PP(16'h17287,4);
TASK_PP(16'h17288,4);
TASK_PP(16'h17289,4);
TASK_PP(16'h1728A,4);
TASK_PP(16'h1728B,4);
TASK_PP(16'h1728C,4);
TASK_PP(16'h1728D,4);
TASK_PP(16'h1728E,4);
TASK_PP(16'h1728F,4);
TASK_PP(16'h17290,4);
TASK_PP(16'h17291,4);
TASK_PP(16'h17292,4);
TASK_PP(16'h17293,4);
TASK_PP(16'h17294,4);
TASK_PP(16'h17295,4);
TASK_PP(16'h17296,4);
TASK_PP(16'h17297,4);
TASK_PP(16'h17298,4);
TASK_PP(16'h17299,4);
TASK_PP(16'h1729A,4);
TASK_PP(16'h1729B,4);
TASK_PP(16'h1729C,4);
TASK_PP(16'h1729D,4);
TASK_PP(16'h1729E,4);
TASK_PP(16'h1729F,4);
TASK_PP(16'h172A0,4);
TASK_PP(16'h172A1,4);
TASK_PP(16'h172A2,4);
TASK_PP(16'h172A3,4);
TASK_PP(16'h172A4,4);
TASK_PP(16'h172A5,4);
TASK_PP(16'h172A6,4);
TASK_PP(16'h172A7,4);
TASK_PP(16'h172A8,4);
TASK_PP(16'h172A9,4);
TASK_PP(16'h172AA,4);
TASK_PP(16'h172AB,4);
TASK_PP(16'h172AC,4);
TASK_PP(16'h172AD,4);
TASK_PP(16'h172AE,4);
TASK_PP(16'h172AF,4);
TASK_PP(16'h172B0,4);
TASK_PP(16'h172B1,4);
TASK_PP(16'h172B2,4);
TASK_PP(16'h172B3,4);
TASK_PP(16'h172B4,4);
TASK_PP(16'h172B5,4);
TASK_PP(16'h172B6,4);
TASK_PP(16'h172B7,4);
TASK_PP(16'h172B8,4);
TASK_PP(16'h172B9,4);
TASK_PP(16'h172BA,4);
TASK_PP(16'h172BB,4);
TASK_PP(16'h172BC,4);
TASK_PP(16'h172BD,4);
TASK_PP(16'h172BE,4);
TASK_PP(16'h172BF,4);
TASK_PP(16'h172C0,4);
TASK_PP(16'h172C1,4);
TASK_PP(16'h172C2,4);
TASK_PP(16'h172C3,4);
TASK_PP(16'h172C4,4);
TASK_PP(16'h172C5,4);
TASK_PP(16'h172C6,4);
TASK_PP(16'h172C7,4);
TASK_PP(16'h172C8,4);
TASK_PP(16'h172C9,4);
TASK_PP(16'h172CA,4);
TASK_PP(16'h172CB,4);
TASK_PP(16'h172CC,4);
TASK_PP(16'h172CD,4);
TASK_PP(16'h172CE,4);
TASK_PP(16'h172CF,4);
TASK_PP(16'h172D0,4);
TASK_PP(16'h172D1,4);
TASK_PP(16'h172D2,4);
TASK_PP(16'h172D3,4);
TASK_PP(16'h172D4,4);
TASK_PP(16'h172D5,4);
TASK_PP(16'h172D6,4);
TASK_PP(16'h172D7,4);
TASK_PP(16'h172D8,4);
TASK_PP(16'h172D9,4);
TASK_PP(16'h172DA,4);
TASK_PP(16'h172DB,4);
TASK_PP(16'h172DC,4);
TASK_PP(16'h172DD,4);
TASK_PP(16'h172DE,4);
TASK_PP(16'h172DF,4);
TASK_PP(16'h172E0,4);
TASK_PP(16'h172E1,4);
TASK_PP(16'h172E2,4);
TASK_PP(16'h172E3,4);
TASK_PP(16'h172E4,4);
TASK_PP(16'h172E5,4);
TASK_PP(16'h172E6,4);
TASK_PP(16'h172E7,4);
TASK_PP(16'h172E8,4);
TASK_PP(16'h172E9,4);
TASK_PP(16'h172EA,4);
TASK_PP(16'h172EB,4);
TASK_PP(16'h172EC,4);
TASK_PP(16'h172ED,4);
TASK_PP(16'h172EE,4);
TASK_PP(16'h172EF,4);
TASK_PP(16'h172F0,4);
TASK_PP(16'h172F1,4);
TASK_PP(16'h172F2,4);
TASK_PP(16'h172F3,4);
TASK_PP(16'h172F4,4);
TASK_PP(16'h172F5,4);
TASK_PP(16'h172F6,4);
TASK_PP(16'h172F7,4);
TASK_PP(16'h172F8,4);
TASK_PP(16'h172F9,4);
TASK_PP(16'h172FA,4);
TASK_PP(16'h172FB,4);
TASK_PP(16'h172FC,4);
TASK_PP(16'h172FD,4);
TASK_PP(16'h172FE,4);
TASK_PP(16'h172FF,4);
TASK_PP(16'h17300,4);
TASK_PP(16'h17301,4);
TASK_PP(16'h17302,4);
TASK_PP(16'h17303,4);
TASK_PP(16'h17304,4);
TASK_PP(16'h17305,4);
TASK_PP(16'h17306,4);
TASK_PP(16'h17307,4);
TASK_PP(16'h17308,4);
TASK_PP(16'h17309,4);
TASK_PP(16'h1730A,4);
TASK_PP(16'h1730B,4);
TASK_PP(16'h1730C,4);
TASK_PP(16'h1730D,4);
TASK_PP(16'h1730E,4);
TASK_PP(16'h1730F,4);
TASK_PP(16'h17310,4);
TASK_PP(16'h17311,4);
TASK_PP(16'h17312,4);
TASK_PP(16'h17313,4);
TASK_PP(16'h17314,4);
TASK_PP(16'h17315,4);
TASK_PP(16'h17316,4);
TASK_PP(16'h17317,4);
TASK_PP(16'h17318,4);
TASK_PP(16'h17319,4);
TASK_PP(16'h1731A,4);
TASK_PP(16'h1731B,4);
TASK_PP(16'h1731C,4);
TASK_PP(16'h1731D,4);
TASK_PP(16'h1731E,4);
TASK_PP(16'h1731F,4);
TASK_PP(16'h17320,4);
TASK_PP(16'h17321,4);
TASK_PP(16'h17322,4);
TASK_PP(16'h17323,4);
TASK_PP(16'h17324,4);
TASK_PP(16'h17325,4);
TASK_PP(16'h17326,4);
TASK_PP(16'h17327,4);
TASK_PP(16'h17328,4);
TASK_PP(16'h17329,4);
TASK_PP(16'h1732A,4);
TASK_PP(16'h1732B,4);
TASK_PP(16'h1732C,4);
TASK_PP(16'h1732D,4);
TASK_PP(16'h1732E,4);
TASK_PP(16'h1732F,4);
TASK_PP(16'h17330,4);
TASK_PP(16'h17331,4);
TASK_PP(16'h17332,4);
TASK_PP(16'h17333,4);
TASK_PP(16'h17334,4);
TASK_PP(16'h17335,4);
TASK_PP(16'h17336,4);
TASK_PP(16'h17337,4);
TASK_PP(16'h17338,4);
TASK_PP(16'h17339,4);
TASK_PP(16'h1733A,4);
TASK_PP(16'h1733B,4);
TASK_PP(16'h1733C,4);
TASK_PP(16'h1733D,4);
TASK_PP(16'h1733E,4);
TASK_PP(16'h1733F,4);
TASK_PP(16'h17340,4);
TASK_PP(16'h17341,4);
TASK_PP(16'h17342,4);
TASK_PP(16'h17343,4);
TASK_PP(16'h17344,4);
TASK_PP(16'h17345,4);
TASK_PP(16'h17346,4);
TASK_PP(16'h17347,4);
TASK_PP(16'h17348,4);
TASK_PP(16'h17349,4);
TASK_PP(16'h1734A,4);
TASK_PP(16'h1734B,4);
TASK_PP(16'h1734C,4);
TASK_PP(16'h1734D,4);
TASK_PP(16'h1734E,4);
TASK_PP(16'h1734F,4);
TASK_PP(16'h17350,4);
TASK_PP(16'h17351,4);
TASK_PP(16'h17352,4);
TASK_PP(16'h17353,4);
TASK_PP(16'h17354,4);
TASK_PP(16'h17355,4);
TASK_PP(16'h17356,4);
TASK_PP(16'h17357,4);
TASK_PP(16'h17358,4);
TASK_PP(16'h17359,4);
TASK_PP(16'h1735A,4);
TASK_PP(16'h1735B,4);
TASK_PP(16'h1735C,4);
TASK_PP(16'h1735D,4);
TASK_PP(16'h1735E,4);
TASK_PP(16'h1735F,4);
TASK_PP(16'h17360,4);
TASK_PP(16'h17361,4);
TASK_PP(16'h17362,4);
TASK_PP(16'h17363,4);
TASK_PP(16'h17364,4);
TASK_PP(16'h17365,4);
TASK_PP(16'h17366,4);
TASK_PP(16'h17367,4);
TASK_PP(16'h17368,4);
TASK_PP(16'h17369,4);
TASK_PP(16'h1736A,4);
TASK_PP(16'h1736B,4);
TASK_PP(16'h1736C,4);
TASK_PP(16'h1736D,4);
TASK_PP(16'h1736E,4);
TASK_PP(16'h1736F,4);
TASK_PP(16'h17370,4);
TASK_PP(16'h17371,4);
TASK_PP(16'h17372,4);
TASK_PP(16'h17373,4);
TASK_PP(16'h17374,4);
TASK_PP(16'h17375,4);
TASK_PP(16'h17376,4);
TASK_PP(16'h17377,4);
TASK_PP(16'h17378,4);
TASK_PP(16'h17379,4);
TASK_PP(16'h1737A,4);
TASK_PP(16'h1737B,4);
TASK_PP(16'h1737C,4);
TASK_PP(16'h1737D,4);
TASK_PP(16'h1737E,4);
TASK_PP(16'h1737F,4);
TASK_PP(16'h17380,4);
TASK_PP(16'h17381,4);
TASK_PP(16'h17382,4);
TASK_PP(16'h17383,4);
TASK_PP(16'h17384,4);
TASK_PP(16'h17385,4);
TASK_PP(16'h17386,4);
TASK_PP(16'h17387,4);
TASK_PP(16'h17388,4);
TASK_PP(16'h17389,4);
TASK_PP(16'h1738A,4);
TASK_PP(16'h1738B,4);
TASK_PP(16'h1738C,4);
TASK_PP(16'h1738D,4);
TASK_PP(16'h1738E,4);
TASK_PP(16'h1738F,4);
TASK_PP(16'h17390,4);
TASK_PP(16'h17391,4);
TASK_PP(16'h17392,4);
TASK_PP(16'h17393,4);
TASK_PP(16'h17394,4);
TASK_PP(16'h17395,4);
TASK_PP(16'h17396,4);
TASK_PP(16'h17397,4);
TASK_PP(16'h17398,4);
TASK_PP(16'h17399,4);
TASK_PP(16'h1739A,4);
TASK_PP(16'h1739B,4);
TASK_PP(16'h1739C,4);
TASK_PP(16'h1739D,4);
TASK_PP(16'h1739E,4);
TASK_PP(16'h1739F,4);
TASK_PP(16'h173A0,4);
TASK_PP(16'h173A1,4);
TASK_PP(16'h173A2,4);
TASK_PP(16'h173A3,4);
TASK_PP(16'h173A4,4);
TASK_PP(16'h173A5,4);
TASK_PP(16'h173A6,4);
TASK_PP(16'h173A7,4);
TASK_PP(16'h173A8,4);
TASK_PP(16'h173A9,4);
TASK_PP(16'h173AA,4);
TASK_PP(16'h173AB,4);
TASK_PP(16'h173AC,4);
TASK_PP(16'h173AD,4);
TASK_PP(16'h173AE,4);
TASK_PP(16'h173AF,4);
TASK_PP(16'h173B0,4);
TASK_PP(16'h173B1,4);
TASK_PP(16'h173B2,4);
TASK_PP(16'h173B3,4);
TASK_PP(16'h173B4,4);
TASK_PP(16'h173B5,4);
TASK_PP(16'h173B6,4);
TASK_PP(16'h173B7,4);
TASK_PP(16'h173B8,4);
TASK_PP(16'h173B9,4);
TASK_PP(16'h173BA,4);
TASK_PP(16'h173BB,4);
TASK_PP(16'h173BC,4);
TASK_PP(16'h173BD,4);
TASK_PP(16'h173BE,4);
TASK_PP(16'h173BF,4);
TASK_PP(16'h173C0,4);
TASK_PP(16'h173C1,4);
TASK_PP(16'h173C2,4);
TASK_PP(16'h173C3,4);
TASK_PP(16'h173C4,4);
TASK_PP(16'h173C5,4);
TASK_PP(16'h173C6,4);
TASK_PP(16'h173C7,4);
TASK_PP(16'h173C8,4);
TASK_PP(16'h173C9,4);
TASK_PP(16'h173CA,4);
TASK_PP(16'h173CB,4);
TASK_PP(16'h173CC,4);
TASK_PP(16'h173CD,4);
TASK_PP(16'h173CE,4);
TASK_PP(16'h173CF,4);
TASK_PP(16'h173D0,4);
TASK_PP(16'h173D1,4);
TASK_PP(16'h173D2,4);
TASK_PP(16'h173D3,4);
TASK_PP(16'h173D4,4);
TASK_PP(16'h173D5,4);
TASK_PP(16'h173D6,4);
TASK_PP(16'h173D7,4);
TASK_PP(16'h173D8,4);
TASK_PP(16'h173D9,4);
TASK_PP(16'h173DA,4);
TASK_PP(16'h173DB,4);
TASK_PP(16'h173DC,4);
TASK_PP(16'h173DD,4);
TASK_PP(16'h173DE,4);
TASK_PP(16'h173DF,4);
TASK_PP(16'h173E0,4);
TASK_PP(16'h173E1,4);
TASK_PP(16'h173E2,4);
TASK_PP(16'h173E3,4);
TASK_PP(16'h173E4,4);
TASK_PP(16'h173E5,4);
TASK_PP(16'h173E6,4);
TASK_PP(16'h173E7,4);
TASK_PP(16'h173E8,4);
TASK_PP(16'h173E9,4);
TASK_PP(16'h173EA,4);
TASK_PP(16'h173EB,4);
TASK_PP(16'h173EC,4);
TASK_PP(16'h173ED,4);
TASK_PP(16'h173EE,4);
TASK_PP(16'h173EF,4);
TASK_PP(16'h173F0,4);
TASK_PP(16'h173F1,4);
TASK_PP(16'h173F2,4);
TASK_PP(16'h173F3,4);
TASK_PP(16'h173F4,4);
TASK_PP(16'h173F5,4);
TASK_PP(16'h173F6,4);
TASK_PP(16'h173F7,4);
TASK_PP(16'h173F8,4);
TASK_PP(16'h173F9,4);
TASK_PP(16'h173FA,4);
TASK_PP(16'h173FB,4);
TASK_PP(16'h173FC,4);
TASK_PP(16'h173FD,4);
TASK_PP(16'h173FE,4);
TASK_PP(16'h173FF,4);
TASK_PP(16'h17400,4);
TASK_PP(16'h17401,4);
TASK_PP(16'h17402,4);
TASK_PP(16'h17403,4);
TASK_PP(16'h17404,4);
TASK_PP(16'h17405,4);
TASK_PP(16'h17406,4);
TASK_PP(16'h17407,4);
TASK_PP(16'h17408,4);
TASK_PP(16'h17409,4);
TASK_PP(16'h1740A,4);
TASK_PP(16'h1740B,4);
TASK_PP(16'h1740C,4);
TASK_PP(16'h1740D,4);
TASK_PP(16'h1740E,4);
TASK_PP(16'h1740F,4);
TASK_PP(16'h17410,4);
TASK_PP(16'h17411,4);
TASK_PP(16'h17412,4);
TASK_PP(16'h17413,4);
TASK_PP(16'h17414,4);
TASK_PP(16'h17415,4);
TASK_PP(16'h17416,4);
TASK_PP(16'h17417,4);
TASK_PP(16'h17418,4);
TASK_PP(16'h17419,4);
TASK_PP(16'h1741A,4);
TASK_PP(16'h1741B,4);
TASK_PP(16'h1741C,4);
TASK_PP(16'h1741D,4);
TASK_PP(16'h1741E,4);
TASK_PP(16'h1741F,4);
TASK_PP(16'h17420,4);
TASK_PP(16'h17421,4);
TASK_PP(16'h17422,4);
TASK_PP(16'h17423,4);
TASK_PP(16'h17424,4);
TASK_PP(16'h17425,4);
TASK_PP(16'h17426,4);
TASK_PP(16'h17427,4);
TASK_PP(16'h17428,4);
TASK_PP(16'h17429,4);
TASK_PP(16'h1742A,4);
TASK_PP(16'h1742B,4);
TASK_PP(16'h1742C,4);
TASK_PP(16'h1742D,4);
TASK_PP(16'h1742E,4);
TASK_PP(16'h1742F,4);
TASK_PP(16'h17430,4);
TASK_PP(16'h17431,4);
TASK_PP(16'h17432,4);
TASK_PP(16'h17433,4);
TASK_PP(16'h17434,4);
TASK_PP(16'h17435,4);
TASK_PP(16'h17436,4);
TASK_PP(16'h17437,4);
TASK_PP(16'h17438,4);
TASK_PP(16'h17439,4);
TASK_PP(16'h1743A,4);
TASK_PP(16'h1743B,4);
TASK_PP(16'h1743C,4);
TASK_PP(16'h1743D,4);
TASK_PP(16'h1743E,4);
TASK_PP(16'h1743F,4);
TASK_PP(16'h17440,4);
TASK_PP(16'h17441,4);
TASK_PP(16'h17442,4);
TASK_PP(16'h17443,4);
TASK_PP(16'h17444,4);
TASK_PP(16'h17445,4);
TASK_PP(16'h17446,4);
TASK_PP(16'h17447,4);
TASK_PP(16'h17448,4);
TASK_PP(16'h17449,4);
TASK_PP(16'h1744A,4);
TASK_PP(16'h1744B,4);
TASK_PP(16'h1744C,4);
TASK_PP(16'h1744D,4);
TASK_PP(16'h1744E,4);
TASK_PP(16'h1744F,4);
TASK_PP(16'h17450,4);
TASK_PP(16'h17451,4);
TASK_PP(16'h17452,4);
TASK_PP(16'h17453,4);
TASK_PP(16'h17454,4);
TASK_PP(16'h17455,4);
TASK_PP(16'h17456,4);
TASK_PP(16'h17457,4);
TASK_PP(16'h17458,4);
TASK_PP(16'h17459,4);
TASK_PP(16'h1745A,4);
TASK_PP(16'h1745B,4);
TASK_PP(16'h1745C,4);
TASK_PP(16'h1745D,4);
TASK_PP(16'h1745E,4);
TASK_PP(16'h1745F,4);
TASK_PP(16'h17460,4);
TASK_PP(16'h17461,4);
TASK_PP(16'h17462,4);
TASK_PP(16'h17463,4);
TASK_PP(16'h17464,4);
TASK_PP(16'h17465,4);
TASK_PP(16'h17466,4);
TASK_PP(16'h17467,4);
TASK_PP(16'h17468,4);
TASK_PP(16'h17469,4);
TASK_PP(16'h1746A,4);
TASK_PP(16'h1746B,4);
TASK_PP(16'h1746C,4);
TASK_PP(16'h1746D,4);
TASK_PP(16'h1746E,4);
TASK_PP(16'h1746F,4);
TASK_PP(16'h17470,4);
TASK_PP(16'h17471,4);
TASK_PP(16'h17472,4);
TASK_PP(16'h17473,4);
TASK_PP(16'h17474,4);
TASK_PP(16'h17475,4);
TASK_PP(16'h17476,4);
TASK_PP(16'h17477,4);
TASK_PP(16'h17478,4);
TASK_PP(16'h17479,4);
TASK_PP(16'h1747A,4);
TASK_PP(16'h1747B,4);
TASK_PP(16'h1747C,4);
TASK_PP(16'h1747D,4);
TASK_PP(16'h1747E,4);
TASK_PP(16'h1747F,4);
TASK_PP(16'h17480,4);
TASK_PP(16'h17481,4);
TASK_PP(16'h17482,4);
TASK_PP(16'h17483,4);
TASK_PP(16'h17484,4);
TASK_PP(16'h17485,4);
TASK_PP(16'h17486,4);
TASK_PP(16'h17487,4);
TASK_PP(16'h17488,4);
TASK_PP(16'h17489,4);
TASK_PP(16'h1748A,4);
TASK_PP(16'h1748B,4);
TASK_PP(16'h1748C,4);
TASK_PP(16'h1748D,4);
TASK_PP(16'h1748E,4);
TASK_PP(16'h1748F,4);
TASK_PP(16'h17490,4);
TASK_PP(16'h17491,4);
TASK_PP(16'h17492,4);
TASK_PP(16'h17493,4);
TASK_PP(16'h17494,4);
TASK_PP(16'h17495,4);
TASK_PP(16'h17496,4);
TASK_PP(16'h17497,4);
TASK_PP(16'h17498,4);
TASK_PP(16'h17499,4);
TASK_PP(16'h1749A,4);
TASK_PP(16'h1749B,4);
TASK_PP(16'h1749C,4);
TASK_PP(16'h1749D,4);
TASK_PP(16'h1749E,4);
TASK_PP(16'h1749F,4);
TASK_PP(16'h174A0,4);
TASK_PP(16'h174A1,4);
TASK_PP(16'h174A2,4);
TASK_PP(16'h174A3,4);
TASK_PP(16'h174A4,4);
TASK_PP(16'h174A5,4);
TASK_PP(16'h174A6,4);
TASK_PP(16'h174A7,4);
TASK_PP(16'h174A8,4);
TASK_PP(16'h174A9,4);
TASK_PP(16'h174AA,4);
TASK_PP(16'h174AB,4);
TASK_PP(16'h174AC,4);
TASK_PP(16'h174AD,4);
TASK_PP(16'h174AE,4);
TASK_PP(16'h174AF,4);
TASK_PP(16'h174B0,4);
TASK_PP(16'h174B1,4);
TASK_PP(16'h174B2,4);
TASK_PP(16'h174B3,4);
TASK_PP(16'h174B4,4);
TASK_PP(16'h174B5,4);
TASK_PP(16'h174B6,4);
TASK_PP(16'h174B7,4);
TASK_PP(16'h174B8,4);
TASK_PP(16'h174B9,4);
TASK_PP(16'h174BA,4);
TASK_PP(16'h174BB,4);
TASK_PP(16'h174BC,4);
TASK_PP(16'h174BD,4);
TASK_PP(16'h174BE,4);
TASK_PP(16'h174BF,4);
TASK_PP(16'h174C0,4);
TASK_PP(16'h174C1,4);
TASK_PP(16'h174C2,4);
TASK_PP(16'h174C3,4);
TASK_PP(16'h174C4,4);
TASK_PP(16'h174C5,4);
TASK_PP(16'h174C6,4);
TASK_PP(16'h174C7,4);
TASK_PP(16'h174C8,4);
TASK_PP(16'h174C9,4);
TASK_PP(16'h174CA,4);
TASK_PP(16'h174CB,4);
TASK_PP(16'h174CC,4);
TASK_PP(16'h174CD,4);
TASK_PP(16'h174CE,4);
TASK_PP(16'h174CF,4);
TASK_PP(16'h174D0,4);
TASK_PP(16'h174D1,4);
TASK_PP(16'h174D2,4);
TASK_PP(16'h174D3,4);
TASK_PP(16'h174D4,4);
TASK_PP(16'h174D5,4);
TASK_PP(16'h174D6,4);
TASK_PP(16'h174D7,4);
TASK_PP(16'h174D8,4);
TASK_PP(16'h174D9,4);
TASK_PP(16'h174DA,4);
TASK_PP(16'h174DB,4);
TASK_PP(16'h174DC,4);
TASK_PP(16'h174DD,4);
TASK_PP(16'h174DE,4);
TASK_PP(16'h174DF,4);
TASK_PP(16'h174E0,4);
TASK_PP(16'h174E1,4);
TASK_PP(16'h174E2,4);
TASK_PP(16'h174E3,4);
TASK_PP(16'h174E4,4);
TASK_PP(16'h174E5,4);
TASK_PP(16'h174E6,4);
TASK_PP(16'h174E7,4);
TASK_PP(16'h174E8,4);
TASK_PP(16'h174E9,4);
TASK_PP(16'h174EA,4);
TASK_PP(16'h174EB,4);
TASK_PP(16'h174EC,4);
TASK_PP(16'h174ED,4);
TASK_PP(16'h174EE,4);
TASK_PP(16'h174EF,4);
TASK_PP(16'h174F0,4);
TASK_PP(16'h174F1,4);
TASK_PP(16'h174F2,4);
TASK_PP(16'h174F3,4);
TASK_PP(16'h174F4,4);
TASK_PP(16'h174F5,4);
TASK_PP(16'h174F6,4);
TASK_PP(16'h174F7,4);
TASK_PP(16'h174F8,4);
TASK_PP(16'h174F9,4);
TASK_PP(16'h174FA,4);
TASK_PP(16'h174FB,4);
TASK_PP(16'h174FC,4);
TASK_PP(16'h174FD,4);
TASK_PP(16'h174FE,4);
TASK_PP(16'h174FF,4);
TASK_PP(16'h17500,4);
TASK_PP(16'h17501,4);
TASK_PP(16'h17502,4);
TASK_PP(16'h17503,4);
TASK_PP(16'h17504,4);
TASK_PP(16'h17505,4);
TASK_PP(16'h17506,4);
TASK_PP(16'h17507,4);
TASK_PP(16'h17508,4);
TASK_PP(16'h17509,4);
TASK_PP(16'h1750A,4);
TASK_PP(16'h1750B,4);
TASK_PP(16'h1750C,4);
TASK_PP(16'h1750D,4);
TASK_PP(16'h1750E,4);
TASK_PP(16'h1750F,4);
TASK_PP(16'h17510,4);
TASK_PP(16'h17511,4);
TASK_PP(16'h17512,4);
TASK_PP(16'h17513,4);
TASK_PP(16'h17514,4);
TASK_PP(16'h17515,4);
TASK_PP(16'h17516,4);
TASK_PP(16'h17517,4);
TASK_PP(16'h17518,4);
TASK_PP(16'h17519,4);
TASK_PP(16'h1751A,4);
TASK_PP(16'h1751B,4);
TASK_PP(16'h1751C,4);
TASK_PP(16'h1751D,4);
TASK_PP(16'h1751E,4);
TASK_PP(16'h1751F,4);
TASK_PP(16'h17520,4);
TASK_PP(16'h17521,4);
TASK_PP(16'h17522,4);
TASK_PP(16'h17523,4);
TASK_PP(16'h17524,4);
TASK_PP(16'h17525,4);
TASK_PP(16'h17526,4);
TASK_PP(16'h17527,4);
TASK_PP(16'h17528,4);
TASK_PP(16'h17529,4);
TASK_PP(16'h1752A,4);
TASK_PP(16'h1752B,4);
TASK_PP(16'h1752C,4);
TASK_PP(16'h1752D,4);
TASK_PP(16'h1752E,4);
TASK_PP(16'h1752F,4);
TASK_PP(16'h17530,4);
TASK_PP(16'h17531,4);
TASK_PP(16'h17532,4);
TASK_PP(16'h17533,4);
TASK_PP(16'h17534,4);
TASK_PP(16'h17535,4);
TASK_PP(16'h17536,4);
TASK_PP(16'h17537,4);
TASK_PP(16'h17538,4);
TASK_PP(16'h17539,4);
TASK_PP(16'h1753A,4);
TASK_PP(16'h1753B,4);
TASK_PP(16'h1753C,4);
TASK_PP(16'h1753D,4);
TASK_PP(16'h1753E,4);
TASK_PP(16'h1753F,4);
TASK_PP(16'h17540,4);
TASK_PP(16'h17541,4);
TASK_PP(16'h17542,4);
TASK_PP(16'h17543,4);
TASK_PP(16'h17544,4);
TASK_PP(16'h17545,4);
TASK_PP(16'h17546,4);
TASK_PP(16'h17547,4);
TASK_PP(16'h17548,4);
TASK_PP(16'h17549,4);
TASK_PP(16'h1754A,4);
TASK_PP(16'h1754B,4);
TASK_PP(16'h1754C,4);
TASK_PP(16'h1754D,4);
TASK_PP(16'h1754E,4);
TASK_PP(16'h1754F,4);
TASK_PP(16'h17550,4);
TASK_PP(16'h17551,4);
TASK_PP(16'h17552,4);
TASK_PP(16'h17553,4);
TASK_PP(16'h17554,4);
TASK_PP(16'h17555,4);
TASK_PP(16'h17556,4);
TASK_PP(16'h17557,4);
TASK_PP(16'h17558,4);
TASK_PP(16'h17559,4);
TASK_PP(16'h1755A,4);
TASK_PP(16'h1755B,4);
TASK_PP(16'h1755C,4);
TASK_PP(16'h1755D,4);
TASK_PP(16'h1755E,4);
TASK_PP(16'h1755F,4);
TASK_PP(16'h17560,4);
TASK_PP(16'h17561,4);
TASK_PP(16'h17562,4);
TASK_PP(16'h17563,4);
TASK_PP(16'h17564,4);
TASK_PP(16'h17565,4);
TASK_PP(16'h17566,4);
TASK_PP(16'h17567,4);
TASK_PP(16'h17568,4);
TASK_PP(16'h17569,4);
TASK_PP(16'h1756A,4);
TASK_PP(16'h1756B,4);
TASK_PP(16'h1756C,4);
TASK_PP(16'h1756D,4);
TASK_PP(16'h1756E,4);
TASK_PP(16'h1756F,4);
TASK_PP(16'h17570,4);
TASK_PP(16'h17571,4);
TASK_PP(16'h17572,4);
TASK_PP(16'h17573,4);
TASK_PP(16'h17574,4);
TASK_PP(16'h17575,4);
TASK_PP(16'h17576,4);
TASK_PP(16'h17577,4);
TASK_PP(16'h17578,4);
TASK_PP(16'h17579,4);
TASK_PP(16'h1757A,4);
TASK_PP(16'h1757B,4);
TASK_PP(16'h1757C,4);
TASK_PP(16'h1757D,4);
TASK_PP(16'h1757E,4);
TASK_PP(16'h1757F,4);
TASK_PP(16'h17580,4);
TASK_PP(16'h17581,4);
TASK_PP(16'h17582,4);
TASK_PP(16'h17583,4);
TASK_PP(16'h17584,4);
TASK_PP(16'h17585,4);
TASK_PP(16'h17586,4);
TASK_PP(16'h17587,4);
TASK_PP(16'h17588,4);
TASK_PP(16'h17589,4);
TASK_PP(16'h1758A,4);
TASK_PP(16'h1758B,4);
TASK_PP(16'h1758C,4);
TASK_PP(16'h1758D,4);
TASK_PP(16'h1758E,4);
TASK_PP(16'h1758F,4);
TASK_PP(16'h17590,4);
TASK_PP(16'h17591,4);
TASK_PP(16'h17592,4);
TASK_PP(16'h17593,4);
TASK_PP(16'h17594,4);
TASK_PP(16'h17595,4);
TASK_PP(16'h17596,4);
TASK_PP(16'h17597,4);
TASK_PP(16'h17598,4);
TASK_PP(16'h17599,4);
TASK_PP(16'h1759A,4);
TASK_PP(16'h1759B,4);
TASK_PP(16'h1759C,4);
TASK_PP(16'h1759D,4);
TASK_PP(16'h1759E,4);
TASK_PP(16'h1759F,4);
TASK_PP(16'h175A0,4);
TASK_PP(16'h175A1,4);
TASK_PP(16'h175A2,4);
TASK_PP(16'h175A3,4);
TASK_PP(16'h175A4,4);
TASK_PP(16'h175A5,4);
TASK_PP(16'h175A6,4);
TASK_PP(16'h175A7,4);
TASK_PP(16'h175A8,4);
TASK_PP(16'h175A9,4);
TASK_PP(16'h175AA,4);
TASK_PP(16'h175AB,4);
TASK_PP(16'h175AC,4);
TASK_PP(16'h175AD,4);
TASK_PP(16'h175AE,4);
TASK_PP(16'h175AF,4);
TASK_PP(16'h175B0,4);
TASK_PP(16'h175B1,4);
TASK_PP(16'h175B2,4);
TASK_PP(16'h175B3,4);
TASK_PP(16'h175B4,4);
TASK_PP(16'h175B5,4);
TASK_PP(16'h175B6,4);
TASK_PP(16'h175B7,4);
TASK_PP(16'h175B8,4);
TASK_PP(16'h175B9,4);
TASK_PP(16'h175BA,4);
TASK_PP(16'h175BB,4);
TASK_PP(16'h175BC,4);
TASK_PP(16'h175BD,4);
TASK_PP(16'h175BE,4);
TASK_PP(16'h175BF,4);
TASK_PP(16'h175C0,4);
TASK_PP(16'h175C1,4);
TASK_PP(16'h175C2,4);
TASK_PP(16'h175C3,4);
TASK_PP(16'h175C4,4);
TASK_PP(16'h175C5,4);
TASK_PP(16'h175C6,4);
TASK_PP(16'h175C7,4);
TASK_PP(16'h175C8,4);
TASK_PP(16'h175C9,4);
TASK_PP(16'h175CA,4);
TASK_PP(16'h175CB,4);
TASK_PP(16'h175CC,4);
TASK_PP(16'h175CD,4);
TASK_PP(16'h175CE,4);
TASK_PP(16'h175CF,4);
TASK_PP(16'h175D0,4);
TASK_PP(16'h175D1,4);
TASK_PP(16'h175D2,4);
TASK_PP(16'h175D3,4);
TASK_PP(16'h175D4,4);
TASK_PP(16'h175D5,4);
TASK_PP(16'h175D6,4);
TASK_PP(16'h175D7,4);
TASK_PP(16'h175D8,4);
TASK_PP(16'h175D9,4);
TASK_PP(16'h175DA,4);
TASK_PP(16'h175DB,4);
TASK_PP(16'h175DC,4);
TASK_PP(16'h175DD,4);
TASK_PP(16'h175DE,4);
TASK_PP(16'h175DF,4);
TASK_PP(16'h175E0,4);
TASK_PP(16'h175E1,4);
TASK_PP(16'h175E2,4);
TASK_PP(16'h175E3,4);
TASK_PP(16'h175E4,4);
TASK_PP(16'h175E5,4);
TASK_PP(16'h175E6,4);
TASK_PP(16'h175E7,4);
TASK_PP(16'h175E8,4);
TASK_PP(16'h175E9,4);
TASK_PP(16'h175EA,4);
TASK_PP(16'h175EB,4);
TASK_PP(16'h175EC,4);
TASK_PP(16'h175ED,4);
TASK_PP(16'h175EE,4);
TASK_PP(16'h175EF,4);
TASK_PP(16'h175F0,4);
TASK_PP(16'h175F1,4);
TASK_PP(16'h175F2,4);
TASK_PP(16'h175F3,4);
TASK_PP(16'h175F4,4);
TASK_PP(16'h175F5,4);
TASK_PP(16'h175F6,4);
TASK_PP(16'h175F7,4);
TASK_PP(16'h175F8,4);
TASK_PP(16'h175F9,4);
TASK_PP(16'h175FA,4);
TASK_PP(16'h175FB,4);
TASK_PP(16'h175FC,4);
TASK_PP(16'h175FD,4);
TASK_PP(16'h175FE,4);
TASK_PP(16'h175FF,4);
TASK_PP(16'h17600,4);
TASK_PP(16'h17601,4);
TASK_PP(16'h17602,4);
TASK_PP(16'h17603,4);
TASK_PP(16'h17604,4);
TASK_PP(16'h17605,4);
TASK_PP(16'h17606,4);
TASK_PP(16'h17607,4);
TASK_PP(16'h17608,4);
TASK_PP(16'h17609,4);
TASK_PP(16'h1760A,4);
TASK_PP(16'h1760B,4);
TASK_PP(16'h1760C,4);
TASK_PP(16'h1760D,4);
TASK_PP(16'h1760E,4);
TASK_PP(16'h1760F,4);
TASK_PP(16'h17610,4);
TASK_PP(16'h17611,4);
TASK_PP(16'h17612,4);
TASK_PP(16'h17613,4);
TASK_PP(16'h17614,4);
TASK_PP(16'h17615,4);
TASK_PP(16'h17616,4);
TASK_PP(16'h17617,4);
TASK_PP(16'h17618,4);
TASK_PP(16'h17619,4);
TASK_PP(16'h1761A,4);
TASK_PP(16'h1761B,4);
TASK_PP(16'h1761C,4);
TASK_PP(16'h1761D,4);
TASK_PP(16'h1761E,4);
TASK_PP(16'h1761F,4);
TASK_PP(16'h17620,4);
TASK_PP(16'h17621,4);
TASK_PP(16'h17622,4);
TASK_PP(16'h17623,4);
TASK_PP(16'h17624,4);
TASK_PP(16'h17625,4);
TASK_PP(16'h17626,4);
TASK_PP(16'h17627,4);
TASK_PP(16'h17628,4);
TASK_PP(16'h17629,4);
TASK_PP(16'h1762A,4);
TASK_PP(16'h1762B,4);
TASK_PP(16'h1762C,4);
TASK_PP(16'h1762D,4);
TASK_PP(16'h1762E,4);
TASK_PP(16'h1762F,4);
TASK_PP(16'h17630,4);
TASK_PP(16'h17631,4);
TASK_PP(16'h17632,4);
TASK_PP(16'h17633,4);
TASK_PP(16'h17634,4);
TASK_PP(16'h17635,4);
TASK_PP(16'h17636,4);
TASK_PP(16'h17637,4);
TASK_PP(16'h17638,4);
TASK_PP(16'h17639,4);
TASK_PP(16'h1763A,4);
TASK_PP(16'h1763B,4);
TASK_PP(16'h1763C,4);
TASK_PP(16'h1763D,4);
TASK_PP(16'h1763E,4);
TASK_PP(16'h1763F,4);
TASK_PP(16'h17640,4);
TASK_PP(16'h17641,4);
TASK_PP(16'h17642,4);
TASK_PP(16'h17643,4);
TASK_PP(16'h17644,4);
TASK_PP(16'h17645,4);
TASK_PP(16'h17646,4);
TASK_PP(16'h17647,4);
TASK_PP(16'h17648,4);
TASK_PP(16'h17649,4);
TASK_PP(16'h1764A,4);
TASK_PP(16'h1764B,4);
TASK_PP(16'h1764C,4);
TASK_PP(16'h1764D,4);
TASK_PP(16'h1764E,4);
TASK_PP(16'h1764F,4);
TASK_PP(16'h17650,4);
TASK_PP(16'h17651,4);
TASK_PP(16'h17652,4);
TASK_PP(16'h17653,4);
TASK_PP(16'h17654,4);
TASK_PP(16'h17655,4);
TASK_PP(16'h17656,4);
TASK_PP(16'h17657,4);
TASK_PP(16'h17658,4);
TASK_PP(16'h17659,4);
TASK_PP(16'h1765A,4);
TASK_PP(16'h1765B,4);
TASK_PP(16'h1765C,4);
TASK_PP(16'h1765D,4);
TASK_PP(16'h1765E,4);
TASK_PP(16'h1765F,4);
TASK_PP(16'h17660,4);
TASK_PP(16'h17661,4);
TASK_PP(16'h17662,4);
TASK_PP(16'h17663,4);
TASK_PP(16'h17664,4);
TASK_PP(16'h17665,4);
TASK_PP(16'h17666,4);
TASK_PP(16'h17667,4);
TASK_PP(16'h17668,4);
TASK_PP(16'h17669,4);
TASK_PP(16'h1766A,4);
TASK_PP(16'h1766B,4);
TASK_PP(16'h1766C,4);
TASK_PP(16'h1766D,4);
TASK_PP(16'h1766E,4);
TASK_PP(16'h1766F,4);
TASK_PP(16'h17670,4);
TASK_PP(16'h17671,4);
TASK_PP(16'h17672,4);
TASK_PP(16'h17673,4);
TASK_PP(16'h17674,4);
TASK_PP(16'h17675,4);
TASK_PP(16'h17676,4);
TASK_PP(16'h17677,4);
TASK_PP(16'h17678,4);
TASK_PP(16'h17679,4);
TASK_PP(16'h1767A,4);
TASK_PP(16'h1767B,4);
TASK_PP(16'h1767C,4);
TASK_PP(16'h1767D,4);
TASK_PP(16'h1767E,4);
TASK_PP(16'h1767F,4);
TASK_PP(16'h17680,4);
TASK_PP(16'h17681,4);
TASK_PP(16'h17682,4);
TASK_PP(16'h17683,4);
TASK_PP(16'h17684,4);
TASK_PP(16'h17685,4);
TASK_PP(16'h17686,4);
TASK_PP(16'h17687,4);
TASK_PP(16'h17688,4);
TASK_PP(16'h17689,4);
TASK_PP(16'h1768A,4);
TASK_PP(16'h1768B,4);
TASK_PP(16'h1768C,4);
TASK_PP(16'h1768D,4);
TASK_PP(16'h1768E,4);
TASK_PP(16'h1768F,4);
TASK_PP(16'h17690,4);
TASK_PP(16'h17691,4);
TASK_PP(16'h17692,4);
TASK_PP(16'h17693,4);
TASK_PP(16'h17694,4);
TASK_PP(16'h17695,4);
TASK_PP(16'h17696,4);
TASK_PP(16'h17697,4);
TASK_PP(16'h17698,4);
TASK_PP(16'h17699,4);
TASK_PP(16'h1769A,4);
TASK_PP(16'h1769B,4);
TASK_PP(16'h1769C,4);
TASK_PP(16'h1769D,4);
TASK_PP(16'h1769E,4);
TASK_PP(16'h1769F,4);
TASK_PP(16'h176A0,4);
TASK_PP(16'h176A1,4);
TASK_PP(16'h176A2,4);
TASK_PP(16'h176A3,4);
TASK_PP(16'h176A4,4);
TASK_PP(16'h176A5,4);
TASK_PP(16'h176A6,4);
TASK_PP(16'h176A7,4);
TASK_PP(16'h176A8,4);
TASK_PP(16'h176A9,4);
TASK_PP(16'h176AA,4);
TASK_PP(16'h176AB,4);
TASK_PP(16'h176AC,4);
TASK_PP(16'h176AD,4);
TASK_PP(16'h176AE,4);
TASK_PP(16'h176AF,4);
TASK_PP(16'h176B0,4);
TASK_PP(16'h176B1,4);
TASK_PP(16'h176B2,4);
TASK_PP(16'h176B3,4);
TASK_PP(16'h176B4,4);
TASK_PP(16'h176B5,4);
TASK_PP(16'h176B6,4);
TASK_PP(16'h176B7,4);
TASK_PP(16'h176B8,4);
TASK_PP(16'h176B9,4);
TASK_PP(16'h176BA,4);
TASK_PP(16'h176BB,4);
TASK_PP(16'h176BC,4);
TASK_PP(16'h176BD,4);
TASK_PP(16'h176BE,4);
TASK_PP(16'h176BF,4);
TASK_PP(16'h176C0,4);
TASK_PP(16'h176C1,4);
TASK_PP(16'h176C2,4);
TASK_PP(16'h176C3,4);
TASK_PP(16'h176C4,4);
TASK_PP(16'h176C5,4);
TASK_PP(16'h176C6,4);
TASK_PP(16'h176C7,4);
TASK_PP(16'h176C8,4);
TASK_PP(16'h176C9,4);
TASK_PP(16'h176CA,4);
TASK_PP(16'h176CB,4);
TASK_PP(16'h176CC,4);
TASK_PP(16'h176CD,4);
TASK_PP(16'h176CE,4);
TASK_PP(16'h176CF,4);
TASK_PP(16'h176D0,4);
TASK_PP(16'h176D1,4);
TASK_PP(16'h176D2,4);
TASK_PP(16'h176D3,4);
TASK_PP(16'h176D4,4);
TASK_PP(16'h176D5,4);
TASK_PP(16'h176D6,4);
TASK_PP(16'h176D7,4);
TASK_PP(16'h176D8,4);
TASK_PP(16'h176D9,4);
TASK_PP(16'h176DA,4);
TASK_PP(16'h176DB,4);
TASK_PP(16'h176DC,4);
TASK_PP(16'h176DD,4);
TASK_PP(16'h176DE,4);
TASK_PP(16'h176DF,4);
TASK_PP(16'h176E0,4);
TASK_PP(16'h176E1,4);
TASK_PP(16'h176E2,4);
TASK_PP(16'h176E3,4);
TASK_PP(16'h176E4,4);
TASK_PP(16'h176E5,4);
TASK_PP(16'h176E6,4);
TASK_PP(16'h176E7,4);
TASK_PP(16'h176E8,4);
TASK_PP(16'h176E9,4);
TASK_PP(16'h176EA,4);
TASK_PP(16'h176EB,4);
TASK_PP(16'h176EC,4);
TASK_PP(16'h176ED,4);
TASK_PP(16'h176EE,4);
TASK_PP(16'h176EF,4);
TASK_PP(16'h176F0,4);
TASK_PP(16'h176F1,4);
TASK_PP(16'h176F2,4);
TASK_PP(16'h176F3,4);
TASK_PP(16'h176F4,4);
TASK_PP(16'h176F5,4);
TASK_PP(16'h176F6,4);
TASK_PP(16'h176F7,4);
TASK_PP(16'h176F8,4);
TASK_PP(16'h176F9,4);
TASK_PP(16'h176FA,4);
TASK_PP(16'h176FB,4);
TASK_PP(16'h176FC,4);
TASK_PP(16'h176FD,4);
TASK_PP(16'h176FE,4);
TASK_PP(16'h176FF,4);
TASK_PP(16'h17700,4);
TASK_PP(16'h17701,4);
TASK_PP(16'h17702,4);
TASK_PP(16'h17703,4);
TASK_PP(16'h17704,4);
TASK_PP(16'h17705,4);
TASK_PP(16'h17706,4);
TASK_PP(16'h17707,4);
TASK_PP(16'h17708,4);
TASK_PP(16'h17709,4);
TASK_PP(16'h1770A,4);
TASK_PP(16'h1770B,4);
TASK_PP(16'h1770C,4);
TASK_PP(16'h1770D,4);
TASK_PP(16'h1770E,4);
TASK_PP(16'h1770F,4);
TASK_PP(16'h17710,4);
TASK_PP(16'h17711,4);
TASK_PP(16'h17712,4);
TASK_PP(16'h17713,4);
TASK_PP(16'h17714,4);
TASK_PP(16'h17715,4);
TASK_PP(16'h17716,4);
TASK_PP(16'h17717,4);
TASK_PP(16'h17718,4);
TASK_PP(16'h17719,4);
TASK_PP(16'h1771A,4);
TASK_PP(16'h1771B,4);
TASK_PP(16'h1771C,4);
TASK_PP(16'h1771D,4);
TASK_PP(16'h1771E,4);
TASK_PP(16'h1771F,4);
TASK_PP(16'h17720,4);
TASK_PP(16'h17721,4);
TASK_PP(16'h17722,4);
TASK_PP(16'h17723,4);
TASK_PP(16'h17724,4);
TASK_PP(16'h17725,4);
TASK_PP(16'h17726,4);
TASK_PP(16'h17727,4);
TASK_PP(16'h17728,4);
TASK_PP(16'h17729,4);
TASK_PP(16'h1772A,4);
TASK_PP(16'h1772B,4);
TASK_PP(16'h1772C,4);
TASK_PP(16'h1772D,4);
TASK_PP(16'h1772E,4);
TASK_PP(16'h1772F,4);
TASK_PP(16'h17730,4);
TASK_PP(16'h17731,4);
TASK_PP(16'h17732,4);
TASK_PP(16'h17733,4);
TASK_PP(16'h17734,4);
TASK_PP(16'h17735,4);
TASK_PP(16'h17736,4);
TASK_PP(16'h17737,4);
TASK_PP(16'h17738,4);
TASK_PP(16'h17739,4);
TASK_PP(16'h1773A,4);
TASK_PP(16'h1773B,4);
TASK_PP(16'h1773C,4);
TASK_PP(16'h1773D,4);
TASK_PP(16'h1773E,4);
TASK_PP(16'h1773F,4);
TASK_PP(16'h17740,4);
TASK_PP(16'h17741,4);
TASK_PP(16'h17742,4);
TASK_PP(16'h17743,4);
TASK_PP(16'h17744,4);
TASK_PP(16'h17745,4);
TASK_PP(16'h17746,4);
TASK_PP(16'h17747,4);
TASK_PP(16'h17748,4);
TASK_PP(16'h17749,4);
TASK_PP(16'h1774A,4);
TASK_PP(16'h1774B,4);
TASK_PP(16'h1774C,4);
TASK_PP(16'h1774D,4);
TASK_PP(16'h1774E,4);
TASK_PP(16'h1774F,4);
TASK_PP(16'h17750,4);
TASK_PP(16'h17751,4);
TASK_PP(16'h17752,4);
TASK_PP(16'h17753,4);
TASK_PP(16'h17754,4);
TASK_PP(16'h17755,4);
TASK_PP(16'h17756,4);
TASK_PP(16'h17757,4);
TASK_PP(16'h17758,4);
TASK_PP(16'h17759,4);
TASK_PP(16'h1775A,4);
TASK_PP(16'h1775B,4);
TASK_PP(16'h1775C,4);
TASK_PP(16'h1775D,4);
TASK_PP(16'h1775E,4);
TASK_PP(16'h1775F,4);
TASK_PP(16'h17760,4);
TASK_PP(16'h17761,4);
TASK_PP(16'h17762,4);
TASK_PP(16'h17763,4);
TASK_PP(16'h17764,4);
TASK_PP(16'h17765,4);
TASK_PP(16'h17766,4);
TASK_PP(16'h17767,4);
TASK_PP(16'h17768,4);
TASK_PP(16'h17769,4);
TASK_PP(16'h1776A,4);
TASK_PP(16'h1776B,4);
TASK_PP(16'h1776C,4);
TASK_PP(16'h1776D,4);
TASK_PP(16'h1776E,4);
TASK_PP(16'h1776F,4);
TASK_PP(16'h17770,4);
TASK_PP(16'h17771,4);
TASK_PP(16'h17772,4);
TASK_PP(16'h17773,4);
TASK_PP(16'h17774,4);
TASK_PP(16'h17775,4);
TASK_PP(16'h17776,4);
TASK_PP(16'h17777,4);
TASK_PP(16'h17778,4);
TASK_PP(16'h17779,4);
TASK_PP(16'h1777A,4);
TASK_PP(16'h1777B,4);
TASK_PP(16'h1777C,4);
TASK_PP(16'h1777D,4);
TASK_PP(16'h1777E,4);
TASK_PP(16'h1777F,4);
TASK_PP(16'h17780,4);
TASK_PP(16'h17781,4);
TASK_PP(16'h17782,4);
TASK_PP(16'h17783,4);
TASK_PP(16'h17784,4);
TASK_PP(16'h17785,4);
TASK_PP(16'h17786,4);
TASK_PP(16'h17787,4);
TASK_PP(16'h17788,4);
TASK_PP(16'h17789,4);
TASK_PP(16'h1778A,4);
TASK_PP(16'h1778B,4);
TASK_PP(16'h1778C,4);
TASK_PP(16'h1778D,4);
TASK_PP(16'h1778E,4);
TASK_PP(16'h1778F,4);
TASK_PP(16'h17790,4);
TASK_PP(16'h17791,4);
TASK_PP(16'h17792,4);
TASK_PP(16'h17793,4);
TASK_PP(16'h17794,4);
TASK_PP(16'h17795,4);
TASK_PP(16'h17796,4);
TASK_PP(16'h17797,4);
TASK_PP(16'h17798,4);
TASK_PP(16'h17799,4);
TASK_PP(16'h1779A,4);
TASK_PP(16'h1779B,4);
TASK_PP(16'h1779C,4);
TASK_PP(16'h1779D,4);
TASK_PP(16'h1779E,4);
TASK_PP(16'h1779F,4);
TASK_PP(16'h177A0,4);
TASK_PP(16'h177A1,4);
TASK_PP(16'h177A2,4);
TASK_PP(16'h177A3,4);
TASK_PP(16'h177A4,4);
TASK_PP(16'h177A5,4);
TASK_PP(16'h177A6,4);
TASK_PP(16'h177A7,4);
TASK_PP(16'h177A8,4);
TASK_PP(16'h177A9,4);
TASK_PP(16'h177AA,4);
TASK_PP(16'h177AB,4);
TASK_PP(16'h177AC,4);
TASK_PP(16'h177AD,4);
TASK_PP(16'h177AE,4);
TASK_PP(16'h177AF,4);
TASK_PP(16'h177B0,4);
TASK_PP(16'h177B1,4);
TASK_PP(16'h177B2,4);
TASK_PP(16'h177B3,4);
TASK_PP(16'h177B4,4);
TASK_PP(16'h177B5,4);
TASK_PP(16'h177B6,4);
TASK_PP(16'h177B7,4);
TASK_PP(16'h177B8,4);
TASK_PP(16'h177B9,4);
TASK_PP(16'h177BA,4);
TASK_PP(16'h177BB,4);
TASK_PP(16'h177BC,4);
TASK_PP(16'h177BD,4);
TASK_PP(16'h177BE,4);
TASK_PP(16'h177BF,4);
TASK_PP(16'h177C0,4);
TASK_PP(16'h177C1,4);
TASK_PP(16'h177C2,4);
TASK_PP(16'h177C3,4);
TASK_PP(16'h177C4,4);
TASK_PP(16'h177C5,4);
TASK_PP(16'h177C6,4);
TASK_PP(16'h177C7,4);
TASK_PP(16'h177C8,4);
TASK_PP(16'h177C9,4);
TASK_PP(16'h177CA,4);
TASK_PP(16'h177CB,4);
TASK_PP(16'h177CC,4);
TASK_PP(16'h177CD,4);
TASK_PP(16'h177CE,4);
TASK_PP(16'h177CF,4);
TASK_PP(16'h177D0,4);
TASK_PP(16'h177D1,4);
TASK_PP(16'h177D2,4);
TASK_PP(16'h177D3,4);
TASK_PP(16'h177D4,4);
TASK_PP(16'h177D5,4);
TASK_PP(16'h177D6,4);
TASK_PP(16'h177D7,4);
TASK_PP(16'h177D8,4);
TASK_PP(16'h177D9,4);
TASK_PP(16'h177DA,4);
TASK_PP(16'h177DB,4);
TASK_PP(16'h177DC,4);
TASK_PP(16'h177DD,4);
TASK_PP(16'h177DE,4);
TASK_PP(16'h177DF,4);
TASK_PP(16'h177E0,4);
TASK_PP(16'h177E1,4);
TASK_PP(16'h177E2,4);
TASK_PP(16'h177E3,4);
TASK_PP(16'h177E4,4);
TASK_PP(16'h177E5,4);
TASK_PP(16'h177E6,4);
TASK_PP(16'h177E7,4);
TASK_PP(16'h177E8,4);
TASK_PP(16'h177E9,4);
TASK_PP(16'h177EA,4);
TASK_PP(16'h177EB,4);
TASK_PP(16'h177EC,4);
TASK_PP(16'h177ED,4);
TASK_PP(16'h177EE,4);
TASK_PP(16'h177EF,4);
TASK_PP(16'h177F0,4);
TASK_PP(16'h177F1,4);
TASK_PP(16'h177F2,4);
TASK_PP(16'h177F3,4);
TASK_PP(16'h177F4,4);
TASK_PP(16'h177F5,4);
TASK_PP(16'h177F6,4);
TASK_PP(16'h177F7,4);
TASK_PP(16'h177F8,4);
TASK_PP(16'h177F9,4);
TASK_PP(16'h177FA,4);
TASK_PP(16'h177FB,4);
TASK_PP(16'h177FC,4);
TASK_PP(16'h177FD,4);
TASK_PP(16'h177FE,4);
TASK_PP(16'h177FF,4);
TASK_PP(16'h17800,4);
TASK_PP(16'h17801,4);
TASK_PP(16'h17802,4);
TASK_PP(16'h17803,4);
TASK_PP(16'h17804,4);
TASK_PP(16'h17805,4);
TASK_PP(16'h17806,4);
TASK_PP(16'h17807,4);
TASK_PP(16'h17808,4);
TASK_PP(16'h17809,4);
TASK_PP(16'h1780A,4);
TASK_PP(16'h1780B,4);
TASK_PP(16'h1780C,4);
TASK_PP(16'h1780D,4);
TASK_PP(16'h1780E,4);
TASK_PP(16'h1780F,4);
TASK_PP(16'h17810,4);
TASK_PP(16'h17811,4);
TASK_PP(16'h17812,4);
TASK_PP(16'h17813,4);
TASK_PP(16'h17814,4);
TASK_PP(16'h17815,4);
TASK_PP(16'h17816,4);
TASK_PP(16'h17817,4);
TASK_PP(16'h17818,4);
TASK_PP(16'h17819,4);
TASK_PP(16'h1781A,4);
TASK_PP(16'h1781B,4);
TASK_PP(16'h1781C,4);
TASK_PP(16'h1781D,4);
TASK_PP(16'h1781E,4);
TASK_PP(16'h1781F,4);
TASK_PP(16'h17820,4);
TASK_PP(16'h17821,4);
TASK_PP(16'h17822,4);
TASK_PP(16'h17823,4);
TASK_PP(16'h17824,4);
TASK_PP(16'h17825,4);
TASK_PP(16'h17826,4);
TASK_PP(16'h17827,4);
TASK_PP(16'h17828,4);
TASK_PP(16'h17829,4);
TASK_PP(16'h1782A,4);
TASK_PP(16'h1782B,4);
TASK_PP(16'h1782C,4);
TASK_PP(16'h1782D,4);
TASK_PP(16'h1782E,4);
TASK_PP(16'h1782F,4);
TASK_PP(16'h17830,4);
TASK_PP(16'h17831,4);
TASK_PP(16'h17832,4);
TASK_PP(16'h17833,4);
TASK_PP(16'h17834,4);
TASK_PP(16'h17835,4);
TASK_PP(16'h17836,4);
TASK_PP(16'h17837,4);
TASK_PP(16'h17838,4);
TASK_PP(16'h17839,4);
TASK_PP(16'h1783A,4);
TASK_PP(16'h1783B,4);
TASK_PP(16'h1783C,4);
TASK_PP(16'h1783D,4);
TASK_PP(16'h1783E,4);
TASK_PP(16'h1783F,4);
TASK_PP(16'h17840,4);
TASK_PP(16'h17841,4);
TASK_PP(16'h17842,4);
TASK_PP(16'h17843,4);
TASK_PP(16'h17844,4);
TASK_PP(16'h17845,4);
TASK_PP(16'h17846,4);
TASK_PP(16'h17847,4);
TASK_PP(16'h17848,4);
TASK_PP(16'h17849,4);
TASK_PP(16'h1784A,4);
TASK_PP(16'h1784B,4);
TASK_PP(16'h1784C,4);
TASK_PP(16'h1784D,4);
TASK_PP(16'h1784E,4);
TASK_PP(16'h1784F,4);
TASK_PP(16'h17850,4);
TASK_PP(16'h17851,4);
TASK_PP(16'h17852,4);
TASK_PP(16'h17853,4);
TASK_PP(16'h17854,4);
TASK_PP(16'h17855,4);
TASK_PP(16'h17856,4);
TASK_PP(16'h17857,4);
TASK_PP(16'h17858,4);
TASK_PP(16'h17859,4);
TASK_PP(16'h1785A,4);
TASK_PP(16'h1785B,4);
TASK_PP(16'h1785C,4);
TASK_PP(16'h1785D,4);
TASK_PP(16'h1785E,4);
TASK_PP(16'h1785F,4);
TASK_PP(16'h17860,4);
TASK_PP(16'h17861,4);
TASK_PP(16'h17862,4);
TASK_PP(16'h17863,4);
TASK_PP(16'h17864,4);
TASK_PP(16'h17865,4);
TASK_PP(16'h17866,4);
TASK_PP(16'h17867,4);
TASK_PP(16'h17868,4);
TASK_PP(16'h17869,4);
TASK_PP(16'h1786A,4);
TASK_PP(16'h1786B,4);
TASK_PP(16'h1786C,4);
TASK_PP(16'h1786D,4);
TASK_PP(16'h1786E,4);
TASK_PP(16'h1786F,4);
TASK_PP(16'h17870,4);
TASK_PP(16'h17871,4);
TASK_PP(16'h17872,4);
TASK_PP(16'h17873,4);
TASK_PP(16'h17874,4);
TASK_PP(16'h17875,4);
TASK_PP(16'h17876,4);
TASK_PP(16'h17877,4);
TASK_PP(16'h17878,4);
TASK_PP(16'h17879,4);
TASK_PP(16'h1787A,4);
TASK_PP(16'h1787B,4);
TASK_PP(16'h1787C,4);
TASK_PP(16'h1787D,4);
TASK_PP(16'h1787E,4);
TASK_PP(16'h1787F,4);
TASK_PP(16'h17880,4);
TASK_PP(16'h17881,4);
TASK_PP(16'h17882,4);
TASK_PP(16'h17883,4);
TASK_PP(16'h17884,4);
TASK_PP(16'h17885,4);
TASK_PP(16'h17886,4);
TASK_PP(16'h17887,4);
TASK_PP(16'h17888,4);
TASK_PP(16'h17889,4);
TASK_PP(16'h1788A,4);
TASK_PP(16'h1788B,4);
TASK_PP(16'h1788C,4);
TASK_PP(16'h1788D,4);
TASK_PP(16'h1788E,4);
TASK_PP(16'h1788F,4);
TASK_PP(16'h17890,4);
TASK_PP(16'h17891,4);
TASK_PP(16'h17892,4);
TASK_PP(16'h17893,4);
TASK_PP(16'h17894,4);
TASK_PP(16'h17895,4);
TASK_PP(16'h17896,4);
TASK_PP(16'h17897,4);
TASK_PP(16'h17898,4);
TASK_PP(16'h17899,4);
TASK_PP(16'h1789A,4);
TASK_PP(16'h1789B,4);
TASK_PP(16'h1789C,4);
TASK_PP(16'h1789D,4);
TASK_PP(16'h1789E,4);
TASK_PP(16'h1789F,4);
TASK_PP(16'h178A0,4);
TASK_PP(16'h178A1,4);
TASK_PP(16'h178A2,4);
TASK_PP(16'h178A3,4);
TASK_PP(16'h178A4,4);
TASK_PP(16'h178A5,4);
TASK_PP(16'h178A6,4);
TASK_PP(16'h178A7,4);
TASK_PP(16'h178A8,4);
TASK_PP(16'h178A9,4);
TASK_PP(16'h178AA,4);
TASK_PP(16'h178AB,4);
TASK_PP(16'h178AC,4);
TASK_PP(16'h178AD,4);
TASK_PP(16'h178AE,4);
TASK_PP(16'h178AF,4);
TASK_PP(16'h178B0,4);
TASK_PP(16'h178B1,4);
TASK_PP(16'h178B2,4);
TASK_PP(16'h178B3,4);
TASK_PP(16'h178B4,4);
TASK_PP(16'h178B5,4);
TASK_PP(16'h178B6,4);
TASK_PP(16'h178B7,4);
TASK_PP(16'h178B8,4);
TASK_PP(16'h178B9,4);
TASK_PP(16'h178BA,4);
TASK_PP(16'h178BB,4);
TASK_PP(16'h178BC,4);
TASK_PP(16'h178BD,4);
TASK_PP(16'h178BE,4);
TASK_PP(16'h178BF,4);
TASK_PP(16'h178C0,4);
TASK_PP(16'h178C1,4);
TASK_PP(16'h178C2,4);
TASK_PP(16'h178C3,4);
TASK_PP(16'h178C4,4);
TASK_PP(16'h178C5,4);
TASK_PP(16'h178C6,4);
TASK_PP(16'h178C7,4);
TASK_PP(16'h178C8,4);
TASK_PP(16'h178C9,4);
TASK_PP(16'h178CA,4);
TASK_PP(16'h178CB,4);
TASK_PP(16'h178CC,4);
TASK_PP(16'h178CD,4);
TASK_PP(16'h178CE,4);
TASK_PP(16'h178CF,4);
TASK_PP(16'h178D0,4);
TASK_PP(16'h178D1,4);
TASK_PP(16'h178D2,4);
TASK_PP(16'h178D3,4);
TASK_PP(16'h178D4,4);
TASK_PP(16'h178D5,4);
TASK_PP(16'h178D6,4);
TASK_PP(16'h178D7,4);
TASK_PP(16'h178D8,4);
TASK_PP(16'h178D9,4);
TASK_PP(16'h178DA,4);
TASK_PP(16'h178DB,4);
TASK_PP(16'h178DC,4);
TASK_PP(16'h178DD,4);
TASK_PP(16'h178DE,4);
TASK_PP(16'h178DF,4);
TASK_PP(16'h178E0,4);
TASK_PP(16'h178E1,4);
TASK_PP(16'h178E2,4);
TASK_PP(16'h178E3,4);
TASK_PP(16'h178E4,4);
TASK_PP(16'h178E5,4);
TASK_PP(16'h178E6,4);
TASK_PP(16'h178E7,4);
TASK_PP(16'h178E8,4);
TASK_PP(16'h178E9,4);
TASK_PP(16'h178EA,4);
TASK_PP(16'h178EB,4);
TASK_PP(16'h178EC,4);
TASK_PP(16'h178ED,4);
TASK_PP(16'h178EE,4);
TASK_PP(16'h178EF,4);
TASK_PP(16'h178F0,4);
TASK_PP(16'h178F1,4);
TASK_PP(16'h178F2,4);
TASK_PP(16'h178F3,4);
TASK_PP(16'h178F4,4);
TASK_PP(16'h178F5,4);
TASK_PP(16'h178F6,4);
TASK_PP(16'h178F7,4);
TASK_PP(16'h178F8,4);
TASK_PP(16'h178F9,4);
TASK_PP(16'h178FA,4);
TASK_PP(16'h178FB,4);
TASK_PP(16'h178FC,4);
TASK_PP(16'h178FD,4);
TASK_PP(16'h178FE,4);
TASK_PP(16'h178FF,4);
TASK_PP(16'h17900,4);
TASK_PP(16'h17901,4);
TASK_PP(16'h17902,4);
TASK_PP(16'h17903,4);
TASK_PP(16'h17904,4);
TASK_PP(16'h17905,4);
TASK_PP(16'h17906,4);
TASK_PP(16'h17907,4);
TASK_PP(16'h17908,4);
TASK_PP(16'h17909,4);
TASK_PP(16'h1790A,4);
TASK_PP(16'h1790B,4);
TASK_PP(16'h1790C,4);
TASK_PP(16'h1790D,4);
TASK_PP(16'h1790E,4);
TASK_PP(16'h1790F,4);
TASK_PP(16'h17910,4);
TASK_PP(16'h17911,4);
TASK_PP(16'h17912,4);
TASK_PP(16'h17913,4);
TASK_PP(16'h17914,4);
TASK_PP(16'h17915,4);
TASK_PP(16'h17916,4);
TASK_PP(16'h17917,4);
TASK_PP(16'h17918,4);
TASK_PP(16'h17919,4);
TASK_PP(16'h1791A,4);
TASK_PP(16'h1791B,4);
TASK_PP(16'h1791C,4);
TASK_PP(16'h1791D,4);
TASK_PP(16'h1791E,4);
TASK_PP(16'h1791F,4);
TASK_PP(16'h17920,4);
TASK_PP(16'h17921,4);
TASK_PP(16'h17922,4);
TASK_PP(16'h17923,4);
TASK_PP(16'h17924,4);
TASK_PP(16'h17925,4);
TASK_PP(16'h17926,4);
TASK_PP(16'h17927,4);
TASK_PP(16'h17928,4);
TASK_PP(16'h17929,4);
TASK_PP(16'h1792A,4);
TASK_PP(16'h1792B,4);
TASK_PP(16'h1792C,4);
TASK_PP(16'h1792D,4);
TASK_PP(16'h1792E,4);
TASK_PP(16'h1792F,4);
TASK_PP(16'h17930,4);
TASK_PP(16'h17931,4);
TASK_PP(16'h17932,4);
TASK_PP(16'h17933,4);
TASK_PP(16'h17934,4);
TASK_PP(16'h17935,4);
TASK_PP(16'h17936,4);
TASK_PP(16'h17937,4);
TASK_PP(16'h17938,4);
TASK_PP(16'h17939,4);
TASK_PP(16'h1793A,4);
TASK_PP(16'h1793B,4);
TASK_PP(16'h1793C,4);
TASK_PP(16'h1793D,4);
TASK_PP(16'h1793E,4);
TASK_PP(16'h1793F,4);
TASK_PP(16'h17940,4);
TASK_PP(16'h17941,4);
TASK_PP(16'h17942,4);
TASK_PP(16'h17943,4);
TASK_PP(16'h17944,4);
TASK_PP(16'h17945,4);
TASK_PP(16'h17946,4);
TASK_PP(16'h17947,4);
TASK_PP(16'h17948,4);
TASK_PP(16'h17949,4);
TASK_PP(16'h1794A,4);
TASK_PP(16'h1794B,4);
TASK_PP(16'h1794C,4);
TASK_PP(16'h1794D,4);
TASK_PP(16'h1794E,4);
TASK_PP(16'h1794F,4);
TASK_PP(16'h17950,4);
TASK_PP(16'h17951,4);
TASK_PP(16'h17952,4);
TASK_PP(16'h17953,4);
TASK_PP(16'h17954,4);
TASK_PP(16'h17955,4);
TASK_PP(16'h17956,4);
TASK_PP(16'h17957,4);
TASK_PP(16'h17958,4);
TASK_PP(16'h17959,4);
TASK_PP(16'h1795A,4);
TASK_PP(16'h1795B,4);
TASK_PP(16'h1795C,4);
TASK_PP(16'h1795D,4);
TASK_PP(16'h1795E,4);
TASK_PP(16'h1795F,4);
TASK_PP(16'h17960,4);
TASK_PP(16'h17961,4);
TASK_PP(16'h17962,4);
TASK_PP(16'h17963,4);
TASK_PP(16'h17964,4);
TASK_PP(16'h17965,4);
TASK_PP(16'h17966,4);
TASK_PP(16'h17967,4);
TASK_PP(16'h17968,4);
TASK_PP(16'h17969,4);
TASK_PP(16'h1796A,4);
TASK_PP(16'h1796B,4);
TASK_PP(16'h1796C,4);
TASK_PP(16'h1796D,4);
TASK_PP(16'h1796E,4);
TASK_PP(16'h1796F,4);
TASK_PP(16'h17970,4);
TASK_PP(16'h17971,4);
TASK_PP(16'h17972,4);
TASK_PP(16'h17973,4);
TASK_PP(16'h17974,4);
TASK_PP(16'h17975,4);
TASK_PP(16'h17976,4);
TASK_PP(16'h17977,4);
TASK_PP(16'h17978,4);
TASK_PP(16'h17979,4);
TASK_PP(16'h1797A,4);
TASK_PP(16'h1797B,4);
TASK_PP(16'h1797C,4);
TASK_PP(16'h1797D,4);
TASK_PP(16'h1797E,4);
TASK_PP(16'h1797F,4);
TASK_PP(16'h17980,4);
TASK_PP(16'h17981,4);
TASK_PP(16'h17982,4);
TASK_PP(16'h17983,4);
TASK_PP(16'h17984,4);
TASK_PP(16'h17985,4);
TASK_PP(16'h17986,4);
TASK_PP(16'h17987,4);
TASK_PP(16'h17988,4);
TASK_PP(16'h17989,4);
TASK_PP(16'h1798A,4);
TASK_PP(16'h1798B,4);
TASK_PP(16'h1798C,4);
TASK_PP(16'h1798D,4);
TASK_PP(16'h1798E,4);
TASK_PP(16'h1798F,4);
TASK_PP(16'h17990,4);
TASK_PP(16'h17991,4);
TASK_PP(16'h17992,4);
TASK_PP(16'h17993,4);
TASK_PP(16'h17994,4);
TASK_PP(16'h17995,4);
TASK_PP(16'h17996,4);
TASK_PP(16'h17997,4);
TASK_PP(16'h17998,4);
TASK_PP(16'h17999,4);
TASK_PP(16'h1799A,4);
TASK_PP(16'h1799B,4);
TASK_PP(16'h1799C,4);
TASK_PP(16'h1799D,4);
TASK_PP(16'h1799E,4);
TASK_PP(16'h1799F,4);
TASK_PP(16'h179A0,4);
TASK_PP(16'h179A1,4);
TASK_PP(16'h179A2,4);
TASK_PP(16'h179A3,4);
TASK_PP(16'h179A4,4);
TASK_PP(16'h179A5,4);
TASK_PP(16'h179A6,4);
TASK_PP(16'h179A7,4);
TASK_PP(16'h179A8,4);
TASK_PP(16'h179A9,4);
TASK_PP(16'h179AA,4);
TASK_PP(16'h179AB,4);
TASK_PP(16'h179AC,4);
TASK_PP(16'h179AD,4);
TASK_PP(16'h179AE,4);
TASK_PP(16'h179AF,4);
TASK_PP(16'h179B0,4);
TASK_PP(16'h179B1,4);
TASK_PP(16'h179B2,4);
TASK_PP(16'h179B3,4);
TASK_PP(16'h179B4,4);
TASK_PP(16'h179B5,4);
TASK_PP(16'h179B6,4);
TASK_PP(16'h179B7,4);
TASK_PP(16'h179B8,4);
TASK_PP(16'h179B9,4);
TASK_PP(16'h179BA,4);
TASK_PP(16'h179BB,4);
TASK_PP(16'h179BC,4);
TASK_PP(16'h179BD,4);
TASK_PP(16'h179BE,4);
TASK_PP(16'h179BF,4);
TASK_PP(16'h179C0,4);
TASK_PP(16'h179C1,4);
TASK_PP(16'h179C2,4);
TASK_PP(16'h179C3,4);
TASK_PP(16'h179C4,4);
TASK_PP(16'h179C5,4);
TASK_PP(16'h179C6,4);
TASK_PP(16'h179C7,4);
TASK_PP(16'h179C8,4);
TASK_PP(16'h179C9,4);
TASK_PP(16'h179CA,4);
TASK_PP(16'h179CB,4);
TASK_PP(16'h179CC,4);
TASK_PP(16'h179CD,4);
TASK_PP(16'h179CE,4);
TASK_PP(16'h179CF,4);
TASK_PP(16'h179D0,4);
TASK_PP(16'h179D1,4);
TASK_PP(16'h179D2,4);
TASK_PP(16'h179D3,4);
TASK_PP(16'h179D4,4);
TASK_PP(16'h179D5,4);
TASK_PP(16'h179D6,4);
TASK_PP(16'h179D7,4);
TASK_PP(16'h179D8,4);
TASK_PP(16'h179D9,4);
TASK_PP(16'h179DA,4);
TASK_PP(16'h179DB,4);
TASK_PP(16'h179DC,4);
TASK_PP(16'h179DD,4);
TASK_PP(16'h179DE,4);
TASK_PP(16'h179DF,4);
TASK_PP(16'h179E0,4);
TASK_PP(16'h179E1,4);
TASK_PP(16'h179E2,4);
TASK_PP(16'h179E3,4);
TASK_PP(16'h179E4,4);
TASK_PP(16'h179E5,4);
TASK_PP(16'h179E6,4);
TASK_PP(16'h179E7,4);
TASK_PP(16'h179E8,4);
TASK_PP(16'h179E9,4);
TASK_PP(16'h179EA,4);
TASK_PP(16'h179EB,4);
TASK_PP(16'h179EC,4);
TASK_PP(16'h179ED,4);
TASK_PP(16'h179EE,4);
TASK_PP(16'h179EF,4);
TASK_PP(16'h179F0,4);
TASK_PP(16'h179F1,4);
TASK_PP(16'h179F2,4);
TASK_PP(16'h179F3,4);
TASK_PP(16'h179F4,4);
TASK_PP(16'h179F5,4);
TASK_PP(16'h179F6,4);
TASK_PP(16'h179F7,4);
TASK_PP(16'h179F8,4);
TASK_PP(16'h179F9,4);
TASK_PP(16'h179FA,4);
TASK_PP(16'h179FB,4);
TASK_PP(16'h179FC,4);
TASK_PP(16'h179FD,4);
TASK_PP(16'h179FE,4);
TASK_PP(16'h179FF,4);
TASK_PP(16'h17A00,4);
TASK_PP(16'h17A01,4);
TASK_PP(16'h17A02,4);
TASK_PP(16'h17A03,4);
TASK_PP(16'h17A04,4);
TASK_PP(16'h17A05,4);
TASK_PP(16'h17A06,4);
TASK_PP(16'h17A07,4);
TASK_PP(16'h17A08,4);
TASK_PP(16'h17A09,4);
TASK_PP(16'h17A0A,4);
TASK_PP(16'h17A0B,4);
TASK_PP(16'h17A0C,4);
TASK_PP(16'h17A0D,4);
TASK_PP(16'h17A0E,4);
TASK_PP(16'h17A0F,4);
TASK_PP(16'h17A10,4);
TASK_PP(16'h17A11,4);
TASK_PP(16'h17A12,4);
TASK_PP(16'h17A13,4);
TASK_PP(16'h17A14,4);
TASK_PP(16'h17A15,4);
TASK_PP(16'h17A16,4);
TASK_PP(16'h17A17,4);
TASK_PP(16'h17A18,4);
TASK_PP(16'h17A19,4);
TASK_PP(16'h17A1A,4);
TASK_PP(16'h17A1B,4);
TASK_PP(16'h17A1C,4);
TASK_PP(16'h17A1D,4);
TASK_PP(16'h17A1E,4);
TASK_PP(16'h17A1F,4);
TASK_PP(16'h17A20,4);
TASK_PP(16'h17A21,4);
TASK_PP(16'h17A22,4);
TASK_PP(16'h17A23,4);
TASK_PP(16'h17A24,4);
TASK_PP(16'h17A25,4);
TASK_PP(16'h17A26,4);
TASK_PP(16'h17A27,4);
TASK_PP(16'h17A28,4);
TASK_PP(16'h17A29,4);
TASK_PP(16'h17A2A,4);
TASK_PP(16'h17A2B,4);
TASK_PP(16'h17A2C,4);
TASK_PP(16'h17A2D,4);
TASK_PP(16'h17A2E,4);
TASK_PP(16'h17A2F,4);
TASK_PP(16'h17A30,4);
TASK_PP(16'h17A31,4);
TASK_PP(16'h17A32,4);
TASK_PP(16'h17A33,4);
TASK_PP(16'h17A34,4);
TASK_PP(16'h17A35,4);
TASK_PP(16'h17A36,4);
TASK_PP(16'h17A37,4);
TASK_PP(16'h17A38,4);
TASK_PP(16'h17A39,4);
TASK_PP(16'h17A3A,4);
TASK_PP(16'h17A3B,4);
TASK_PP(16'h17A3C,4);
TASK_PP(16'h17A3D,4);
TASK_PP(16'h17A3E,4);
TASK_PP(16'h17A3F,4);
TASK_PP(16'h17A40,4);
TASK_PP(16'h17A41,4);
TASK_PP(16'h17A42,4);
TASK_PP(16'h17A43,4);
TASK_PP(16'h17A44,4);
TASK_PP(16'h17A45,4);
TASK_PP(16'h17A46,4);
TASK_PP(16'h17A47,4);
TASK_PP(16'h17A48,4);
TASK_PP(16'h17A49,4);
TASK_PP(16'h17A4A,4);
TASK_PP(16'h17A4B,4);
TASK_PP(16'h17A4C,4);
TASK_PP(16'h17A4D,4);
TASK_PP(16'h17A4E,4);
TASK_PP(16'h17A4F,4);
TASK_PP(16'h17A50,4);
TASK_PP(16'h17A51,4);
TASK_PP(16'h17A52,4);
TASK_PP(16'h17A53,4);
TASK_PP(16'h17A54,4);
TASK_PP(16'h17A55,4);
TASK_PP(16'h17A56,4);
TASK_PP(16'h17A57,4);
TASK_PP(16'h17A58,4);
TASK_PP(16'h17A59,4);
TASK_PP(16'h17A5A,4);
TASK_PP(16'h17A5B,4);
TASK_PP(16'h17A5C,4);
TASK_PP(16'h17A5D,4);
TASK_PP(16'h17A5E,4);
TASK_PP(16'h17A5F,4);
TASK_PP(16'h17A60,4);
TASK_PP(16'h17A61,4);
TASK_PP(16'h17A62,4);
TASK_PP(16'h17A63,4);
TASK_PP(16'h17A64,4);
TASK_PP(16'h17A65,4);
TASK_PP(16'h17A66,4);
TASK_PP(16'h17A67,4);
TASK_PP(16'h17A68,4);
TASK_PP(16'h17A69,4);
TASK_PP(16'h17A6A,4);
TASK_PP(16'h17A6B,4);
TASK_PP(16'h17A6C,4);
TASK_PP(16'h17A6D,4);
TASK_PP(16'h17A6E,4);
TASK_PP(16'h17A6F,4);
TASK_PP(16'h17A70,4);
TASK_PP(16'h17A71,4);
TASK_PP(16'h17A72,4);
TASK_PP(16'h17A73,4);
TASK_PP(16'h17A74,4);
TASK_PP(16'h17A75,4);
TASK_PP(16'h17A76,4);
TASK_PP(16'h17A77,4);
TASK_PP(16'h17A78,4);
TASK_PP(16'h17A79,4);
TASK_PP(16'h17A7A,4);
TASK_PP(16'h17A7B,4);
TASK_PP(16'h17A7C,4);
TASK_PP(16'h17A7D,4);
TASK_PP(16'h17A7E,4);
TASK_PP(16'h17A7F,4);
TASK_PP(16'h17A80,4);
TASK_PP(16'h17A81,4);
TASK_PP(16'h17A82,4);
TASK_PP(16'h17A83,4);
TASK_PP(16'h17A84,4);
TASK_PP(16'h17A85,4);
TASK_PP(16'h17A86,4);
TASK_PP(16'h17A87,4);
TASK_PP(16'h17A88,4);
TASK_PP(16'h17A89,4);
TASK_PP(16'h17A8A,4);
TASK_PP(16'h17A8B,4);
TASK_PP(16'h17A8C,4);
TASK_PP(16'h17A8D,4);
TASK_PP(16'h17A8E,4);
TASK_PP(16'h17A8F,4);
TASK_PP(16'h17A90,4);
TASK_PP(16'h17A91,4);
TASK_PP(16'h17A92,4);
TASK_PP(16'h17A93,4);
TASK_PP(16'h17A94,4);
TASK_PP(16'h17A95,4);
TASK_PP(16'h17A96,4);
TASK_PP(16'h17A97,4);
TASK_PP(16'h17A98,4);
TASK_PP(16'h17A99,4);
TASK_PP(16'h17A9A,4);
TASK_PP(16'h17A9B,4);
TASK_PP(16'h17A9C,4);
TASK_PP(16'h17A9D,4);
TASK_PP(16'h17A9E,4);
TASK_PP(16'h17A9F,4);
TASK_PP(16'h17AA0,4);
TASK_PP(16'h17AA1,4);
TASK_PP(16'h17AA2,4);
TASK_PP(16'h17AA3,4);
TASK_PP(16'h17AA4,4);
TASK_PP(16'h17AA5,4);
TASK_PP(16'h17AA6,4);
TASK_PP(16'h17AA7,4);
TASK_PP(16'h17AA8,4);
TASK_PP(16'h17AA9,4);
TASK_PP(16'h17AAA,4);
TASK_PP(16'h17AAB,4);
TASK_PP(16'h17AAC,4);
TASK_PP(16'h17AAD,4);
TASK_PP(16'h17AAE,4);
TASK_PP(16'h17AAF,4);
TASK_PP(16'h17AB0,4);
TASK_PP(16'h17AB1,4);
TASK_PP(16'h17AB2,4);
TASK_PP(16'h17AB3,4);
TASK_PP(16'h17AB4,4);
TASK_PP(16'h17AB5,4);
TASK_PP(16'h17AB6,4);
TASK_PP(16'h17AB7,4);
TASK_PP(16'h17AB8,4);
TASK_PP(16'h17AB9,4);
TASK_PP(16'h17ABA,4);
TASK_PP(16'h17ABB,4);
TASK_PP(16'h17ABC,4);
TASK_PP(16'h17ABD,4);
TASK_PP(16'h17ABE,4);
TASK_PP(16'h17ABF,4);
TASK_PP(16'h17AC0,4);
TASK_PP(16'h17AC1,4);
TASK_PP(16'h17AC2,4);
TASK_PP(16'h17AC3,4);
TASK_PP(16'h17AC4,4);
TASK_PP(16'h17AC5,4);
TASK_PP(16'h17AC6,4);
TASK_PP(16'h17AC7,4);
TASK_PP(16'h17AC8,4);
TASK_PP(16'h17AC9,4);
TASK_PP(16'h17ACA,4);
TASK_PP(16'h17ACB,4);
TASK_PP(16'h17ACC,4);
TASK_PP(16'h17ACD,4);
TASK_PP(16'h17ACE,4);
TASK_PP(16'h17ACF,4);
TASK_PP(16'h17AD0,4);
TASK_PP(16'h17AD1,4);
TASK_PP(16'h17AD2,4);
TASK_PP(16'h17AD3,4);
TASK_PP(16'h17AD4,4);
TASK_PP(16'h17AD5,4);
TASK_PP(16'h17AD6,4);
TASK_PP(16'h17AD7,4);
TASK_PP(16'h17AD8,4);
TASK_PP(16'h17AD9,4);
TASK_PP(16'h17ADA,4);
TASK_PP(16'h17ADB,4);
TASK_PP(16'h17ADC,4);
TASK_PP(16'h17ADD,4);
TASK_PP(16'h17ADE,4);
TASK_PP(16'h17ADF,4);
TASK_PP(16'h17AE0,4);
TASK_PP(16'h17AE1,4);
TASK_PP(16'h17AE2,4);
TASK_PP(16'h17AE3,4);
TASK_PP(16'h17AE4,4);
TASK_PP(16'h17AE5,4);
TASK_PP(16'h17AE6,4);
TASK_PP(16'h17AE7,4);
TASK_PP(16'h17AE8,4);
TASK_PP(16'h17AE9,4);
TASK_PP(16'h17AEA,4);
TASK_PP(16'h17AEB,4);
TASK_PP(16'h17AEC,4);
TASK_PP(16'h17AED,4);
TASK_PP(16'h17AEE,4);
TASK_PP(16'h17AEF,4);
TASK_PP(16'h17AF0,4);
TASK_PP(16'h17AF1,4);
TASK_PP(16'h17AF2,4);
TASK_PP(16'h17AF3,4);
TASK_PP(16'h17AF4,4);
TASK_PP(16'h17AF5,4);
TASK_PP(16'h17AF6,4);
TASK_PP(16'h17AF7,4);
TASK_PP(16'h17AF8,4);
TASK_PP(16'h17AF9,4);
TASK_PP(16'h17AFA,4);
TASK_PP(16'h17AFB,4);
TASK_PP(16'h17AFC,4);
TASK_PP(16'h17AFD,4);
TASK_PP(16'h17AFE,4);
TASK_PP(16'h17AFF,4);
TASK_PP(16'h17B00,4);
TASK_PP(16'h17B01,4);
TASK_PP(16'h17B02,4);
TASK_PP(16'h17B03,4);
TASK_PP(16'h17B04,4);
TASK_PP(16'h17B05,4);
TASK_PP(16'h17B06,4);
TASK_PP(16'h17B07,4);
TASK_PP(16'h17B08,4);
TASK_PP(16'h17B09,4);
TASK_PP(16'h17B0A,4);
TASK_PP(16'h17B0B,4);
TASK_PP(16'h17B0C,4);
TASK_PP(16'h17B0D,4);
TASK_PP(16'h17B0E,4);
TASK_PP(16'h17B0F,4);
TASK_PP(16'h17B10,4);
TASK_PP(16'h17B11,4);
TASK_PP(16'h17B12,4);
TASK_PP(16'h17B13,4);
TASK_PP(16'h17B14,4);
TASK_PP(16'h17B15,4);
TASK_PP(16'h17B16,4);
TASK_PP(16'h17B17,4);
TASK_PP(16'h17B18,4);
TASK_PP(16'h17B19,4);
TASK_PP(16'h17B1A,4);
TASK_PP(16'h17B1B,4);
TASK_PP(16'h17B1C,4);
TASK_PP(16'h17B1D,4);
TASK_PP(16'h17B1E,4);
TASK_PP(16'h17B1F,4);
TASK_PP(16'h17B20,4);
TASK_PP(16'h17B21,4);
TASK_PP(16'h17B22,4);
TASK_PP(16'h17B23,4);
TASK_PP(16'h17B24,4);
TASK_PP(16'h17B25,4);
TASK_PP(16'h17B26,4);
TASK_PP(16'h17B27,4);
TASK_PP(16'h17B28,4);
TASK_PP(16'h17B29,4);
TASK_PP(16'h17B2A,4);
TASK_PP(16'h17B2B,4);
TASK_PP(16'h17B2C,4);
TASK_PP(16'h17B2D,4);
TASK_PP(16'h17B2E,4);
TASK_PP(16'h17B2F,4);
TASK_PP(16'h17B30,4);
TASK_PP(16'h17B31,4);
TASK_PP(16'h17B32,4);
TASK_PP(16'h17B33,4);
TASK_PP(16'h17B34,4);
TASK_PP(16'h17B35,4);
TASK_PP(16'h17B36,4);
TASK_PP(16'h17B37,4);
TASK_PP(16'h17B38,4);
TASK_PP(16'h17B39,4);
TASK_PP(16'h17B3A,4);
TASK_PP(16'h17B3B,4);
TASK_PP(16'h17B3C,4);
TASK_PP(16'h17B3D,4);
TASK_PP(16'h17B3E,4);
TASK_PP(16'h17B3F,4);
TASK_PP(16'h17B40,4);
TASK_PP(16'h17B41,4);
TASK_PP(16'h17B42,4);
TASK_PP(16'h17B43,4);
TASK_PP(16'h17B44,4);
TASK_PP(16'h17B45,4);
TASK_PP(16'h17B46,4);
TASK_PP(16'h17B47,4);
TASK_PP(16'h17B48,4);
TASK_PP(16'h17B49,4);
TASK_PP(16'h17B4A,4);
TASK_PP(16'h17B4B,4);
TASK_PP(16'h17B4C,4);
TASK_PP(16'h17B4D,4);
TASK_PP(16'h17B4E,4);
TASK_PP(16'h17B4F,4);
TASK_PP(16'h17B50,4);
TASK_PP(16'h17B51,4);
TASK_PP(16'h17B52,4);
TASK_PP(16'h17B53,4);
TASK_PP(16'h17B54,4);
TASK_PP(16'h17B55,4);
TASK_PP(16'h17B56,4);
TASK_PP(16'h17B57,4);
TASK_PP(16'h17B58,4);
TASK_PP(16'h17B59,4);
TASK_PP(16'h17B5A,4);
TASK_PP(16'h17B5B,4);
TASK_PP(16'h17B5C,4);
TASK_PP(16'h17B5D,4);
TASK_PP(16'h17B5E,4);
TASK_PP(16'h17B5F,4);
TASK_PP(16'h17B60,4);
TASK_PP(16'h17B61,4);
TASK_PP(16'h17B62,4);
TASK_PP(16'h17B63,4);
TASK_PP(16'h17B64,4);
TASK_PP(16'h17B65,4);
TASK_PP(16'h17B66,4);
TASK_PP(16'h17B67,4);
TASK_PP(16'h17B68,4);
TASK_PP(16'h17B69,4);
TASK_PP(16'h17B6A,4);
TASK_PP(16'h17B6B,4);
TASK_PP(16'h17B6C,4);
TASK_PP(16'h17B6D,4);
TASK_PP(16'h17B6E,4);
TASK_PP(16'h17B6F,4);
TASK_PP(16'h17B70,4);
TASK_PP(16'h17B71,4);
TASK_PP(16'h17B72,4);
TASK_PP(16'h17B73,4);
TASK_PP(16'h17B74,4);
TASK_PP(16'h17B75,4);
TASK_PP(16'h17B76,4);
TASK_PP(16'h17B77,4);
TASK_PP(16'h17B78,4);
TASK_PP(16'h17B79,4);
TASK_PP(16'h17B7A,4);
TASK_PP(16'h17B7B,4);
TASK_PP(16'h17B7C,4);
TASK_PP(16'h17B7D,4);
TASK_PP(16'h17B7E,4);
TASK_PP(16'h17B7F,4);
TASK_PP(16'h17B80,4);
TASK_PP(16'h17B81,4);
TASK_PP(16'h17B82,4);
TASK_PP(16'h17B83,4);
TASK_PP(16'h17B84,4);
TASK_PP(16'h17B85,4);
TASK_PP(16'h17B86,4);
TASK_PP(16'h17B87,4);
TASK_PP(16'h17B88,4);
TASK_PP(16'h17B89,4);
TASK_PP(16'h17B8A,4);
TASK_PP(16'h17B8B,4);
TASK_PP(16'h17B8C,4);
TASK_PP(16'h17B8D,4);
TASK_PP(16'h17B8E,4);
TASK_PP(16'h17B8F,4);
TASK_PP(16'h17B90,4);
TASK_PP(16'h17B91,4);
TASK_PP(16'h17B92,4);
TASK_PP(16'h17B93,4);
TASK_PP(16'h17B94,4);
TASK_PP(16'h17B95,4);
TASK_PP(16'h17B96,4);
TASK_PP(16'h17B97,4);
TASK_PP(16'h17B98,4);
TASK_PP(16'h17B99,4);
TASK_PP(16'h17B9A,4);
TASK_PP(16'h17B9B,4);
TASK_PP(16'h17B9C,4);
TASK_PP(16'h17B9D,4);
TASK_PP(16'h17B9E,4);
TASK_PP(16'h17B9F,4);
TASK_PP(16'h17BA0,4);
TASK_PP(16'h17BA1,4);
TASK_PP(16'h17BA2,4);
TASK_PP(16'h17BA3,4);
TASK_PP(16'h17BA4,4);
TASK_PP(16'h17BA5,4);
TASK_PP(16'h17BA6,4);
TASK_PP(16'h17BA7,4);
TASK_PP(16'h17BA8,4);
TASK_PP(16'h17BA9,4);
TASK_PP(16'h17BAA,4);
TASK_PP(16'h17BAB,4);
TASK_PP(16'h17BAC,4);
TASK_PP(16'h17BAD,4);
TASK_PP(16'h17BAE,4);
TASK_PP(16'h17BAF,4);
TASK_PP(16'h17BB0,4);
TASK_PP(16'h17BB1,4);
TASK_PP(16'h17BB2,4);
TASK_PP(16'h17BB3,4);
TASK_PP(16'h17BB4,4);
TASK_PP(16'h17BB5,4);
TASK_PP(16'h17BB6,4);
TASK_PP(16'h17BB7,4);
TASK_PP(16'h17BB8,4);
TASK_PP(16'h17BB9,4);
TASK_PP(16'h17BBA,4);
TASK_PP(16'h17BBB,4);
TASK_PP(16'h17BBC,4);
TASK_PP(16'h17BBD,4);
TASK_PP(16'h17BBE,4);
TASK_PP(16'h17BBF,4);
TASK_PP(16'h17BC0,4);
TASK_PP(16'h17BC1,4);
TASK_PP(16'h17BC2,4);
TASK_PP(16'h17BC3,4);
TASK_PP(16'h17BC4,4);
TASK_PP(16'h17BC5,4);
TASK_PP(16'h17BC6,4);
TASK_PP(16'h17BC7,4);
TASK_PP(16'h17BC8,4);
TASK_PP(16'h17BC9,4);
TASK_PP(16'h17BCA,4);
TASK_PP(16'h17BCB,4);
TASK_PP(16'h17BCC,4);
TASK_PP(16'h17BCD,4);
TASK_PP(16'h17BCE,4);
TASK_PP(16'h17BCF,4);
TASK_PP(16'h17BD0,4);
TASK_PP(16'h17BD1,4);
TASK_PP(16'h17BD2,4);
TASK_PP(16'h17BD3,4);
TASK_PP(16'h17BD4,4);
TASK_PP(16'h17BD5,4);
TASK_PP(16'h17BD6,4);
TASK_PP(16'h17BD7,4);
TASK_PP(16'h17BD8,4);
TASK_PP(16'h17BD9,4);
TASK_PP(16'h17BDA,4);
TASK_PP(16'h17BDB,4);
TASK_PP(16'h17BDC,4);
TASK_PP(16'h17BDD,4);
TASK_PP(16'h17BDE,4);
TASK_PP(16'h17BDF,4);
TASK_PP(16'h17BE0,4);
TASK_PP(16'h17BE1,4);
TASK_PP(16'h17BE2,4);
TASK_PP(16'h17BE3,4);
TASK_PP(16'h17BE4,4);
TASK_PP(16'h17BE5,4);
TASK_PP(16'h17BE6,4);
TASK_PP(16'h17BE7,4);
TASK_PP(16'h17BE8,4);
TASK_PP(16'h17BE9,4);
TASK_PP(16'h17BEA,4);
TASK_PP(16'h17BEB,4);
TASK_PP(16'h17BEC,4);
TASK_PP(16'h17BED,4);
TASK_PP(16'h17BEE,4);
TASK_PP(16'h17BEF,4);
TASK_PP(16'h17BF0,4);
TASK_PP(16'h17BF1,4);
TASK_PP(16'h17BF2,4);
TASK_PP(16'h17BF3,4);
TASK_PP(16'h17BF4,4);
TASK_PP(16'h17BF5,4);
TASK_PP(16'h17BF6,4);
TASK_PP(16'h17BF7,4);
TASK_PP(16'h17BF8,4);
TASK_PP(16'h17BF9,4);
TASK_PP(16'h17BFA,4);
TASK_PP(16'h17BFB,4);
TASK_PP(16'h17BFC,4);
TASK_PP(16'h17BFD,4);
TASK_PP(16'h17BFE,4);
TASK_PP(16'h17BFF,4);
TASK_PP(16'h17C00,4);
TASK_PP(16'h17C01,4);
TASK_PP(16'h17C02,4);
TASK_PP(16'h17C03,4);
TASK_PP(16'h17C04,4);
TASK_PP(16'h17C05,4);
TASK_PP(16'h17C06,4);
TASK_PP(16'h17C07,4);
TASK_PP(16'h17C08,4);
TASK_PP(16'h17C09,4);
TASK_PP(16'h17C0A,4);
TASK_PP(16'h17C0B,4);
TASK_PP(16'h17C0C,4);
TASK_PP(16'h17C0D,4);
TASK_PP(16'h17C0E,4);
TASK_PP(16'h17C0F,4);
TASK_PP(16'h17C10,4);
TASK_PP(16'h17C11,4);
TASK_PP(16'h17C12,4);
TASK_PP(16'h17C13,4);
TASK_PP(16'h17C14,4);
TASK_PP(16'h17C15,4);
TASK_PP(16'h17C16,4);
TASK_PP(16'h17C17,4);
TASK_PP(16'h17C18,4);
TASK_PP(16'h17C19,4);
TASK_PP(16'h17C1A,4);
TASK_PP(16'h17C1B,4);
TASK_PP(16'h17C1C,4);
TASK_PP(16'h17C1D,4);
TASK_PP(16'h17C1E,4);
TASK_PP(16'h17C1F,4);
TASK_PP(16'h17C20,4);
TASK_PP(16'h17C21,4);
TASK_PP(16'h17C22,4);
TASK_PP(16'h17C23,4);
TASK_PP(16'h17C24,4);
TASK_PP(16'h17C25,4);
TASK_PP(16'h17C26,4);
TASK_PP(16'h17C27,4);
TASK_PP(16'h17C28,4);
TASK_PP(16'h17C29,4);
TASK_PP(16'h17C2A,4);
TASK_PP(16'h17C2B,4);
TASK_PP(16'h17C2C,4);
TASK_PP(16'h17C2D,4);
TASK_PP(16'h17C2E,4);
TASK_PP(16'h17C2F,4);
TASK_PP(16'h17C30,4);
TASK_PP(16'h17C31,4);
TASK_PP(16'h17C32,4);
TASK_PP(16'h17C33,4);
TASK_PP(16'h17C34,4);
TASK_PP(16'h17C35,4);
TASK_PP(16'h17C36,4);
TASK_PP(16'h17C37,4);
TASK_PP(16'h17C38,4);
TASK_PP(16'h17C39,4);
TASK_PP(16'h17C3A,4);
TASK_PP(16'h17C3B,4);
TASK_PP(16'h17C3C,4);
TASK_PP(16'h17C3D,4);
TASK_PP(16'h17C3E,4);
TASK_PP(16'h17C3F,4);
TASK_PP(16'h17C40,4);
TASK_PP(16'h17C41,4);
TASK_PP(16'h17C42,4);
TASK_PP(16'h17C43,4);
TASK_PP(16'h17C44,4);
TASK_PP(16'h17C45,4);
TASK_PP(16'h17C46,4);
TASK_PP(16'h17C47,4);
TASK_PP(16'h17C48,4);
TASK_PP(16'h17C49,4);
TASK_PP(16'h17C4A,4);
TASK_PP(16'h17C4B,4);
TASK_PP(16'h17C4C,4);
TASK_PP(16'h17C4D,4);
TASK_PP(16'h17C4E,4);
TASK_PP(16'h17C4F,4);
TASK_PP(16'h17C50,4);
TASK_PP(16'h17C51,4);
TASK_PP(16'h17C52,4);
TASK_PP(16'h17C53,4);
TASK_PP(16'h17C54,4);
TASK_PP(16'h17C55,4);
TASK_PP(16'h17C56,4);
TASK_PP(16'h17C57,4);
TASK_PP(16'h17C58,4);
TASK_PP(16'h17C59,4);
TASK_PP(16'h17C5A,4);
TASK_PP(16'h17C5B,4);
TASK_PP(16'h17C5C,4);
TASK_PP(16'h17C5D,4);
TASK_PP(16'h17C5E,4);
TASK_PP(16'h17C5F,4);
TASK_PP(16'h17C60,4);
TASK_PP(16'h17C61,4);
TASK_PP(16'h17C62,4);
TASK_PP(16'h17C63,4);
TASK_PP(16'h17C64,4);
TASK_PP(16'h17C65,4);
TASK_PP(16'h17C66,4);
TASK_PP(16'h17C67,4);
TASK_PP(16'h17C68,4);
TASK_PP(16'h17C69,4);
TASK_PP(16'h17C6A,4);
TASK_PP(16'h17C6B,4);
TASK_PP(16'h17C6C,4);
TASK_PP(16'h17C6D,4);
TASK_PP(16'h17C6E,4);
TASK_PP(16'h17C6F,4);
TASK_PP(16'h17C70,4);
TASK_PP(16'h17C71,4);
TASK_PP(16'h17C72,4);
TASK_PP(16'h17C73,4);
TASK_PP(16'h17C74,4);
TASK_PP(16'h17C75,4);
TASK_PP(16'h17C76,4);
TASK_PP(16'h17C77,4);
TASK_PP(16'h17C78,4);
TASK_PP(16'h17C79,4);
TASK_PP(16'h17C7A,4);
TASK_PP(16'h17C7B,4);
TASK_PP(16'h17C7C,4);
TASK_PP(16'h17C7D,4);
TASK_PP(16'h17C7E,4);
TASK_PP(16'h17C7F,4);
TASK_PP(16'h17C80,4);
TASK_PP(16'h17C81,4);
TASK_PP(16'h17C82,4);
TASK_PP(16'h17C83,4);
TASK_PP(16'h17C84,4);
TASK_PP(16'h17C85,4);
TASK_PP(16'h17C86,4);
TASK_PP(16'h17C87,4);
TASK_PP(16'h17C88,4);
TASK_PP(16'h17C89,4);
TASK_PP(16'h17C8A,4);
TASK_PP(16'h17C8B,4);
TASK_PP(16'h17C8C,4);
TASK_PP(16'h17C8D,4);
TASK_PP(16'h17C8E,4);
TASK_PP(16'h17C8F,4);
TASK_PP(16'h17C90,4);
TASK_PP(16'h17C91,4);
TASK_PP(16'h17C92,4);
TASK_PP(16'h17C93,4);
TASK_PP(16'h17C94,4);
TASK_PP(16'h17C95,4);
TASK_PP(16'h17C96,4);
TASK_PP(16'h17C97,4);
TASK_PP(16'h17C98,4);
TASK_PP(16'h17C99,4);
TASK_PP(16'h17C9A,4);
TASK_PP(16'h17C9B,4);
TASK_PP(16'h17C9C,4);
TASK_PP(16'h17C9D,4);
TASK_PP(16'h17C9E,4);
TASK_PP(16'h17C9F,4);
TASK_PP(16'h17CA0,4);
TASK_PP(16'h17CA1,4);
TASK_PP(16'h17CA2,4);
TASK_PP(16'h17CA3,4);
TASK_PP(16'h17CA4,4);
TASK_PP(16'h17CA5,4);
TASK_PP(16'h17CA6,4);
TASK_PP(16'h17CA7,4);
TASK_PP(16'h17CA8,4);
TASK_PP(16'h17CA9,4);
TASK_PP(16'h17CAA,4);
TASK_PP(16'h17CAB,4);
TASK_PP(16'h17CAC,4);
TASK_PP(16'h17CAD,4);
TASK_PP(16'h17CAE,4);
TASK_PP(16'h17CAF,4);
TASK_PP(16'h17CB0,4);
TASK_PP(16'h17CB1,4);
TASK_PP(16'h17CB2,4);
TASK_PP(16'h17CB3,4);
TASK_PP(16'h17CB4,4);
TASK_PP(16'h17CB5,4);
TASK_PP(16'h17CB6,4);
TASK_PP(16'h17CB7,4);
TASK_PP(16'h17CB8,4);
TASK_PP(16'h17CB9,4);
TASK_PP(16'h17CBA,4);
TASK_PP(16'h17CBB,4);
TASK_PP(16'h17CBC,4);
TASK_PP(16'h17CBD,4);
TASK_PP(16'h17CBE,4);
TASK_PP(16'h17CBF,4);
TASK_PP(16'h17CC0,4);
TASK_PP(16'h17CC1,4);
TASK_PP(16'h17CC2,4);
TASK_PP(16'h17CC3,4);
TASK_PP(16'h17CC4,4);
TASK_PP(16'h17CC5,4);
TASK_PP(16'h17CC6,4);
TASK_PP(16'h17CC7,4);
TASK_PP(16'h17CC8,4);
TASK_PP(16'h17CC9,4);
TASK_PP(16'h17CCA,4);
TASK_PP(16'h17CCB,4);
TASK_PP(16'h17CCC,4);
TASK_PP(16'h17CCD,4);
TASK_PP(16'h17CCE,4);
TASK_PP(16'h17CCF,4);
TASK_PP(16'h17CD0,4);
TASK_PP(16'h17CD1,4);
TASK_PP(16'h17CD2,4);
TASK_PP(16'h17CD3,4);
TASK_PP(16'h17CD4,4);
TASK_PP(16'h17CD5,4);
TASK_PP(16'h17CD6,4);
TASK_PP(16'h17CD7,4);
TASK_PP(16'h17CD8,4);
TASK_PP(16'h17CD9,4);
TASK_PP(16'h17CDA,4);
TASK_PP(16'h17CDB,4);
TASK_PP(16'h17CDC,4);
TASK_PP(16'h17CDD,4);
TASK_PP(16'h17CDE,4);
TASK_PP(16'h17CDF,4);
TASK_PP(16'h17CE0,4);
TASK_PP(16'h17CE1,4);
TASK_PP(16'h17CE2,4);
TASK_PP(16'h17CE3,4);
TASK_PP(16'h17CE4,4);
TASK_PP(16'h17CE5,4);
TASK_PP(16'h17CE6,4);
TASK_PP(16'h17CE7,4);
TASK_PP(16'h17CE8,4);
TASK_PP(16'h17CE9,4);
TASK_PP(16'h17CEA,4);
TASK_PP(16'h17CEB,4);
TASK_PP(16'h17CEC,4);
TASK_PP(16'h17CED,4);
TASK_PP(16'h17CEE,4);
TASK_PP(16'h17CEF,4);
TASK_PP(16'h17CF0,4);
TASK_PP(16'h17CF1,4);
TASK_PP(16'h17CF2,4);
TASK_PP(16'h17CF3,4);
TASK_PP(16'h17CF4,4);
TASK_PP(16'h17CF5,4);
TASK_PP(16'h17CF6,4);
TASK_PP(16'h17CF7,4);
TASK_PP(16'h17CF8,4);
TASK_PP(16'h17CF9,4);
TASK_PP(16'h17CFA,4);
TASK_PP(16'h17CFB,4);
TASK_PP(16'h17CFC,4);
TASK_PP(16'h17CFD,4);
TASK_PP(16'h17CFE,4);
TASK_PP(16'h17CFF,4);
TASK_PP(16'h17D00,4);
TASK_PP(16'h17D01,4);
TASK_PP(16'h17D02,4);
TASK_PP(16'h17D03,4);
TASK_PP(16'h17D04,4);
TASK_PP(16'h17D05,4);
TASK_PP(16'h17D06,4);
TASK_PP(16'h17D07,4);
TASK_PP(16'h17D08,4);
TASK_PP(16'h17D09,4);
TASK_PP(16'h17D0A,4);
TASK_PP(16'h17D0B,4);
TASK_PP(16'h17D0C,4);
TASK_PP(16'h17D0D,4);
TASK_PP(16'h17D0E,4);
TASK_PP(16'h17D0F,4);
TASK_PP(16'h17D10,4);
TASK_PP(16'h17D11,4);
TASK_PP(16'h17D12,4);
TASK_PP(16'h17D13,4);
TASK_PP(16'h17D14,4);
TASK_PP(16'h17D15,4);
TASK_PP(16'h17D16,4);
TASK_PP(16'h17D17,4);
TASK_PP(16'h17D18,4);
TASK_PP(16'h17D19,4);
TASK_PP(16'h17D1A,4);
TASK_PP(16'h17D1B,4);
TASK_PP(16'h17D1C,4);
TASK_PP(16'h17D1D,4);
TASK_PP(16'h17D1E,4);
TASK_PP(16'h17D1F,4);
TASK_PP(16'h17D20,4);
TASK_PP(16'h17D21,4);
TASK_PP(16'h17D22,4);
TASK_PP(16'h17D23,4);
TASK_PP(16'h17D24,4);
TASK_PP(16'h17D25,4);
TASK_PP(16'h17D26,4);
TASK_PP(16'h17D27,4);
TASK_PP(16'h17D28,4);
TASK_PP(16'h17D29,4);
TASK_PP(16'h17D2A,4);
TASK_PP(16'h17D2B,4);
TASK_PP(16'h17D2C,4);
TASK_PP(16'h17D2D,4);
TASK_PP(16'h17D2E,4);
TASK_PP(16'h17D2F,4);
TASK_PP(16'h17D30,4);
TASK_PP(16'h17D31,4);
TASK_PP(16'h17D32,4);
TASK_PP(16'h17D33,4);
TASK_PP(16'h17D34,4);
TASK_PP(16'h17D35,4);
TASK_PP(16'h17D36,4);
TASK_PP(16'h17D37,4);
TASK_PP(16'h17D38,4);
TASK_PP(16'h17D39,4);
TASK_PP(16'h17D3A,4);
TASK_PP(16'h17D3B,4);
TASK_PP(16'h17D3C,4);
TASK_PP(16'h17D3D,4);
TASK_PP(16'h17D3E,4);
TASK_PP(16'h17D3F,4);
TASK_PP(16'h17D40,4);
TASK_PP(16'h17D41,4);
TASK_PP(16'h17D42,4);
TASK_PP(16'h17D43,4);
TASK_PP(16'h17D44,4);
TASK_PP(16'h17D45,4);
TASK_PP(16'h17D46,4);
TASK_PP(16'h17D47,4);
TASK_PP(16'h17D48,4);
TASK_PP(16'h17D49,4);
TASK_PP(16'h17D4A,4);
TASK_PP(16'h17D4B,4);
TASK_PP(16'h17D4C,4);
TASK_PP(16'h17D4D,4);
TASK_PP(16'h17D4E,4);
TASK_PP(16'h17D4F,4);
TASK_PP(16'h17D50,4);
TASK_PP(16'h17D51,4);
TASK_PP(16'h17D52,4);
TASK_PP(16'h17D53,4);
TASK_PP(16'h17D54,4);
TASK_PP(16'h17D55,4);
TASK_PP(16'h17D56,4);
TASK_PP(16'h17D57,4);
TASK_PP(16'h17D58,4);
TASK_PP(16'h17D59,4);
TASK_PP(16'h17D5A,4);
TASK_PP(16'h17D5B,4);
TASK_PP(16'h17D5C,4);
TASK_PP(16'h17D5D,4);
TASK_PP(16'h17D5E,4);
TASK_PP(16'h17D5F,4);
TASK_PP(16'h17D60,4);
TASK_PP(16'h17D61,4);
TASK_PP(16'h17D62,4);
TASK_PP(16'h17D63,4);
TASK_PP(16'h17D64,4);
TASK_PP(16'h17D65,4);
TASK_PP(16'h17D66,4);
TASK_PP(16'h17D67,4);
TASK_PP(16'h17D68,4);
TASK_PP(16'h17D69,4);
TASK_PP(16'h17D6A,4);
TASK_PP(16'h17D6B,4);
TASK_PP(16'h17D6C,4);
TASK_PP(16'h17D6D,4);
TASK_PP(16'h17D6E,4);
TASK_PP(16'h17D6F,4);
TASK_PP(16'h17D70,4);
TASK_PP(16'h17D71,4);
TASK_PP(16'h17D72,4);
TASK_PP(16'h17D73,4);
TASK_PP(16'h17D74,4);
TASK_PP(16'h17D75,4);
TASK_PP(16'h17D76,4);
TASK_PP(16'h17D77,4);
TASK_PP(16'h17D78,4);
TASK_PP(16'h17D79,4);
TASK_PP(16'h17D7A,4);
TASK_PP(16'h17D7B,4);
TASK_PP(16'h17D7C,4);
TASK_PP(16'h17D7D,4);
TASK_PP(16'h17D7E,4);
TASK_PP(16'h17D7F,4);
TASK_PP(16'h17D80,4);
TASK_PP(16'h17D81,4);
TASK_PP(16'h17D82,4);
TASK_PP(16'h17D83,4);
TASK_PP(16'h17D84,4);
TASK_PP(16'h17D85,4);
TASK_PP(16'h17D86,4);
TASK_PP(16'h17D87,4);
TASK_PP(16'h17D88,4);
TASK_PP(16'h17D89,4);
TASK_PP(16'h17D8A,4);
TASK_PP(16'h17D8B,4);
TASK_PP(16'h17D8C,4);
TASK_PP(16'h17D8D,4);
TASK_PP(16'h17D8E,4);
TASK_PP(16'h17D8F,4);
TASK_PP(16'h17D90,4);
TASK_PP(16'h17D91,4);
TASK_PP(16'h17D92,4);
TASK_PP(16'h17D93,4);
TASK_PP(16'h17D94,4);
TASK_PP(16'h17D95,4);
TASK_PP(16'h17D96,4);
TASK_PP(16'h17D97,4);
TASK_PP(16'h17D98,4);
TASK_PP(16'h17D99,4);
TASK_PP(16'h17D9A,4);
TASK_PP(16'h17D9B,4);
TASK_PP(16'h17D9C,4);
TASK_PP(16'h17D9D,4);
TASK_PP(16'h17D9E,4);
TASK_PP(16'h17D9F,4);
TASK_PP(16'h17DA0,4);
TASK_PP(16'h17DA1,4);
TASK_PP(16'h17DA2,4);
TASK_PP(16'h17DA3,4);
TASK_PP(16'h17DA4,4);
TASK_PP(16'h17DA5,4);
TASK_PP(16'h17DA6,4);
TASK_PP(16'h17DA7,4);
TASK_PP(16'h17DA8,4);
TASK_PP(16'h17DA9,4);
TASK_PP(16'h17DAA,4);
TASK_PP(16'h17DAB,4);
TASK_PP(16'h17DAC,4);
TASK_PP(16'h17DAD,4);
TASK_PP(16'h17DAE,4);
TASK_PP(16'h17DAF,4);
TASK_PP(16'h17DB0,4);
TASK_PP(16'h17DB1,4);
TASK_PP(16'h17DB2,4);
TASK_PP(16'h17DB3,4);
TASK_PP(16'h17DB4,4);
TASK_PP(16'h17DB5,4);
TASK_PP(16'h17DB6,4);
TASK_PP(16'h17DB7,4);
TASK_PP(16'h17DB8,4);
TASK_PP(16'h17DB9,4);
TASK_PP(16'h17DBA,4);
TASK_PP(16'h17DBB,4);
TASK_PP(16'h17DBC,4);
TASK_PP(16'h17DBD,4);
TASK_PP(16'h17DBE,4);
TASK_PP(16'h17DBF,4);
TASK_PP(16'h17DC0,4);
TASK_PP(16'h17DC1,4);
TASK_PP(16'h17DC2,4);
TASK_PP(16'h17DC3,4);
TASK_PP(16'h17DC4,4);
TASK_PP(16'h17DC5,4);
TASK_PP(16'h17DC6,4);
TASK_PP(16'h17DC7,4);
TASK_PP(16'h17DC8,4);
TASK_PP(16'h17DC9,4);
TASK_PP(16'h17DCA,4);
TASK_PP(16'h17DCB,4);
TASK_PP(16'h17DCC,4);
TASK_PP(16'h17DCD,4);
TASK_PP(16'h17DCE,4);
TASK_PP(16'h17DCF,4);
TASK_PP(16'h17DD0,4);
TASK_PP(16'h17DD1,4);
TASK_PP(16'h17DD2,4);
TASK_PP(16'h17DD3,4);
TASK_PP(16'h17DD4,4);
TASK_PP(16'h17DD5,4);
TASK_PP(16'h17DD6,4);
TASK_PP(16'h17DD7,4);
TASK_PP(16'h17DD8,4);
TASK_PP(16'h17DD9,4);
TASK_PP(16'h17DDA,4);
TASK_PP(16'h17DDB,4);
TASK_PP(16'h17DDC,4);
TASK_PP(16'h17DDD,4);
TASK_PP(16'h17DDE,4);
TASK_PP(16'h17DDF,4);
TASK_PP(16'h17DE0,4);
TASK_PP(16'h17DE1,4);
TASK_PP(16'h17DE2,4);
TASK_PP(16'h17DE3,4);
TASK_PP(16'h17DE4,4);
TASK_PP(16'h17DE5,4);
TASK_PP(16'h17DE6,4);
TASK_PP(16'h17DE7,4);
TASK_PP(16'h17DE8,4);
TASK_PP(16'h17DE9,4);
TASK_PP(16'h17DEA,4);
TASK_PP(16'h17DEB,4);
TASK_PP(16'h17DEC,4);
TASK_PP(16'h17DED,4);
TASK_PP(16'h17DEE,4);
TASK_PP(16'h17DEF,4);
TASK_PP(16'h17DF0,4);
TASK_PP(16'h17DF1,4);
TASK_PP(16'h17DF2,4);
TASK_PP(16'h17DF3,4);
TASK_PP(16'h17DF4,4);
TASK_PP(16'h17DF5,4);
TASK_PP(16'h17DF6,4);
TASK_PP(16'h17DF7,4);
TASK_PP(16'h17DF8,4);
TASK_PP(16'h17DF9,4);
TASK_PP(16'h17DFA,4);
TASK_PP(16'h17DFB,4);
TASK_PP(16'h17DFC,4);
TASK_PP(16'h17DFD,4);
TASK_PP(16'h17DFE,4);
TASK_PP(16'h17DFF,4);
TASK_PP(16'h17E00,4);
TASK_PP(16'h17E01,4);
TASK_PP(16'h17E02,4);
TASK_PP(16'h17E03,4);
TASK_PP(16'h17E04,4);
TASK_PP(16'h17E05,4);
TASK_PP(16'h17E06,4);
TASK_PP(16'h17E07,4);
TASK_PP(16'h17E08,4);
TASK_PP(16'h17E09,4);
TASK_PP(16'h17E0A,4);
TASK_PP(16'h17E0B,4);
TASK_PP(16'h17E0C,4);
TASK_PP(16'h17E0D,4);
TASK_PP(16'h17E0E,4);
TASK_PP(16'h17E0F,4);
TASK_PP(16'h17E10,4);
TASK_PP(16'h17E11,4);
TASK_PP(16'h17E12,4);
TASK_PP(16'h17E13,4);
TASK_PP(16'h17E14,4);
TASK_PP(16'h17E15,4);
TASK_PP(16'h17E16,4);
TASK_PP(16'h17E17,4);
TASK_PP(16'h17E18,4);
TASK_PP(16'h17E19,4);
TASK_PP(16'h17E1A,4);
TASK_PP(16'h17E1B,4);
TASK_PP(16'h17E1C,4);
TASK_PP(16'h17E1D,4);
TASK_PP(16'h17E1E,4);
TASK_PP(16'h17E1F,4);
TASK_PP(16'h17E20,4);
TASK_PP(16'h17E21,4);
TASK_PP(16'h17E22,4);
TASK_PP(16'h17E23,4);
TASK_PP(16'h17E24,4);
TASK_PP(16'h17E25,4);
TASK_PP(16'h17E26,4);
TASK_PP(16'h17E27,4);
TASK_PP(16'h17E28,4);
TASK_PP(16'h17E29,4);
TASK_PP(16'h17E2A,4);
TASK_PP(16'h17E2B,4);
TASK_PP(16'h17E2C,4);
TASK_PP(16'h17E2D,4);
TASK_PP(16'h17E2E,4);
TASK_PP(16'h17E2F,4);
TASK_PP(16'h17E30,4);
TASK_PP(16'h17E31,4);
TASK_PP(16'h17E32,4);
TASK_PP(16'h17E33,4);
TASK_PP(16'h17E34,4);
TASK_PP(16'h17E35,4);
TASK_PP(16'h17E36,4);
TASK_PP(16'h17E37,4);
TASK_PP(16'h17E38,4);
TASK_PP(16'h17E39,4);
TASK_PP(16'h17E3A,4);
TASK_PP(16'h17E3B,4);
TASK_PP(16'h17E3C,4);
TASK_PP(16'h17E3D,4);
TASK_PP(16'h17E3E,4);
TASK_PP(16'h17E3F,4);
TASK_PP(16'h17E40,4);
TASK_PP(16'h17E41,4);
TASK_PP(16'h17E42,4);
TASK_PP(16'h17E43,4);
TASK_PP(16'h17E44,4);
TASK_PP(16'h17E45,4);
TASK_PP(16'h17E46,4);
TASK_PP(16'h17E47,4);
TASK_PP(16'h17E48,4);
TASK_PP(16'h17E49,4);
TASK_PP(16'h17E4A,4);
TASK_PP(16'h17E4B,4);
TASK_PP(16'h17E4C,4);
TASK_PP(16'h17E4D,4);
TASK_PP(16'h17E4E,4);
TASK_PP(16'h17E4F,4);
TASK_PP(16'h17E50,4);
TASK_PP(16'h17E51,4);
TASK_PP(16'h17E52,4);
TASK_PP(16'h17E53,4);
TASK_PP(16'h17E54,4);
TASK_PP(16'h17E55,4);
TASK_PP(16'h17E56,4);
TASK_PP(16'h17E57,4);
TASK_PP(16'h17E58,4);
TASK_PP(16'h17E59,4);
TASK_PP(16'h17E5A,4);
TASK_PP(16'h17E5B,4);
TASK_PP(16'h17E5C,4);
TASK_PP(16'h17E5D,4);
TASK_PP(16'h17E5E,4);
TASK_PP(16'h17E5F,4);
TASK_PP(16'h17E60,4);
TASK_PP(16'h17E61,4);
TASK_PP(16'h17E62,4);
TASK_PP(16'h17E63,4);
TASK_PP(16'h17E64,4);
TASK_PP(16'h17E65,4);
TASK_PP(16'h17E66,4);
TASK_PP(16'h17E67,4);
TASK_PP(16'h17E68,4);
TASK_PP(16'h17E69,4);
TASK_PP(16'h17E6A,4);
TASK_PP(16'h17E6B,4);
TASK_PP(16'h17E6C,4);
TASK_PP(16'h17E6D,4);
TASK_PP(16'h17E6E,4);
TASK_PP(16'h17E6F,4);
TASK_PP(16'h17E70,4);
TASK_PP(16'h17E71,4);
TASK_PP(16'h17E72,4);
TASK_PP(16'h17E73,4);
TASK_PP(16'h17E74,4);
TASK_PP(16'h17E75,4);
TASK_PP(16'h17E76,4);
TASK_PP(16'h17E77,4);
TASK_PP(16'h17E78,4);
TASK_PP(16'h17E79,4);
TASK_PP(16'h17E7A,4);
TASK_PP(16'h17E7B,4);
TASK_PP(16'h17E7C,4);
TASK_PP(16'h17E7D,4);
TASK_PP(16'h17E7E,4);
TASK_PP(16'h17E7F,4);
TASK_PP(16'h17E80,4);
TASK_PP(16'h17E81,4);
TASK_PP(16'h17E82,4);
TASK_PP(16'h17E83,4);
TASK_PP(16'h17E84,4);
TASK_PP(16'h17E85,4);
TASK_PP(16'h17E86,4);
TASK_PP(16'h17E87,4);
TASK_PP(16'h17E88,4);
TASK_PP(16'h17E89,4);
TASK_PP(16'h17E8A,4);
TASK_PP(16'h17E8B,4);
TASK_PP(16'h17E8C,4);
TASK_PP(16'h17E8D,4);
TASK_PP(16'h17E8E,4);
TASK_PP(16'h17E8F,4);
TASK_PP(16'h17E90,4);
TASK_PP(16'h17E91,4);
TASK_PP(16'h17E92,4);
TASK_PP(16'h17E93,4);
TASK_PP(16'h17E94,4);
TASK_PP(16'h17E95,4);
TASK_PP(16'h17E96,4);
TASK_PP(16'h17E97,4);
TASK_PP(16'h17E98,4);
TASK_PP(16'h17E99,4);
TASK_PP(16'h17E9A,4);
TASK_PP(16'h17E9B,4);
TASK_PP(16'h17E9C,4);
TASK_PP(16'h17E9D,4);
TASK_PP(16'h17E9E,4);
TASK_PP(16'h17E9F,4);
TASK_PP(16'h17EA0,4);
TASK_PP(16'h17EA1,4);
TASK_PP(16'h17EA2,4);
TASK_PP(16'h17EA3,4);
TASK_PP(16'h17EA4,4);
TASK_PP(16'h17EA5,4);
TASK_PP(16'h17EA6,4);
TASK_PP(16'h17EA7,4);
TASK_PP(16'h17EA8,4);
TASK_PP(16'h17EA9,4);
TASK_PP(16'h17EAA,4);
TASK_PP(16'h17EAB,4);
TASK_PP(16'h17EAC,4);
TASK_PP(16'h17EAD,4);
TASK_PP(16'h17EAE,4);
TASK_PP(16'h17EAF,4);
TASK_PP(16'h17EB0,4);
TASK_PP(16'h17EB1,4);
TASK_PP(16'h17EB2,4);
TASK_PP(16'h17EB3,4);
TASK_PP(16'h17EB4,4);
TASK_PP(16'h17EB5,4);
TASK_PP(16'h17EB6,4);
TASK_PP(16'h17EB7,4);
TASK_PP(16'h17EB8,4);
TASK_PP(16'h17EB9,4);
TASK_PP(16'h17EBA,4);
TASK_PP(16'h17EBB,4);
TASK_PP(16'h17EBC,4);
TASK_PP(16'h17EBD,4);
TASK_PP(16'h17EBE,4);
TASK_PP(16'h17EBF,4);
TASK_PP(16'h17EC0,4);
TASK_PP(16'h17EC1,4);
TASK_PP(16'h17EC2,4);
TASK_PP(16'h17EC3,4);
TASK_PP(16'h17EC4,4);
TASK_PP(16'h17EC5,4);
TASK_PP(16'h17EC6,4);
TASK_PP(16'h17EC7,4);
TASK_PP(16'h17EC8,4);
TASK_PP(16'h17EC9,4);
TASK_PP(16'h17ECA,4);
TASK_PP(16'h17ECB,4);
TASK_PP(16'h17ECC,4);
TASK_PP(16'h17ECD,4);
TASK_PP(16'h17ECE,4);
TASK_PP(16'h17ECF,4);
TASK_PP(16'h17ED0,4);
TASK_PP(16'h17ED1,4);
TASK_PP(16'h17ED2,4);
TASK_PP(16'h17ED3,4);
TASK_PP(16'h17ED4,4);
TASK_PP(16'h17ED5,4);
TASK_PP(16'h17ED6,4);
TASK_PP(16'h17ED7,4);
TASK_PP(16'h17ED8,4);
TASK_PP(16'h17ED9,4);
TASK_PP(16'h17EDA,4);
TASK_PP(16'h17EDB,4);
TASK_PP(16'h17EDC,4);
TASK_PP(16'h17EDD,4);
TASK_PP(16'h17EDE,4);
TASK_PP(16'h17EDF,4);
TASK_PP(16'h17EE0,4);
TASK_PP(16'h17EE1,4);
TASK_PP(16'h17EE2,4);
TASK_PP(16'h17EE3,4);
TASK_PP(16'h17EE4,4);
TASK_PP(16'h17EE5,4);
TASK_PP(16'h17EE6,4);
TASK_PP(16'h17EE7,4);
TASK_PP(16'h17EE8,4);
TASK_PP(16'h17EE9,4);
TASK_PP(16'h17EEA,4);
TASK_PP(16'h17EEB,4);
TASK_PP(16'h17EEC,4);
TASK_PP(16'h17EED,4);
TASK_PP(16'h17EEE,4);
TASK_PP(16'h17EEF,4);
TASK_PP(16'h17EF0,4);
TASK_PP(16'h17EF1,4);
TASK_PP(16'h17EF2,4);
TASK_PP(16'h17EF3,4);
TASK_PP(16'h17EF4,4);
TASK_PP(16'h17EF5,4);
TASK_PP(16'h17EF6,4);
TASK_PP(16'h17EF7,4);
TASK_PP(16'h17EF8,4);
TASK_PP(16'h17EF9,4);
TASK_PP(16'h17EFA,4);
TASK_PP(16'h17EFB,4);
TASK_PP(16'h17EFC,4);
TASK_PP(16'h17EFD,4);
TASK_PP(16'h17EFE,4);
TASK_PP(16'h17EFF,4);
TASK_PP(16'h17F00,4);
TASK_PP(16'h17F01,4);
TASK_PP(16'h17F02,4);
TASK_PP(16'h17F03,4);
TASK_PP(16'h17F04,4);
TASK_PP(16'h17F05,4);
TASK_PP(16'h17F06,4);
TASK_PP(16'h17F07,4);
TASK_PP(16'h17F08,4);
TASK_PP(16'h17F09,4);
TASK_PP(16'h17F0A,4);
TASK_PP(16'h17F0B,4);
TASK_PP(16'h17F0C,4);
TASK_PP(16'h17F0D,4);
TASK_PP(16'h17F0E,4);
TASK_PP(16'h17F0F,4);
TASK_PP(16'h17F10,4);
TASK_PP(16'h17F11,4);
TASK_PP(16'h17F12,4);
TASK_PP(16'h17F13,4);
TASK_PP(16'h17F14,4);
TASK_PP(16'h17F15,4);
TASK_PP(16'h17F16,4);
TASK_PP(16'h17F17,4);
TASK_PP(16'h17F18,4);
TASK_PP(16'h17F19,4);
TASK_PP(16'h17F1A,4);
TASK_PP(16'h17F1B,4);
TASK_PP(16'h17F1C,4);
TASK_PP(16'h17F1D,4);
TASK_PP(16'h17F1E,4);
TASK_PP(16'h17F1F,4);
TASK_PP(16'h17F20,4);
TASK_PP(16'h17F21,4);
TASK_PP(16'h17F22,4);
TASK_PP(16'h17F23,4);
TASK_PP(16'h17F24,4);
TASK_PP(16'h17F25,4);
TASK_PP(16'h17F26,4);
TASK_PP(16'h17F27,4);
TASK_PP(16'h17F28,4);
TASK_PP(16'h17F29,4);
TASK_PP(16'h17F2A,4);
TASK_PP(16'h17F2B,4);
TASK_PP(16'h17F2C,4);
TASK_PP(16'h17F2D,4);
TASK_PP(16'h17F2E,4);
TASK_PP(16'h17F2F,4);
TASK_PP(16'h17F30,4);
TASK_PP(16'h17F31,4);
TASK_PP(16'h17F32,4);
TASK_PP(16'h17F33,4);
TASK_PP(16'h17F34,4);
TASK_PP(16'h17F35,4);
TASK_PP(16'h17F36,4);
TASK_PP(16'h17F37,4);
TASK_PP(16'h17F38,4);
TASK_PP(16'h17F39,4);
TASK_PP(16'h17F3A,4);
TASK_PP(16'h17F3B,4);
TASK_PP(16'h17F3C,4);
TASK_PP(16'h17F3D,4);
TASK_PP(16'h17F3E,4);
TASK_PP(16'h17F3F,4);
TASK_PP(16'h17F40,4);
TASK_PP(16'h17F41,4);
TASK_PP(16'h17F42,4);
TASK_PP(16'h17F43,4);
TASK_PP(16'h17F44,4);
TASK_PP(16'h17F45,4);
TASK_PP(16'h17F46,4);
TASK_PP(16'h17F47,4);
TASK_PP(16'h17F48,4);
TASK_PP(16'h17F49,4);
TASK_PP(16'h17F4A,4);
TASK_PP(16'h17F4B,4);
TASK_PP(16'h17F4C,4);
TASK_PP(16'h17F4D,4);
TASK_PP(16'h17F4E,4);
TASK_PP(16'h17F4F,4);
TASK_PP(16'h17F50,4);
TASK_PP(16'h17F51,4);
TASK_PP(16'h17F52,4);
TASK_PP(16'h17F53,4);
TASK_PP(16'h17F54,4);
TASK_PP(16'h17F55,4);
TASK_PP(16'h17F56,4);
TASK_PP(16'h17F57,4);
TASK_PP(16'h17F58,4);
TASK_PP(16'h17F59,4);
TASK_PP(16'h17F5A,4);
TASK_PP(16'h17F5B,4);
TASK_PP(16'h17F5C,4);
TASK_PP(16'h17F5D,4);
TASK_PP(16'h17F5E,4);
TASK_PP(16'h17F5F,4);
TASK_PP(16'h17F60,4);
TASK_PP(16'h17F61,4);
TASK_PP(16'h17F62,4);
TASK_PP(16'h17F63,4);
TASK_PP(16'h17F64,4);
TASK_PP(16'h17F65,4);
TASK_PP(16'h17F66,4);
TASK_PP(16'h17F67,4);
TASK_PP(16'h17F68,4);
TASK_PP(16'h17F69,4);
TASK_PP(16'h17F6A,4);
TASK_PP(16'h17F6B,4);
TASK_PP(16'h17F6C,4);
TASK_PP(16'h17F6D,4);
TASK_PP(16'h17F6E,4);
TASK_PP(16'h17F6F,4);
TASK_PP(16'h17F70,4);
TASK_PP(16'h17F71,4);
TASK_PP(16'h17F72,4);
TASK_PP(16'h17F73,4);
TASK_PP(16'h17F74,4);
TASK_PP(16'h17F75,4);
TASK_PP(16'h17F76,4);
TASK_PP(16'h17F77,4);
TASK_PP(16'h17F78,4);
TASK_PP(16'h17F79,4);
TASK_PP(16'h17F7A,4);
TASK_PP(16'h17F7B,4);
TASK_PP(16'h17F7C,4);
TASK_PP(16'h17F7D,4);
TASK_PP(16'h17F7E,4);
TASK_PP(16'h17F7F,4);
TASK_PP(16'h17F80,4);
TASK_PP(16'h17F81,4);
TASK_PP(16'h17F82,4);
TASK_PP(16'h17F83,4);
TASK_PP(16'h17F84,4);
TASK_PP(16'h17F85,4);
TASK_PP(16'h17F86,4);
TASK_PP(16'h17F87,4);
TASK_PP(16'h17F88,4);
TASK_PP(16'h17F89,4);
TASK_PP(16'h17F8A,4);
TASK_PP(16'h17F8B,4);
TASK_PP(16'h17F8C,4);
TASK_PP(16'h17F8D,4);
TASK_PP(16'h17F8E,4);
TASK_PP(16'h17F8F,4);
TASK_PP(16'h17F90,4);
TASK_PP(16'h17F91,4);
TASK_PP(16'h17F92,4);
TASK_PP(16'h17F93,4);
TASK_PP(16'h17F94,4);
TASK_PP(16'h17F95,4);
TASK_PP(16'h17F96,4);
TASK_PP(16'h17F97,4);
TASK_PP(16'h17F98,4);
TASK_PP(16'h17F99,4);
TASK_PP(16'h17F9A,4);
TASK_PP(16'h17F9B,4);
TASK_PP(16'h17F9C,4);
TASK_PP(16'h17F9D,4);
TASK_PP(16'h17F9E,4);
TASK_PP(16'h17F9F,4);
TASK_PP(16'h17FA0,4);
TASK_PP(16'h17FA1,4);
TASK_PP(16'h17FA2,4);
TASK_PP(16'h17FA3,4);
TASK_PP(16'h17FA4,4);
TASK_PP(16'h17FA5,4);
TASK_PP(16'h17FA6,4);
TASK_PP(16'h17FA7,4);
TASK_PP(16'h17FA8,4);
TASK_PP(16'h17FA9,4);
TASK_PP(16'h17FAA,4);
TASK_PP(16'h17FAB,4);
TASK_PP(16'h17FAC,4);
TASK_PP(16'h17FAD,4);
TASK_PP(16'h17FAE,4);
TASK_PP(16'h17FAF,4);
TASK_PP(16'h17FB0,4);
TASK_PP(16'h17FB1,4);
TASK_PP(16'h17FB2,4);
TASK_PP(16'h17FB3,4);
TASK_PP(16'h17FB4,4);
TASK_PP(16'h17FB5,4);
TASK_PP(16'h17FB6,4);
TASK_PP(16'h17FB7,4);
TASK_PP(16'h17FB8,4);
TASK_PP(16'h17FB9,4);
TASK_PP(16'h17FBA,4);
TASK_PP(16'h17FBB,4);
TASK_PP(16'h17FBC,4);
TASK_PP(16'h17FBD,4);
TASK_PP(16'h17FBE,4);
TASK_PP(16'h17FBF,4);
TASK_PP(16'h17FC0,4);
TASK_PP(16'h17FC1,4);
TASK_PP(16'h17FC2,4);
TASK_PP(16'h17FC3,4);
TASK_PP(16'h17FC4,4);
TASK_PP(16'h17FC5,4);
TASK_PP(16'h17FC6,4);
TASK_PP(16'h17FC7,4);
TASK_PP(16'h17FC8,4);
TASK_PP(16'h17FC9,4);
TASK_PP(16'h17FCA,4);
TASK_PP(16'h17FCB,4);
TASK_PP(16'h17FCC,4);
TASK_PP(16'h17FCD,4);
TASK_PP(16'h17FCE,4);
TASK_PP(16'h17FCF,4);
TASK_PP(16'h17FD0,4);
TASK_PP(16'h17FD1,4);
TASK_PP(16'h17FD2,4);
TASK_PP(16'h17FD3,4);
TASK_PP(16'h17FD4,4);
TASK_PP(16'h17FD5,4);
TASK_PP(16'h17FD6,4);
TASK_PP(16'h17FD7,4);
TASK_PP(16'h17FD8,4);
TASK_PP(16'h17FD9,4);
TASK_PP(16'h17FDA,4);
TASK_PP(16'h17FDB,4);
TASK_PP(16'h17FDC,4);
TASK_PP(16'h17FDD,4);
TASK_PP(16'h17FDE,4);
TASK_PP(16'h17FDF,4);
TASK_PP(16'h17FE0,4);
TASK_PP(16'h17FE1,4);
TASK_PP(16'h17FE2,4);
TASK_PP(16'h17FE3,4);
TASK_PP(16'h17FE4,4);
TASK_PP(16'h17FE5,4);
TASK_PP(16'h17FE6,4);
TASK_PP(16'h17FE7,4);
TASK_PP(16'h17FE8,4);
TASK_PP(16'h17FE9,4);
TASK_PP(16'h17FEA,4);
TASK_PP(16'h17FEB,4);
TASK_PP(16'h17FEC,4);
TASK_PP(16'h17FED,4);
TASK_PP(16'h17FEE,4);
TASK_PP(16'h17FEF,4);
TASK_PP(16'h17FF0,4);
TASK_PP(16'h17FF1,4);
TASK_PP(16'h17FF2,4);
TASK_PP(16'h17FF3,4);
TASK_PP(16'h17FF4,4);
TASK_PP(16'h17FF5,4);
TASK_PP(16'h17FF6,4);
TASK_PP(16'h17FF7,4);
TASK_PP(16'h17FF8,4);
TASK_PP(16'h17FF9,4);
TASK_PP(16'h17FFA,4);
TASK_PP(16'h17FFB,4);
TASK_PP(16'h17FFC,4);
TASK_PP(16'h17FFD,4);
TASK_PP(16'h17FFE,4);
TASK_PP(16'h17FFF,4);
TASK_PP(16'h18000,4);
TASK_PP(16'h18001,4);
TASK_PP(16'h18002,4);
TASK_PP(16'h18003,4);
TASK_PP(16'h18004,4);
TASK_PP(16'h18005,4);
TASK_PP(16'h18006,4);
TASK_PP(16'h18007,4);
TASK_PP(16'h18008,4);
TASK_PP(16'h18009,4);
TASK_PP(16'h1800A,4);
TASK_PP(16'h1800B,4);
TASK_PP(16'h1800C,4);
TASK_PP(16'h1800D,4);
TASK_PP(16'h1800E,4);
TASK_PP(16'h1800F,4);
TASK_PP(16'h18010,4);
TASK_PP(16'h18011,4);
TASK_PP(16'h18012,4);
TASK_PP(16'h18013,4);
TASK_PP(16'h18014,4);
TASK_PP(16'h18015,4);
TASK_PP(16'h18016,4);
TASK_PP(16'h18017,4);
TASK_PP(16'h18018,4);
TASK_PP(16'h18019,4);
TASK_PP(16'h1801A,4);
TASK_PP(16'h1801B,4);
TASK_PP(16'h1801C,4);
TASK_PP(16'h1801D,4);
TASK_PP(16'h1801E,4);
TASK_PP(16'h1801F,4);
TASK_PP(16'h18020,4);
TASK_PP(16'h18021,4);
TASK_PP(16'h18022,4);
TASK_PP(16'h18023,4);
TASK_PP(16'h18024,4);
TASK_PP(16'h18025,4);
TASK_PP(16'h18026,4);
TASK_PP(16'h18027,4);
TASK_PP(16'h18028,4);
TASK_PP(16'h18029,4);
TASK_PP(16'h1802A,4);
TASK_PP(16'h1802B,4);
TASK_PP(16'h1802C,4);
TASK_PP(16'h1802D,4);
TASK_PP(16'h1802E,4);
TASK_PP(16'h1802F,4);
TASK_PP(16'h18030,4);
TASK_PP(16'h18031,4);
TASK_PP(16'h18032,4);
TASK_PP(16'h18033,4);
TASK_PP(16'h18034,4);
TASK_PP(16'h18035,4);
TASK_PP(16'h18036,4);
TASK_PP(16'h18037,4);
TASK_PP(16'h18038,4);
TASK_PP(16'h18039,4);
TASK_PP(16'h1803A,4);
TASK_PP(16'h1803B,4);
TASK_PP(16'h1803C,4);
TASK_PP(16'h1803D,4);
TASK_PP(16'h1803E,4);
TASK_PP(16'h1803F,4);
TASK_PP(16'h18040,4);
TASK_PP(16'h18041,4);
TASK_PP(16'h18042,4);
TASK_PP(16'h18043,4);
TASK_PP(16'h18044,4);
TASK_PP(16'h18045,4);
TASK_PP(16'h18046,4);
TASK_PP(16'h18047,4);
TASK_PP(16'h18048,4);
TASK_PP(16'h18049,4);
TASK_PP(16'h1804A,4);
TASK_PP(16'h1804B,4);
TASK_PP(16'h1804C,4);
TASK_PP(16'h1804D,4);
TASK_PP(16'h1804E,4);
TASK_PP(16'h1804F,4);
TASK_PP(16'h18050,4);
TASK_PP(16'h18051,4);
TASK_PP(16'h18052,4);
TASK_PP(16'h18053,4);
TASK_PP(16'h18054,4);
TASK_PP(16'h18055,4);
TASK_PP(16'h18056,4);
TASK_PP(16'h18057,4);
TASK_PP(16'h18058,4);
TASK_PP(16'h18059,4);
TASK_PP(16'h1805A,4);
TASK_PP(16'h1805B,4);
TASK_PP(16'h1805C,4);
TASK_PP(16'h1805D,4);
TASK_PP(16'h1805E,4);
TASK_PP(16'h1805F,4);
TASK_PP(16'h18060,4);
TASK_PP(16'h18061,4);
TASK_PP(16'h18062,4);
TASK_PP(16'h18063,4);
TASK_PP(16'h18064,4);
TASK_PP(16'h18065,4);
TASK_PP(16'h18066,4);
TASK_PP(16'h18067,4);
TASK_PP(16'h18068,4);
TASK_PP(16'h18069,4);
TASK_PP(16'h1806A,4);
TASK_PP(16'h1806B,4);
TASK_PP(16'h1806C,4);
TASK_PP(16'h1806D,4);
TASK_PP(16'h1806E,4);
TASK_PP(16'h1806F,4);
TASK_PP(16'h18070,4);
TASK_PP(16'h18071,4);
TASK_PP(16'h18072,4);
TASK_PP(16'h18073,4);
TASK_PP(16'h18074,4);
TASK_PP(16'h18075,4);
TASK_PP(16'h18076,4);
TASK_PP(16'h18077,4);
TASK_PP(16'h18078,4);
TASK_PP(16'h18079,4);
TASK_PP(16'h1807A,4);
TASK_PP(16'h1807B,4);
TASK_PP(16'h1807C,4);
TASK_PP(16'h1807D,4);
TASK_PP(16'h1807E,4);
TASK_PP(16'h1807F,4);
TASK_PP(16'h18080,4);
TASK_PP(16'h18081,4);
TASK_PP(16'h18082,4);
TASK_PP(16'h18083,4);
TASK_PP(16'h18084,4);
TASK_PP(16'h18085,4);
TASK_PP(16'h18086,4);
TASK_PP(16'h18087,4);
TASK_PP(16'h18088,4);
TASK_PP(16'h18089,4);
TASK_PP(16'h1808A,4);
TASK_PP(16'h1808B,4);
TASK_PP(16'h1808C,4);
TASK_PP(16'h1808D,4);
TASK_PP(16'h1808E,4);
TASK_PP(16'h1808F,4);
TASK_PP(16'h18090,4);
TASK_PP(16'h18091,4);
TASK_PP(16'h18092,4);
TASK_PP(16'h18093,4);
TASK_PP(16'h18094,4);
TASK_PP(16'h18095,4);
TASK_PP(16'h18096,4);
TASK_PP(16'h18097,4);
TASK_PP(16'h18098,4);
TASK_PP(16'h18099,4);
TASK_PP(16'h1809A,4);
TASK_PP(16'h1809B,4);
TASK_PP(16'h1809C,4);
TASK_PP(16'h1809D,4);
TASK_PP(16'h1809E,4);
TASK_PP(16'h1809F,4);
TASK_PP(16'h180A0,4);
TASK_PP(16'h180A1,4);
TASK_PP(16'h180A2,4);
TASK_PP(16'h180A3,4);
TASK_PP(16'h180A4,4);
TASK_PP(16'h180A5,4);
TASK_PP(16'h180A6,4);
TASK_PP(16'h180A7,4);
TASK_PP(16'h180A8,4);
TASK_PP(16'h180A9,4);
TASK_PP(16'h180AA,4);
TASK_PP(16'h180AB,4);
TASK_PP(16'h180AC,4);
TASK_PP(16'h180AD,4);
TASK_PP(16'h180AE,4);
TASK_PP(16'h180AF,4);
TASK_PP(16'h180B0,4);
TASK_PP(16'h180B1,4);
TASK_PP(16'h180B2,4);
TASK_PP(16'h180B3,4);
TASK_PP(16'h180B4,4);
TASK_PP(16'h180B5,4);
TASK_PP(16'h180B6,4);
TASK_PP(16'h180B7,4);
TASK_PP(16'h180B8,4);
TASK_PP(16'h180B9,4);
TASK_PP(16'h180BA,4);
TASK_PP(16'h180BB,4);
TASK_PP(16'h180BC,4);
TASK_PP(16'h180BD,4);
TASK_PP(16'h180BE,4);
TASK_PP(16'h180BF,4);
TASK_PP(16'h180C0,4);
TASK_PP(16'h180C1,4);
TASK_PP(16'h180C2,4);
TASK_PP(16'h180C3,4);
TASK_PP(16'h180C4,4);
TASK_PP(16'h180C5,4);
TASK_PP(16'h180C6,4);
TASK_PP(16'h180C7,4);
TASK_PP(16'h180C8,4);
TASK_PP(16'h180C9,4);
TASK_PP(16'h180CA,4);
TASK_PP(16'h180CB,4);
TASK_PP(16'h180CC,4);
TASK_PP(16'h180CD,4);
TASK_PP(16'h180CE,4);
TASK_PP(16'h180CF,4);
TASK_PP(16'h180D0,4);
TASK_PP(16'h180D1,4);
TASK_PP(16'h180D2,4);
TASK_PP(16'h180D3,4);
TASK_PP(16'h180D4,4);
TASK_PP(16'h180D5,4);
TASK_PP(16'h180D6,4);
TASK_PP(16'h180D7,4);
TASK_PP(16'h180D8,4);
TASK_PP(16'h180D9,4);
TASK_PP(16'h180DA,4);
TASK_PP(16'h180DB,4);
TASK_PP(16'h180DC,4);
TASK_PP(16'h180DD,4);
TASK_PP(16'h180DE,4);
TASK_PP(16'h180DF,4);
TASK_PP(16'h180E0,4);
TASK_PP(16'h180E1,4);
TASK_PP(16'h180E2,4);
TASK_PP(16'h180E3,4);
TASK_PP(16'h180E4,4);
TASK_PP(16'h180E5,4);
TASK_PP(16'h180E6,4);
TASK_PP(16'h180E7,4);
TASK_PP(16'h180E8,4);
TASK_PP(16'h180E9,4);
TASK_PP(16'h180EA,4);
TASK_PP(16'h180EB,4);
TASK_PP(16'h180EC,4);
TASK_PP(16'h180ED,4);
TASK_PP(16'h180EE,4);
TASK_PP(16'h180EF,4);
TASK_PP(16'h180F0,4);
TASK_PP(16'h180F1,4);
TASK_PP(16'h180F2,4);
TASK_PP(16'h180F3,4);
TASK_PP(16'h180F4,4);
TASK_PP(16'h180F5,4);
TASK_PP(16'h180F6,4);
TASK_PP(16'h180F7,4);
TASK_PP(16'h180F8,4);
TASK_PP(16'h180F9,4);
TASK_PP(16'h180FA,4);
TASK_PP(16'h180FB,4);
TASK_PP(16'h180FC,4);
TASK_PP(16'h180FD,4);
TASK_PP(16'h180FE,4);
TASK_PP(16'h180FF,4);
TASK_PP(16'h18100,4);
TASK_PP(16'h18101,4);
TASK_PP(16'h18102,4);
TASK_PP(16'h18103,4);
TASK_PP(16'h18104,4);
TASK_PP(16'h18105,4);
TASK_PP(16'h18106,4);
TASK_PP(16'h18107,4);
TASK_PP(16'h18108,4);
TASK_PP(16'h18109,4);
TASK_PP(16'h1810A,4);
TASK_PP(16'h1810B,4);
TASK_PP(16'h1810C,4);
TASK_PP(16'h1810D,4);
TASK_PP(16'h1810E,4);
TASK_PP(16'h1810F,4);
TASK_PP(16'h18110,4);
TASK_PP(16'h18111,4);
TASK_PP(16'h18112,4);
TASK_PP(16'h18113,4);
TASK_PP(16'h18114,4);
TASK_PP(16'h18115,4);
TASK_PP(16'h18116,4);
TASK_PP(16'h18117,4);
TASK_PP(16'h18118,4);
TASK_PP(16'h18119,4);
TASK_PP(16'h1811A,4);
TASK_PP(16'h1811B,4);
TASK_PP(16'h1811C,4);
TASK_PP(16'h1811D,4);
TASK_PP(16'h1811E,4);
TASK_PP(16'h1811F,4);
TASK_PP(16'h18120,4);
TASK_PP(16'h18121,4);
TASK_PP(16'h18122,4);
TASK_PP(16'h18123,4);
TASK_PP(16'h18124,4);
TASK_PP(16'h18125,4);
TASK_PP(16'h18126,4);
TASK_PP(16'h18127,4);
TASK_PP(16'h18128,4);
TASK_PP(16'h18129,4);
TASK_PP(16'h1812A,4);
TASK_PP(16'h1812B,4);
TASK_PP(16'h1812C,4);
TASK_PP(16'h1812D,4);
TASK_PP(16'h1812E,4);
TASK_PP(16'h1812F,4);
TASK_PP(16'h18130,4);
TASK_PP(16'h18131,4);
TASK_PP(16'h18132,4);
TASK_PP(16'h18133,4);
TASK_PP(16'h18134,4);
TASK_PP(16'h18135,4);
TASK_PP(16'h18136,4);
TASK_PP(16'h18137,4);
TASK_PP(16'h18138,4);
TASK_PP(16'h18139,4);
TASK_PP(16'h1813A,4);
TASK_PP(16'h1813B,4);
TASK_PP(16'h1813C,4);
TASK_PP(16'h1813D,4);
TASK_PP(16'h1813E,4);
TASK_PP(16'h1813F,4);
TASK_PP(16'h18140,4);
TASK_PP(16'h18141,4);
TASK_PP(16'h18142,4);
TASK_PP(16'h18143,4);
TASK_PP(16'h18144,4);
TASK_PP(16'h18145,4);
TASK_PP(16'h18146,4);
TASK_PP(16'h18147,4);
TASK_PP(16'h18148,4);
TASK_PP(16'h18149,4);
TASK_PP(16'h1814A,4);
TASK_PP(16'h1814B,4);
TASK_PP(16'h1814C,4);
TASK_PP(16'h1814D,4);
TASK_PP(16'h1814E,4);
TASK_PP(16'h1814F,4);
TASK_PP(16'h18150,4);
TASK_PP(16'h18151,4);
TASK_PP(16'h18152,4);
TASK_PP(16'h18153,4);
TASK_PP(16'h18154,4);
TASK_PP(16'h18155,4);
TASK_PP(16'h18156,4);
TASK_PP(16'h18157,4);
TASK_PP(16'h18158,4);
TASK_PP(16'h18159,4);
TASK_PP(16'h1815A,4);
TASK_PP(16'h1815B,4);
TASK_PP(16'h1815C,4);
TASK_PP(16'h1815D,4);
TASK_PP(16'h1815E,4);
TASK_PP(16'h1815F,4);
TASK_PP(16'h18160,4);
TASK_PP(16'h18161,4);
TASK_PP(16'h18162,4);
TASK_PP(16'h18163,4);
TASK_PP(16'h18164,4);
TASK_PP(16'h18165,4);
TASK_PP(16'h18166,4);
TASK_PP(16'h18167,4);
TASK_PP(16'h18168,4);
TASK_PP(16'h18169,4);
TASK_PP(16'h1816A,4);
TASK_PP(16'h1816B,4);
TASK_PP(16'h1816C,4);
TASK_PP(16'h1816D,4);
TASK_PP(16'h1816E,4);
TASK_PP(16'h1816F,4);
TASK_PP(16'h18170,4);
TASK_PP(16'h18171,4);
TASK_PP(16'h18172,4);
TASK_PP(16'h18173,4);
TASK_PP(16'h18174,4);
TASK_PP(16'h18175,4);
TASK_PP(16'h18176,4);
TASK_PP(16'h18177,4);
TASK_PP(16'h18178,4);
TASK_PP(16'h18179,4);
TASK_PP(16'h1817A,4);
TASK_PP(16'h1817B,4);
TASK_PP(16'h1817C,4);
TASK_PP(16'h1817D,4);
TASK_PP(16'h1817E,4);
TASK_PP(16'h1817F,4);
TASK_PP(16'h18180,4);
TASK_PP(16'h18181,4);
TASK_PP(16'h18182,4);
TASK_PP(16'h18183,4);
TASK_PP(16'h18184,4);
TASK_PP(16'h18185,4);
TASK_PP(16'h18186,4);
TASK_PP(16'h18187,4);
TASK_PP(16'h18188,4);
TASK_PP(16'h18189,4);
TASK_PP(16'h1818A,4);
TASK_PP(16'h1818B,4);
TASK_PP(16'h1818C,4);
TASK_PP(16'h1818D,4);
TASK_PP(16'h1818E,4);
TASK_PP(16'h1818F,4);
TASK_PP(16'h18190,4);
TASK_PP(16'h18191,4);
TASK_PP(16'h18192,4);
TASK_PP(16'h18193,4);
TASK_PP(16'h18194,4);
TASK_PP(16'h18195,4);
TASK_PP(16'h18196,4);
TASK_PP(16'h18197,4);
TASK_PP(16'h18198,4);
TASK_PP(16'h18199,4);
TASK_PP(16'h1819A,4);
TASK_PP(16'h1819B,4);
TASK_PP(16'h1819C,4);
TASK_PP(16'h1819D,4);
TASK_PP(16'h1819E,4);
TASK_PP(16'h1819F,4);
TASK_PP(16'h181A0,4);
TASK_PP(16'h181A1,4);
TASK_PP(16'h181A2,4);
TASK_PP(16'h181A3,4);
TASK_PP(16'h181A4,4);
TASK_PP(16'h181A5,4);
TASK_PP(16'h181A6,4);
TASK_PP(16'h181A7,4);
TASK_PP(16'h181A8,4);
TASK_PP(16'h181A9,4);
TASK_PP(16'h181AA,4);
TASK_PP(16'h181AB,4);
TASK_PP(16'h181AC,4);
TASK_PP(16'h181AD,4);
TASK_PP(16'h181AE,4);
TASK_PP(16'h181AF,4);
TASK_PP(16'h181B0,4);
TASK_PP(16'h181B1,4);
TASK_PP(16'h181B2,4);
TASK_PP(16'h181B3,4);
TASK_PP(16'h181B4,4);
TASK_PP(16'h181B5,4);
TASK_PP(16'h181B6,4);
TASK_PP(16'h181B7,4);
TASK_PP(16'h181B8,4);
TASK_PP(16'h181B9,4);
TASK_PP(16'h181BA,4);
TASK_PP(16'h181BB,4);
TASK_PP(16'h181BC,4);
TASK_PP(16'h181BD,4);
TASK_PP(16'h181BE,4);
TASK_PP(16'h181BF,4);
TASK_PP(16'h181C0,4);
TASK_PP(16'h181C1,4);
TASK_PP(16'h181C2,4);
TASK_PP(16'h181C3,4);
TASK_PP(16'h181C4,4);
TASK_PP(16'h181C5,4);
TASK_PP(16'h181C6,4);
TASK_PP(16'h181C7,4);
TASK_PP(16'h181C8,4);
TASK_PP(16'h181C9,4);
TASK_PP(16'h181CA,4);
TASK_PP(16'h181CB,4);
TASK_PP(16'h181CC,4);
TASK_PP(16'h181CD,4);
TASK_PP(16'h181CE,4);
TASK_PP(16'h181CF,4);
TASK_PP(16'h181D0,4);
TASK_PP(16'h181D1,4);
TASK_PP(16'h181D2,4);
TASK_PP(16'h181D3,4);
TASK_PP(16'h181D4,4);
TASK_PP(16'h181D5,4);
TASK_PP(16'h181D6,4);
TASK_PP(16'h181D7,4);
TASK_PP(16'h181D8,4);
TASK_PP(16'h181D9,4);
TASK_PP(16'h181DA,4);
TASK_PP(16'h181DB,4);
TASK_PP(16'h181DC,4);
TASK_PP(16'h181DD,4);
TASK_PP(16'h181DE,4);
TASK_PP(16'h181DF,4);
TASK_PP(16'h181E0,4);
TASK_PP(16'h181E1,4);
TASK_PP(16'h181E2,4);
TASK_PP(16'h181E3,4);
TASK_PP(16'h181E4,4);
TASK_PP(16'h181E5,4);
TASK_PP(16'h181E6,4);
TASK_PP(16'h181E7,4);
TASK_PP(16'h181E8,4);
TASK_PP(16'h181E9,4);
TASK_PP(16'h181EA,4);
TASK_PP(16'h181EB,4);
TASK_PP(16'h181EC,4);
TASK_PP(16'h181ED,4);
TASK_PP(16'h181EE,4);
TASK_PP(16'h181EF,4);
TASK_PP(16'h181F0,4);
TASK_PP(16'h181F1,4);
TASK_PP(16'h181F2,4);
TASK_PP(16'h181F3,4);
TASK_PP(16'h181F4,4);
TASK_PP(16'h181F5,4);
TASK_PP(16'h181F6,4);
TASK_PP(16'h181F7,4);
TASK_PP(16'h181F8,4);
TASK_PP(16'h181F9,4);
TASK_PP(16'h181FA,4);
TASK_PP(16'h181FB,4);
TASK_PP(16'h181FC,4);
TASK_PP(16'h181FD,4);
TASK_PP(16'h181FE,4);
TASK_PP(16'h181FF,4);
TASK_PP(16'h18200,4);
TASK_PP(16'h18201,4);
TASK_PP(16'h18202,4);
TASK_PP(16'h18203,4);
TASK_PP(16'h18204,4);
TASK_PP(16'h18205,4);
TASK_PP(16'h18206,4);
TASK_PP(16'h18207,4);
TASK_PP(16'h18208,4);
TASK_PP(16'h18209,4);
TASK_PP(16'h1820A,4);
TASK_PP(16'h1820B,4);
TASK_PP(16'h1820C,4);
TASK_PP(16'h1820D,4);
TASK_PP(16'h1820E,4);
TASK_PP(16'h1820F,4);
TASK_PP(16'h18210,4);
TASK_PP(16'h18211,4);
TASK_PP(16'h18212,4);
TASK_PP(16'h18213,4);
TASK_PP(16'h18214,4);
TASK_PP(16'h18215,4);
TASK_PP(16'h18216,4);
TASK_PP(16'h18217,4);
TASK_PP(16'h18218,4);
TASK_PP(16'h18219,4);
TASK_PP(16'h1821A,4);
TASK_PP(16'h1821B,4);
TASK_PP(16'h1821C,4);
TASK_PP(16'h1821D,4);
TASK_PP(16'h1821E,4);
TASK_PP(16'h1821F,4);
TASK_PP(16'h18220,4);
TASK_PP(16'h18221,4);
TASK_PP(16'h18222,4);
TASK_PP(16'h18223,4);
TASK_PP(16'h18224,4);
TASK_PP(16'h18225,4);
TASK_PP(16'h18226,4);
TASK_PP(16'h18227,4);
TASK_PP(16'h18228,4);
TASK_PP(16'h18229,4);
TASK_PP(16'h1822A,4);
TASK_PP(16'h1822B,4);
TASK_PP(16'h1822C,4);
TASK_PP(16'h1822D,4);
TASK_PP(16'h1822E,4);
TASK_PP(16'h1822F,4);
TASK_PP(16'h18230,4);
TASK_PP(16'h18231,4);
TASK_PP(16'h18232,4);
TASK_PP(16'h18233,4);
TASK_PP(16'h18234,4);
TASK_PP(16'h18235,4);
TASK_PP(16'h18236,4);
TASK_PP(16'h18237,4);
TASK_PP(16'h18238,4);
TASK_PP(16'h18239,4);
TASK_PP(16'h1823A,4);
TASK_PP(16'h1823B,4);
TASK_PP(16'h1823C,4);
TASK_PP(16'h1823D,4);
TASK_PP(16'h1823E,4);
TASK_PP(16'h1823F,4);
TASK_PP(16'h18240,4);
TASK_PP(16'h18241,4);
TASK_PP(16'h18242,4);
TASK_PP(16'h18243,4);
TASK_PP(16'h18244,4);
TASK_PP(16'h18245,4);
TASK_PP(16'h18246,4);
TASK_PP(16'h18247,4);
TASK_PP(16'h18248,4);
TASK_PP(16'h18249,4);
TASK_PP(16'h1824A,4);
TASK_PP(16'h1824B,4);
TASK_PP(16'h1824C,4);
TASK_PP(16'h1824D,4);
TASK_PP(16'h1824E,4);
TASK_PP(16'h1824F,4);
TASK_PP(16'h18250,4);
TASK_PP(16'h18251,4);
TASK_PP(16'h18252,4);
TASK_PP(16'h18253,4);
TASK_PP(16'h18254,4);
TASK_PP(16'h18255,4);
TASK_PP(16'h18256,4);
TASK_PP(16'h18257,4);
TASK_PP(16'h18258,4);
TASK_PP(16'h18259,4);
TASK_PP(16'h1825A,4);
TASK_PP(16'h1825B,4);
TASK_PP(16'h1825C,4);
TASK_PP(16'h1825D,4);
TASK_PP(16'h1825E,4);
TASK_PP(16'h1825F,4);
TASK_PP(16'h18260,4);
TASK_PP(16'h18261,4);
TASK_PP(16'h18262,4);
TASK_PP(16'h18263,4);
TASK_PP(16'h18264,4);
TASK_PP(16'h18265,4);
TASK_PP(16'h18266,4);
TASK_PP(16'h18267,4);
TASK_PP(16'h18268,4);
TASK_PP(16'h18269,4);
TASK_PP(16'h1826A,4);
TASK_PP(16'h1826B,4);
TASK_PP(16'h1826C,4);
TASK_PP(16'h1826D,4);
TASK_PP(16'h1826E,4);
TASK_PP(16'h1826F,4);
TASK_PP(16'h18270,4);
TASK_PP(16'h18271,4);
TASK_PP(16'h18272,4);
TASK_PP(16'h18273,4);
TASK_PP(16'h18274,4);
TASK_PP(16'h18275,4);
TASK_PP(16'h18276,4);
TASK_PP(16'h18277,4);
TASK_PP(16'h18278,4);
TASK_PP(16'h18279,4);
TASK_PP(16'h1827A,4);
TASK_PP(16'h1827B,4);
TASK_PP(16'h1827C,4);
TASK_PP(16'h1827D,4);
TASK_PP(16'h1827E,4);
TASK_PP(16'h1827F,4);
TASK_PP(16'h18280,4);
TASK_PP(16'h18281,4);
TASK_PP(16'h18282,4);
TASK_PP(16'h18283,4);
TASK_PP(16'h18284,4);
TASK_PP(16'h18285,4);
TASK_PP(16'h18286,4);
TASK_PP(16'h18287,4);
TASK_PP(16'h18288,4);
TASK_PP(16'h18289,4);
TASK_PP(16'h1828A,4);
TASK_PP(16'h1828B,4);
TASK_PP(16'h1828C,4);
TASK_PP(16'h1828D,4);
TASK_PP(16'h1828E,4);
TASK_PP(16'h1828F,4);
TASK_PP(16'h18290,4);
TASK_PP(16'h18291,4);
TASK_PP(16'h18292,4);
TASK_PP(16'h18293,4);
TASK_PP(16'h18294,4);
TASK_PP(16'h18295,4);
TASK_PP(16'h18296,4);
TASK_PP(16'h18297,4);
TASK_PP(16'h18298,4);
TASK_PP(16'h18299,4);
TASK_PP(16'h1829A,4);
TASK_PP(16'h1829B,4);
TASK_PP(16'h1829C,4);
TASK_PP(16'h1829D,4);
TASK_PP(16'h1829E,4);
TASK_PP(16'h1829F,4);
TASK_PP(16'h182A0,4);
TASK_PP(16'h182A1,4);
TASK_PP(16'h182A2,4);
TASK_PP(16'h182A3,4);
TASK_PP(16'h182A4,4);
TASK_PP(16'h182A5,4);
TASK_PP(16'h182A6,4);
TASK_PP(16'h182A7,4);
TASK_PP(16'h182A8,4);
TASK_PP(16'h182A9,4);
TASK_PP(16'h182AA,4);
TASK_PP(16'h182AB,4);
TASK_PP(16'h182AC,4);
TASK_PP(16'h182AD,4);
TASK_PP(16'h182AE,4);
TASK_PP(16'h182AF,4);
TASK_PP(16'h182B0,4);
TASK_PP(16'h182B1,4);
TASK_PP(16'h182B2,4);
TASK_PP(16'h182B3,4);
TASK_PP(16'h182B4,4);
TASK_PP(16'h182B5,4);
TASK_PP(16'h182B6,4);
TASK_PP(16'h182B7,4);
TASK_PP(16'h182B8,4);
TASK_PP(16'h182B9,4);
TASK_PP(16'h182BA,4);
TASK_PP(16'h182BB,4);
TASK_PP(16'h182BC,4);
TASK_PP(16'h182BD,4);
TASK_PP(16'h182BE,4);
TASK_PP(16'h182BF,4);
TASK_PP(16'h182C0,4);
TASK_PP(16'h182C1,4);
TASK_PP(16'h182C2,4);
TASK_PP(16'h182C3,4);
TASK_PP(16'h182C4,4);
TASK_PP(16'h182C5,4);
TASK_PP(16'h182C6,4);
TASK_PP(16'h182C7,4);
TASK_PP(16'h182C8,4);
TASK_PP(16'h182C9,4);
TASK_PP(16'h182CA,4);
TASK_PP(16'h182CB,4);
TASK_PP(16'h182CC,4);
TASK_PP(16'h182CD,4);
TASK_PP(16'h182CE,4);
TASK_PP(16'h182CF,4);
TASK_PP(16'h182D0,4);
TASK_PP(16'h182D1,4);
TASK_PP(16'h182D2,4);
TASK_PP(16'h182D3,4);
TASK_PP(16'h182D4,4);
TASK_PP(16'h182D5,4);
TASK_PP(16'h182D6,4);
TASK_PP(16'h182D7,4);
TASK_PP(16'h182D8,4);
TASK_PP(16'h182D9,4);
TASK_PP(16'h182DA,4);
TASK_PP(16'h182DB,4);
TASK_PP(16'h182DC,4);
TASK_PP(16'h182DD,4);
TASK_PP(16'h182DE,4);
TASK_PP(16'h182DF,4);
TASK_PP(16'h182E0,4);
TASK_PP(16'h182E1,4);
TASK_PP(16'h182E2,4);
TASK_PP(16'h182E3,4);
TASK_PP(16'h182E4,4);
TASK_PP(16'h182E5,4);
TASK_PP(16'h182E6,4);
TASK_PP(16'h182E7,4);
TASK_PP(16'h182E8,4);
TASK_PP(16'h182E9,4);
TASK_PP(16'h182EA,4);
TASK_PP(16'h182EB,4);
TASK_PP(16'h182EC,4);
TASK_PP(16'h182ED,4);
TASK_PP(16'h182EE,4);
TASK_PP(16'h182EF,4);
TASK_PP(16'h182F0,4);
TASK_PP(16'h182F1,4);
TASK_PP(16'h182F2,4);
TASK_PP(16'h182F3,4);
TASK_PP(16'h182F4,4);
TASK_PP(16'h182F5,4);
TASK_PP(16'h182F6,4);
TASK_PP(16'h182F7,4);
TASK_PP(16'h182F8,4);
TASK_PP(16'h182F9,4);
TASK_PP(16'h182FA,4);
TASK_PP(16'h182FB,4);
TASK_PP(16'h182FC,4);
TASK_PP(16'h182FD,4);
TASK_PP(16'h182FE,4);
TASK_PP(16'h182FF,4);
TASK_PP(16'h18300,4);
TASK_PP(16'h18301,4);
TASK_PP(16'h18302,4);
TASK_PP(16'h18303,4);
TASK_PP(16'h18304,4);
TASK_PP(16'h18305,4);
TASK_PP(16'h18306,4);
TASK_PP(16'h18307,4);
TASK_PP(16'h18308,4);
TASK_PP(16'h18309,4);
TASK_PP(16'h1830A,4);
TASK_PP(16'h1830B,4);
TASK_PP(16'h1830C,4);
TASK_PP(16'h1830D,4);
TASK_PP(16'h1830E,4);
TASK_PP(16'h1830F,4);
TASK_PP(16'h18310,4);
TASK_PP(16'h18311,4);
TASK_PP(16'h18312,4);
TASK_PP(16'h18313,4);
TASK_PP(16'h18314,4);
TASK_PP(16'h18315,4);
TASK_PP(16'h18316,4);
TASK_PP(16'h18317,4);
TASK_PP(16'h18318,4);
TASK_PP(16'h18319,4);
TASK_PP(16'h1831A,4);
TASK_PP(16'h1831B,4);
TASK_PP(16'h1831C,4);
TASK_PP(16'h1831D,4);
TASK_PP(16'h1831E,4);
TASK_PP(16'h1831F,4);
TASK_PP(16'h18320,4);
TASK_PP(16'h18321,4);
TASK_PP(16'h18322,4);
TASK_PP(16'h18323,4);
TASK_PP(16'h18324,4);
TASK_PP(16'h18325,4);
TASK_PP(16'h18326,4);
TASK_PP(16'h18327,4);
TASK_PP(16'h18328,4);
TASK_PP(16'h18329,4);
TASK_PP(16'h1832A,4);
TASK_PP(16'h1832B,4);
TASK_PP(16'h1832C,4);
TASK_PP(16'h1832D,4);
TASK_PP(16'h1832E,4);
TASK_PP(16'h1832F,4);
TASK_PP(16'h18330,4);
TASK_PP(16'h18331,4);
TASK_PP(16'h18332,4);
TASK_PP(16'h18333,4);
TASK_PP(16'h18334,4);
TASK_PP(16'h18335,4);
TASK_PP(16'h18336,4);
TASK_PP(16'h18337,4);
TASK_PP(16'h18338,4);
TASK_PP(16'h18339,4);
TASK_PP(16'h1833A,4);
TASK_PP(16'h1833B,4);
TASK_PP(16'h1833C,4);
TASK_PP(16'h1833D,4);
TASK_PP(16'h1833E,4);
TASK_PP(16'h1833F,4);
TASK_PP(16'h18340,4);
TASK_PP(16'h18341,4);
TASK_PP(16'h18342,4);
TASK_PP(16'h18343,4);
TASK_PP(16'h18344,4);
TASK_PP(16'h18345,4);
TASK_PP(16'h18346,4);
TASK_PP(16'h18347,4);
TASK_PP(16'h18348,4);
TASK_PP(16'h18349,4);
TASK_PP(16'h1834A,4);
TASK_PP(16'h1834B,4);
TASK_PP(16'h1834C,4);
TASK_PP(16'h1834D,4);
TASK_PP(16'h1834E,4);
TASK_PP(16'h1834F,4);
TASK_PP(16'h18350,4);
TASK_PP(16'h18351,4);
TASK_PP(16'h18352,4);
TASK_PP(16'h18353,4);
TASK_PP(16'h18354,4);
TASK_PP(16'h18355,4);
TASK_PP(16'h18356,4);
TASK_PP(16'h18357,4);
TASK_PP(16'h18358,4);
TASK_PP(16'h18359,4);
TASK_PP(16'h1835A,4);
TASK_PP(16'h1835B,4);
TASK_PP(16'h1835C,4);
TASK_PP(16'h1835D,4);
TASK_PP(16'h1835E,4);
TASK_PP(16'h1835F,4);
TASK_PP(16'h18360,4);
TASK_PP(16'h18361,4);
TASK_PP(16'h18362,4);
TASK_PP(16'h18363,4);
TASK_PP(16'h18364,4);
TASK_PP(16'h18365,4);
TASK_PP(16'h18366,4);
TASK_PP(16'h18367,4);
TASK_PP(16'h18368,4);
TASK_PP(16'h18369,4);
TASK_PP(16'h1836A,4);
TASK_PP(16'h1836B,4);
TASK_PP(16'h1836C,4);
TASK_PP(16'h1836D,4);
TASK_PP(16'h1836E,4);
TASK_PP(16'h1836F,4);
TASK_PP(16'h18370,4);
TASK_PP(16'h18371,4);
TASK_PP(16'h18372,4);
TASK_PP(16'h18373,4);
TASK_PP(16'h18374,4);
TASK_PP(16'h18375,4);
TASK_PP(16'h18376,4);
TASK_PP(16'h18377,4);
TASK_PP(16'h18378,4);
TASK_PP(16'h18379,4);
TASK_PP(16'h1837A,4);
TASK_PP(16'h1837B,4);
TASK_PP(16'h1837C,4);
TASK_PP(16'h1837D,4);
TASK_PP(16'h1837E,4);
TASK_PP(16'h1837F,4);
TASK_PP(16'h18380,4);
TASK_PP(16'h18381,4);
TASK_PP(16'h18382,4);
TASK_PP(16'h18383,4);
TASK_PP(16'h18384,4);
TASK_PP(16'h18385,4);
TASK_PP(16'h18386,4);
TASK_PP(16'h18387,4);
TASK_PP(16'h18388,4);
TASK_PP(16'h18389,4);
TASK_PP(16'h1838A,4);
TASK_PP(16'h1838B,4);
TASK_PP(16'h1838C,4);
TASK_PP(16'h1838D,4);
TASK_PP(16'h1838E,4);
TASK_PP(16'h1838F,4);
TASK_PP(16'h18390,4);
TASK_PP(16'h18391,4);
TASK_PP(16'h18392,4);
TASK_PP(16'h18393,4);
TASK_PP(16'h18394,4);
TASK_PP(16'h18395,4);
TASK_PP(16'h18396,4);
TASK_PP(16'h18397,4);
TASK_PP(16'h18398,4);
TASK_PP(16'h18399,4);
TASK_PP(16'h1839A,4);
TASK_PP(16'h1839B,4);
TASK_PP(16'h1839C,4);
TASK_PP(16'h1839D,4);
TASK_PP(16'h1839E,4);
TASK_PP(16'h1839F,4);
TASK_PP(16'h183A0,4);
TASK_PP(16'h183A1,4);
TASK_PP(16'h183A2,4);
TASK_PP(16'h183A3,4);
TASK_PP(16'h183A4,4);
TASK_PP(16'h183A5,4);
TASK_PP(16'h183A6,4);
TASK_PP(16'h183A7,4);
TASK_PP(16'h183A8,4);
TASK_PP(16'h183A9,4);
TASK_PP(16'h183AA,4);
TASK_PP(16'h183AB,4);
TASK_PP(16'h183AC,4);
TASK_PP(16'h183AD,4);
TASK_PP(16'h183AE,4);
TASK_PP(16'h183AF,4);
TASK_PP(16'h183B0,4);
TASK_PP(16'h183B1,4);
TASK_PP(16'h183B2,4);
TASK_PP(16'h183B3,4);
TASK_PP(16'h183B4,4);
TASK_PP(16'h183B5,4);
TASK_PP(16'h183B6,4);
TASK_PP(16'h183B7,4);
TASK_PP(16'h183B8,4);
TASK_PP(16'h183B9,4);
TASK_PP(16'h183BA,4);
TASK_PP(16'h183BB,4);
TASK_PP(16'h183BC,4);
TASK_PP(16'h183BD,4);
TASK_PP(16'h183BE,4);
TASK_PP(16'h183BF,4);
TASK_PP(16'h183C0,4);
TASK_PP(16'h183C1,4);
TASK_PP(16'h183C2,4);
TASK_PP(16'h183C3,4);
TASK_PP(16'h183C4,4);
TASK_PP(16'h183C5,4);
TASK_PP(16'h183C6,4);
TASK_PP(16'h183C7,4);
TASK_PP(16'h183C8,4);
TASK_PP(16'h183C9,4);
TASK_PP(16'h183CA,4);
TASK_PP(16'h183CB,4);
TASK_PP(16'h183CC,4);
TASK_PP(16'h183CD,4);
TASK_PP(16'h183CE,4);
TASK_PP(16'h183CF,4);
TASK_PP(16'h183D0,4);
TASK_PP(16'h183D1,4);
TASK_PP(16'h183D2,4);
TASK_PP(16'h183D3,4);
TASK_PP(16'h183D4,4);
TASK_PP(16'h183D5,4);
TASK_PP(16'h183D6,4);
TASK_PP(16'h183D7,4);
TASK_PP(16'h183D8,4);
TASK_PP(16'h183D9,4);
TASK_PP(16'h183DA,4);
TASK_PP(16'h183DB,4);
TASK_PP(16'h183DC,4);
TASK_PP(16'h183DD,4);
TASK_PP(16'h183DE,4);
TASK_PP(16'h183DF,4);
TASK_PP(16'h183E0,4);
TASK_PP(16'h183E1,4);
TASK_PP(16'h183E2,4);
TASK_PP(16'h183E3,4);
TASK_PP(16'h183E4,4);
TASK_PP(16'h183E5,4);
TASK_PP(16'h183E6,4);
TASK_PP(16'h183E7,4);
TASK_PP(16'h183E8,4);
TASK_PP(16'h183E9,4);
TASK_PP(16'h183EA,4);
TASK_PP(16'h183EB,4);
TASK_PP(16'h183EC,4);
TASK_PP(16'h183ED,4);
TASK_PP(16'h183EE,4);
TASK_PP(16'h183EF,4);
TASK_PP(16'h183F0,4);
TASK_PP(16'h183F1,4);
TASK_PP(16'h183F2,4);
TASK_PP(16'h183F3,4);
TASK_PP(16'h183F4,4);
TASK_PP(16'h183F5,4);
TASK_PP(16'h183F6,4);
TASK_PP(16'h183F7,4);
TASK_PP(16'h183F8,4);
TASK_PP(16'h183F9,4);
TASK_PP(16'h183FA,4);
TASK_PP(16'h183FB,4);
TASK_PP(16'h183FC,4);
TASK_PP(16'h183FD,4);
TASK_PP(16'h183FE,4);
TASK_PP(16'h183FF,4);
TASK_PP(16'h18400,4);
TASK_PP(16'h18401,4);
TASK_PP(16'h18402,4);
TASK_PP(16'h18403,4);
TASK_PP(16'h18404,4);
TASK_PP(16'h18405,4);
TASK_PP(16'h18406,4);
TASK_PP(16'h18407,4);
TASK_PP(16'h18408,4);
TASK_PP(16'h18409,4);
TASK_PP(16'h1840A,4);
TASK_PP(16'h1840B,4);
TASK_PP(16'h1840C,4);
TASK_PP(16'h1840D,4);
TASK_PP(16'h1840E,4);
TASK_PP(16'h1840F,4);
TASK_PP(16'h18410,4);
TASK_PP(16'h18411,4);
TASK_PP(16'h18412,4);
TASK_PP(16'h18413,4);
TASK_PP(16'h18414,4);
TASK_PP(16'h18415,4);
TASK_PP(16'h18416,4);
TASK_PP(16'h18417,4);
TASK_PP(16'h18418,4);
TASK_PP(16'h18419,4);
TASK_PP(16'h1841A,4);
TASK_PP(16'h1841B,4);
TASK_PP(16'h1841C,4);
TASK_PP(16'h1841D,4);
TASK_PP(16'h1841E,4);
TASK_PP(16'h1841F,4);
TASK_PP(16'h18420,4);
TASK_PP(16'h18421,4);
TASK_PP(16'h18422,4);
TASK_PP(16'h18423,4);
TASK_PP(16'h18424,4);
TASK_PP(16'h18425,4);
TASK_PP(16'h18426,4);
TASK_PP(16'h18427,4);
TASK_PP(16'h18428,4);
TASK_PP(16'h18429,4);
TASK_PP(16'h1842A,4);
TASK_PP(16'h1842B,4);
TASK_PP(16'h1842C,4);
TASK_PP(16'h1842D,4);
TASK_PP(16'h1842E,4);
TASK_PP(16'h1842F,4);
TASK_PP(16'h18430,4);
TASK_PP(16'h18431,4);
TASK_PP(16'h18432,4);
TASK_PP(16'h18433,4);
TASK_PP(16'h18434,4);
TASK_PP(16'h18435,4);
TASK_PP(16'h18436,4);
TASK_PP(16'h18437,4);
TASK_PP(16'h18438,4);
TASK_PP(16'h18439,4);
TASK_PP(16'h1843A,4);
TASK_PP(16'h1843B,4);
TASK_PP(16'h1843C,4);
TASK_PP(16'h1843D,4);
TASK_PP(16'h1843E,4);
TASK_PP(16'h1843F,4);
TASK_PP(16'h18440,4);
TASK_PP(16'h18441,4);
TASK_PP(16'h18442,4);
TASK_PP(16'h18443,4);
TASK_PP(16'h18444,4);
TASK_PP(16'h18445,4);
TASK_PP(16'h18446,4);
TASK_PP(16'h18447,4);
TASK_PP(16'h18448,4);
TASK_PP(16'h18449,4);
TASK_PP(16'h1844A,4);
TASK_PP(16'h1844B,4);
TASK_PP(16'h1844C,4);
TASK_PP(16'h1844D,4);
TASK_PP(16'h1844E,4);
TASK_PP(16'h1844F,4);
TASK_PP(16'h18450,4);
TASK_PP(16'h18451,4);
TASK_PP(16'h18452,4);
TASK_PP(16'h18453,4);
TASK_PP(16'h18454,4);
TASK_PP(16'h18455,4);
TASK_PP(16'h18456,4);
TASK_PP(16'h18457,4);
TASK_PP(16'h18458,4);
TASK_PP(16'h18459,4);
TASK_PP(16'h1845A,4);
TASK_PP(16'h1845B,4);
TASK_PP(16'h1845C,4);
TASK_PP(16'h1845D,4);
TASK_PP(16'h1845E,4);
TASK_PP(16'h1845F,4);
TASK_PP(16'h18460,4);
TASK_PP(16'h18461,4);
TASK_PP(16'h18462,4);
TASK_PP(16'h18463,4);
TASK_PP(16'h18464,4);
TASK_PP(16'h18465,4);
TASK_PP(16'h18466,4);
TASK_PP(16'h18467,4);
TASK_PP(16'h18468,4);
TASK_PP(16'h18469,4);
TASK_PP(16'h1846A,4);
TASK_PP(16'h1846B,4);
TASK_PP(16'h1846C,4);
TASK_PP(16'h1846D,4);
TASK_PP(16'h1846E,4);
TASK_PP(16'h1846F,4);
TASK_PP(16'h18470,4);
TASK_PP(16'h18471,4);
TASK_PP(16'h18472,4);
TASK_PP(16'h18473,4);
TASK_PP(16'h18474,4);
TASK_PP(16'h18475,4);
TASK_PP(16'h18476,4);
TASK_PP(16'h18477,4);
TASK_PP(16'h18478,4);
TASK_PP(16'h18479,4);
TASK_PP(16'h1847A,4);
TASK_PP(16'h1847B,4);
TASK_PP(16'h1847C,4);
TASK_PP(16'h1847D,4);
TASK_PP(16'h1847E,4);
TASK_PP(16'h1847F,4);
TASK_PP(16'h18480,4);
TASK_PP(16'h18481,4);
TASK_PP(16'h18482,4);
TASK_PP(16'h18483,4);
TASK_PP(16'h18484,4);
TASK_PP(16'h18485,4);
TASK_PP(16'h18486,4);
TASK_PP(16'h18487,4);
TASK_PP(16'h18488,4);
TASK_PP(16'h18489,4);
TASK_PP(16'h1848A,4);
TASK_PP(16'h1848B,4);
TASK_PP(16'h1848C,4);
TASK_PP(16'h1848D,4);
TASK_PP(16'h1848E,4);
TASK_PP(16'h1848F,4);
TASK_PP(16'h18490,4);
TASK_PP(16'h18491,4);
TASK_PP(16'h18492,4);
TASK_PP(16'h18493,4);
TASK_PP(16'h18494,4);
TASK_PP(16'h18495,4);
TASK_PP(16'h18496,4);
TASK_PP(16'h18497,4);
TASK_PP(16'h18498,4);
TASK_PP(16'h18499,4);
TASK_PP(16'h1849A,4);
TASK_PP(16'h1849B,4);
TASK_PP(16'h1849C,4);
TASK_PP(16'h1849D,4);
TASK_PP(16'h1849E,4);
TASK_PP(16'h1849F,4);
TASK_PP(16'h184A0,4);
TASK_PP(16'h184A1,4);
TASK_PP(16'h184A2,4);
TASK_PP(16'h184A3,4);
TASK_PP(16'h184A4,4);
TASK_PP(16'h184A5,4);
TASK_PP(16'h184A6,4);
TASK_PP(16'h184A7,4);
TASK_PP(16'h184A8,4);
TASK_PP(16'h184A9,4);
TASK_PP(16'h184AA,4);
TASK_PP(16'h184AB,4);
TASK_PP(16'h184AC,4);
TASK_PP(16'h184AD,4);
TASK_PP(16'h184AE,4);
TASK_PP(16'h184AF,4);
TASK_PP(16'h184B0,4);
TASK_PP(16'h184B1,4);
TASK_PP(16'h184B2,4);
TASK_PP(16'h184B3,4);
TASK_PP(16'h184B4,4);
TASK_PP(16'h184B5,4);
TASK_PP(16'h184B6,4);
TASK_PP(16'h184B7,4);
TASK_PP(16'h184B8,4);
TASK_PP(16'h184B9,4);
TASK_PP(16'h184BA,4);
TASK_PP(16'h184BB,4);
TASK_PP(16'h184BC,4);
TASK_PP(16'h184BD,4);
TASK_PP(16'h184BE,4);
TASK_PP(16'h184BF,4);
TASK_PP(16'h184C0,4);
TASK_PP(16'h184C1,4);
TASK_PP(16'h184C2,4);
TASK_PP(16'h184C3,4);
TASK_PP(16'h184C4,4);
TASK_PP(16'h184C5,4);
TASK_PP(16'h184C6,4);
TASK_PP(16'h184C7,4);
TASK_PP(16'h184C8,4);
TASK_PP(16'h184C9,4);
TASK_PP(16'h184CA,4);
TASK_PP(16'h184CB,4);
TASK_PP(16'h184CC,4);
TASK_PP(16'h184CD,4);
TASK_PP(16'h184CE,4);
TASK_PP(16'h184CF,4);
TASK_PP(16'h184D0,4);
TASK_PP(16'h184D1,4);
TASK_PP(16'h184D2,4);
TASK_PP(16'h184D3,4);
TASK_PP(16'h184D4,4);
TASK_PP(16'h184D5,4);
TASK_PP(16'h184D6,4);
TASK_PP(16'h184D7,4);
TASK_PP(16'h184D8,4);
TASK_PP(16'h184D9,4);
TASK_PP(16'h184DA,4);
TASK_PP(16'h184DB,4);
TASK_PP(16'h184DC,4);
TASK_PP(16'h184DD,4);
TASK_PP(16'h184DE,4);
TASK_PP(16'h184DF,4);
TASK_PP(16'h184E0,4);
TASK_PP(16'h184E1,4);
TASK_PP(16'h184E2,4);
TASK_PP(16'h184E3,4);
TASK_PP(16'h184E4,4);
TASK_PP(16'h184E5,4);
TASK_PP(16'h184E6,4);
TASK_PP(16'h184E7,4);
TASK_PP(16'h184E8,4);
TASK_PP(16'h184E9,4);
TASK_PP(16'h184EA,4);
TASK_PP(16'h184EB,4);
TASK_PP(16'h184EC,4);
TASK_PP(16'h184ED,4);
TASK_PP(16'h184EE,4);
TASK_PP(16'h184EF,4);
TASK_PP(16'h184F0,4);
TASK_PP(16'h184F1,4);
TASK_PP(16'h184F2,4);
TASK_PP(16'h184F3,4);
TASK_PP(16'h184F4,4);
TASK_PP(16'h184F5,4);
TASK_PP(16'h184F6,4);
TASK_PP(16'h184F7,4);
TASK_PP(16'h184F8,4);
TASK_PP(16'h184F9,4);
TASK_PP(16'h184FA,4);
TASK_PP(16'h184FB,4);
TASK_PP(16'h184FC,4);
TASK_PP(16'h184FD,4);
TASK_PP(16'h184FE,4);
TASK_PP(16'h184FF,4);
TASK_PP(16'h18500,4);
TASK_PP(16'h18501,4);
TASK_PP(16'h18502,4);
TASK_PP(16'h18503,4);
TASK_PP(16'h18504,4);
TASK_PP(16'h18505,4);
TASK_PP(16'h18506,4);
TASK_PP(16'h18507,4);
TASK_PP(16'h18508,4);
TASK_PP(16'h18509,4);
TASK_PP(16'h1850A,4);
TASK_PP(16'h1850B,4);
TASK_PP(16'h1850C,4);
TASK_PP(16'h1850D,4);
TASK_PP(16'h1850E,4);
TASK_PP(16'h1850F,4);
TASK_PP(16'h18510,4);
TASK_PP(16'h18511,4);
TASK_PP(16'h18512,4);
TASK_PP(16'h18513,4);
TASK_PP(16'h18514,4);
TASK_PP(16'h18515,4);
TASK_PP(16'h18516,4);
TASK_PP(16'h18517,4);
TASK_PP(16'h18518,4);
TASK_PP(16'h18519,4);
TASK_PP(16'h1851A,4);
TASK_PP(16'h1851B,4);
TASK_PP(16'h1851C,4);
TASK_PP(16'h1851D,4);
TASK_PP(16'h1851E,4);
TASK_PP(16'h1851F,4);
TASK_PP(16'h18520,4);
TASK_PP(16'h18521,4);
TASK_PP(16'h18522,4);
TASK_PP(16'h18523,4);
TASK_PP(16'h18524,4);
TASK_PP(16'h18525,4);
TASK_PP(16'h18526,4);
TASK_PP(16'h18527,4);
TASK_PP(16'h18528,4);
TASK_PP(16'h18529,4);
TASK_PP(16'h1852A,4);
TASK_PP(16'h1852B,4);
TASK_PP(16'h1852C,4);
TASK_PP(16'h1852D,4);
TASK_PP(16'h1852E,4);
TASK_PP(16'h1852F,4);
TASK_PP(16'h18530,4);
TASK_PP(16'h18531,4);
TASK_PP(16'h18532,4);
TASK_PP(16'h18533,4);
TASK_PP(16'h18534,4);
TASK_PP(16'h18535,4);
TASK_PP(16'h18536,4);
TASK_PP(16'h18537,4);
TASK_PP(16'h18538,4);
TASK_PP(16'h18539,4);
TASK_PP(16'h1853A,4);
TASK_PP(16'h1853B,4);
TASK_PP(16'h1853C,4);
TASK_PP(16'h1853D,4);
TASK_PP(16'h1853E,4);
TASK_PP(16'h1853F,4);
TASK_PP(16'h18540,4);
TASK_PP(16'h18541,4);
TASK_PP(16'h18542,4);
TASK_PP(16'h18543,4);
TASK_PP(16'h18544,4);
TASK_PP(16'h18545,4);
TASK_PP(16'h18546,4);
TASK_PP(16'h18547,4);
TASK_PP(16'h18548,4);
TASK_PP(16'h18549,4);
TASK_PP(16'h1854A,4);
TASK_PP(16'h1854B,4);
TASK_PP(16'h1854C,4);
TASK_PP(16'h1854D,4);
TASK_PP(16'h1854E,4);
TASK_PP(16'h1854F,4);
TASK_PP(16'h18550,4);
TASK_PP(16'h18551,4);
TASK_PP(16'h18552,4);
TASK_PP(16'h18553,4);
TASK_PP(16'h18554,4);
TASK_PP(16'h18555,4);
TASK_PP(16'h18556,4);
TASK_PP(16'h18557,4);
TASK_PP(16'h18558,4);
TASK_PP(16'h18559,4);
TASK_PP(16'h1855A,4);
TASK_PP(16'h1855B,4);
TASK_PP(16'h1855C,4);
TASK_PP(16'h1855D,4);
TASK_PP(16'h1855E,4);
TASK_PP(16'h1855F,4);
TASK_PP(16'h18560,4);
TASK_PP(16'h18561,4);
TASK_PP(16'h18562,4);
TASK_PP(16'h18563,4);
TASK_PP(16'h18564,4);
TASK_PP(16'h18565,4);
TASK_PP(16'h18566,4);
TASK_PP(16'h18567,4);
TASK_PP(16'h18568,4);
TASK_PP(16'h18569,4);
TASK_PP(16'h1856A,4);
TASK_PP(16'h1856B,4);
TASK_PP(16'h1856C,4);
TASK_PP(16'h1856D,4);
TASK_PP(16'h1856E,4);
TASK_PP(16'h1856F,4);
TASK_PP(16'h18570,4);
TASK_PP(16'h18571,4);
TASK_PP(16'h18572,4);
TASK_PP(16'h18573,4);
TASK_PP(16'h18574,4);
TASK_PP(16'h18575,4);
TASK_PP(16'h18576,4);
TASK_PP(16'h18577,4);
TASK_PP(16'h18578,4);
TASK_PP(16'h18579,4);
TASK_PP(16'h1857A,4);
TASK_PP(16'h1857B,4);
TASK_PP(16'h1857C,4);
TASK_PP(16'h1857D,4);
TASK_PP(16'h1857E,4);
TASK_PP(16'h1857F,4);
TASK_PP(16'h18580,4);
TASK_PP(16'h18581,4);
TASK_PP(16'h18582,4);
TASK_PP(16'h18583,4);
TASK_PP(16'h18584,4);
TASK_PP(16'h18585,4);
TASK_PP(16'h18586,4);
TASK_PP(16'h18587,4);
TASK_PP(16'h18588,4);
TASK_PP(16'h18589,4);
TASK_PP(16'h1858A,4);
TASK_PP(16'h1858B,4);
TASK_PP(16'h1858C,4);
TASK_PP(16'h1858D,4);
TASK_PP(16'h1858E,4);
TASK_PP(16'h1858F,4);
TASK_PP(16'h18590,4);
TASK_PP(16'h18591,4);
TASK_PP(16'h18592,4);
TASK_PP(16'h18593,4);
TASK_PP(16'h18594,4);
TASK_PP(16'h18595,4);
TASK_PP(16'h18596,4);
TASK_PP(16'h18597,4);
TASK_PP(16'h18598,4);
TASK_PP(16'h18599,4);
TASK_PP(16'h1859A,4);
TASK_PP(16'h1859B,4);
TASK_PP(16'h1859C,4);
TASK_PP(16'h1859D,4);
TASK_PP(16'h1859E,4);
TASK_PP(16'h1859F,4);
TASK_PP(16'h185A0,4);
TASK_PP(16'h185A1,4);
TASK_PP(16'h185A2,4);
TASK_PP(16'h185A3,4);
TASK_PP(16'h185A4,4);
TASK_PP(16'h185A5,4);
TASK_PP(16'h185A6,4);
TASK_PP(16'h185A7,4);
TASK_PP(16'h185A8,4);
TASK_PP(16'h185A9,4);
TASK_PP(16'h185AA,4);
TASK_PP(16'h185AB,4);
TASK_PP(16'h185AC,4);
TASK_PP(16'h185AD,4);
TASK_PP(16'h185AE,4);
TASK_PP(16'h185AF,4);
TASK_PP(16'h185B0,4);
TASK_PP(16'h185B1,4);
TASK_PP(16'h185B2,4);
TASK_PP(16'h185B3,4);
TASK_PP(16'h185B4,4);
TASK_PP(16'h185B5,4);
TASK_PP(16'h185B6,4);
TASK_PP(16'h185B7,4);
TASK_PP(16'h185B8,4);
TASK_PP(16'h185B9,4);
TASK_PP(16'h185BA,4);
TASK_PP(16'h185BB,4);
TASK_PP(16'h185BC,4);
TASK_PP(16'h185BD,4);
TASK_PP(16'h185BE,4);
TASK_PP(16'h185BF,4);
TASK_PP(16'h185C0,4);
TASK_PP(16'h185C1,4);
TASK_PP(16'h185C2,4);
TASK_PP(16'h185C3,4);
TASK_PP(16'h185C4,4);
TASK_PP(16'h185C5,4);
TASK_PP(16'h185C6,4);
TASK_PP(16'h185C7,4);
TASK_PP(16'h185C8,4);
TASK_PP(16'h185C9,4);
TASK_PP(16'h185CA,4);
TASK_PP(16'h185CB,4);
TASK_PP(16'h185CC,4);
TASK_PP(16'h185CD,4);
TASK_PP(16'h185CE,4);
TASK_PP(16'h185CF,4);
TASK_PP(16'h185D0,4);
TASK_PP(16'h185D1,4);
TASK_PP(16'h185D2,4);
TASK_PP(16'h185D3,4);
TASK_PP(16'h185D4,4);
TASK_PP(16'h185D5,4);
TASK_PP(16'h185D6,4);
TASK_PP(16'h185D7,4);
TASK_PP(16'h185D8,4);
TASK_PP(16'h185D9,4);
TASK_PP(16'h185DA,4);
TASK_PP(16'h185DB,4);
TASK_PP(16'h185DC,4);
TASK_PP(16'h185DD,4);
TASK_PP(16'h185DE,4);
TASK_PP(16'h185DF,4);
TASK_PP(16'h185E0,4);
TASK_PP(16'h185E1,4);
TASK_PP(16'h185E2,4);
TASK_PP(16'h185E3,4);
TASK_PP(16'h185E4,4);
TASK_PP(16'h185E5,4);
TASK_PP(16'h185E6,4);
TASK_PP(16'h185E7,4);
TASK_PP(16'h185E8,4);
TASK_PP(16'h185E9,4);
TASK_PP(16'h185EA,4);
TASK_PP(16'h185EB,4);
TASK_PP(16'h185EC,4);
TASK_PP(16'h185ED,4);
TASK_PP(16'h185EE,4);
TASK_PP(16'h185EF,4);
TASK_PP(16'h185F0,4);
TASK_PP(16'h185F1,4);
TASK_PP(16'h185F2,4);
TASK_PP(16'h185F3,4);
TASK_PP(16'h185F4,4);
TASK_PP(16'h185F5,4);
TASK_PP(16'h185F6,4);
TASK_PP(16'h185F7,4);
TASK_PP(16'h185F8,4);
TASK_PP(16'h185F9,4);
TASK_PP(16'h185FA,4);
TASK_PP(16'h185FB,4);
TASK_PP(16'h185FC,4);
TASK_PP(16'h185FD,4);
TASK_PP(16'h185FE,4);
TASK_PP(16'h185FF,4);
TASK_PP(16'h18600,4);
TASK_PP(16'h18601,4);
TASK_PP(16'h18602,4);
TASK_PP(16'h18603,4);
TASK_PP(16'h18604,4);
TASK_PP(16'h18605,4);
TASK_PP(16'h18606,4);
TASK_PP(16'h18607,4);
TASK_PP(16'h18608,4);
TASK_PP(16'h18609,4);
TASK_PP(16'h1860A,4);
TASK_PP(16'h1860B,4);
TASK_PP(16'h1860C,4);
TASK_PP(16'h1860D,4);
TASK_PP(16'h1860E,4);
TASK_PP(16'h1860F,4);
TASK_PP(16'h18610,4);
TASK_PP(16'h18611,4);
TASK_PP(16'h18612,4);
TASK_PP(16'h18613,4);
TASK_PP(16'h18614,4);
TASK_PP(16'h18615,4);
TASK_PP(16'h18616,4);
TASK_PP(16'h18617,4);
TASK_PP(16'h18618,4);
TASK_PP(16'h18619,4);
TASK_PP(16'h1861A,4);
TASK_PP(16'h1861B,4);
TASK_PP(16'h1861C,4);
TASK_PP(16'h1861D,4);
TASK_PP(16'h1861E,4);
TASK_PP(16'h1861F,4);
TASK_PP(16'h18620,4);
TASK_PP(16'h18621,4);
TASK_PP(16'h18622,4);
TASK_PP(16'h18623,4);
TASK_PP(16'h18624,4);
TASK_PP(16'h18625,4);
TASK_PP(16'h18626,4);
TASK_PP(16'h18627,4);
TASK_PP(16'h18628,4);
TASK_PP(16'h18629,4);
TASK_PP(16'h1862A,4);
TASK_PP(16'h1862B,4);
TASK_PP(16'h1862C,4);
TASK_PP(16'h1862D,4);
TASK_PP(16'h1862E,4);
TASK_PP(16'h1862F,4);
TASK_PP(16'h18630,4);
TASK_PP(16'h18631,4);
TASK_PP(16'h18632,4);
TASK_PP(16'h18633,4);
TASK_PP(16'h18634,4);
TASK_PP(16'h18635,4);
TASK_PP(16'h18636,4);
TASK_PP(16'h18637,4);
TASK_PP(16'h18638,4);
TASK_PP(16'h18639,4);
TASK_PP(16'h1863A,4);
TASK_PP(16'h1863B,4);
TASK_PP(16'h1863C,4);
TASK_PP(16'h1863D,4);
TASK_PP(16'h1863E,4);
TASK_PP(16'h1863F,4);
TASK_PP(16'h18640,4);
TASK_PP(16'h18641,4);
TASK_PP(16'h18642,4);
TASK_PP(16'h18643,4);
TASK_PP(16'h18644,4);
TASK_PP(16'h18645,4);
TASK_PP(16'h18646,4);
TASK_PP(16'h18647,4);
TASK_PP(16'h18648,4);
TASK_PP(16'h18649,4);
TASK_PP(16'h1864A,4);
TASK_PP(16'h1864B,4);
TASK_PP(16'h1864C,4);
TASK_PP(16'h1864D,4);
TASK_PP(16'h1864E,4);
TASK_PP(16'h1864F,4);
TASK_PP(16'h18650,4);
TASK_PP(16'h18651,4);
TASK_PP(16'h18652,4);
TASK_PP(16'h18653,4);
TASK_PP(16'h18654,4);
TASK_PP(16'h18655,4);
TASK_PP(16'h18656,4);
TASK_PP(16'h18657,4);
TASK_PP(16'h18658,4);
TASK_PP(16'h18659,4);
TASK_PP(16'h1865A,4);
TASK_PP(16'h1865B,4);
TASK_PP(16'h1865C,4);
TASK_PP(16'h1865D,4);
TASK_PP(16'h1865E,4);
TASK_PP(16'h1865F,4);
TASK_PP(16'h18660,4);
TASK_PP(16'h18661,4);
TASK_PP(16'h18662,4);
TASK_PP(16'h18663,4);
TASK_PP(16'h18664,4);
TASK_PP(16'h18665,4);
TASK_PP(16'h18666,4);
TASK_PP(16'h18667,4);
TASK_PP(16'h18668,4);
TASK_PP(16'h18669,4);
TASK_PP(16'h1866A,4);
TASK_PP(16'h1866B,4);
TASK_PP(16'h1866C,4);
TASK_PP(16'h1866D,4);
TASK_PP(16'h1866E,4);
TASK_PP(16'h1866F,4);
TASK_PP(16'h18670,4);
TASK_PP(16'h18671,4);
TASK_PP(16'h18672,4);
TASK_PP(16'h18673,4);
TASK_PP(16'h18674,4);
TASK_PP(16'h18675,4);
TASK_PP(16'h18676,4);
TASK_PP(16'h18677,4);
TASK_PP(16'h18678,4);
TASK_PP(16'h18679,4);
TASK_PP(16'h1867A,4);
TASK_PP(16'h1867B,4);
TASK_PP(16'h1867C,4);
TASK_PP(16'h1867D,4);
TASK_PP(16'h1867E,4);
TASK_PP(16'h1867F,4);
TASK_PP(16'h18680,4);
TASK_PP(16'h18681,4);
TASK_PP(16'h18682,4);
TASK_PP(16'h18683,4);
TASK_PP(16'h18684,4);
TASK_PP(16'h18685,4);
TASK_PP(16'h18686,4);
TASK_PP(16'h18687,4);
TASK_PP(16'h18688,4);
TASK_PP(16'h18689,4);
TASK_PP(16'h1868A,4);
TASK_PP(16'h1868B,4);
TASK_PP(16'h1868C,4);
TASK_PP(16'h1868D,4);
TASK_PP(16'h1868E,4);
TASK_PP(16'h1868F,4);
TASK_PP(16'h18690,4);
TASK_PP(16'h18691,4);
TASK_PP(16'h18692,4);
TASK_PP(16'h18693,4);
TASK_PP(16'h18694,4);
TASK_PP(16'h18695,4);
TASK_PP(16'h18696,4);
TASK_PP(16'h18697,4);
TASK_PP(16'h18698,4);
TASK_PP(16'h18699,4);
TASK_PP(16'h1869A,4);
TASK_PP(16'h1869B,4);
TASK_PP(16'h1869C,4);
TASK_PP(16'h1869D,4);
TASK_PP(16'h1869E,4);
TASK_PP(16'h1869F,4);
TASK_PP(16'h186A0,4);
TASK_PP(16'h186A1,4);
TASK_PP(16'h186A2,4);
TASK_PP(16'h186A3,4);
TASK_PP(16'h186A4,4);
TASK_PP(16'h186A5,4);
TASK_PP(16'h186A6,4);
TASK_PP(16'h186A7,4);
TASK_PP(16'h186A8,4);
TASK_PP(16'h186A9,4);
TASK_PP(16'h186AA,4);
TASK_PP(16'h186AB,4);
TASK_PP(16'h186AC,4);
TASK_PP(16'h186AD,4);
TASK_PP(16'h186AE,4);
TASK_PP(16'h186AF,4);
TASK_PP(16'h186B0,4);
TASK_PP(16'h186B1,4);
TASK_PP(16'h186B2,4);
TASK_PP(16'h186B3,4);
TASK_PP(16'h186B4,4);
TASK_PP(16'h186B5,4);
TASK_PP(16'h186B6,4);
TASK_PP(16'h186B7,4);
TASK_PP(16'h186B8,4);
TASK_PP(16'h186B9,4);
TASK_PP(16'h186BA,4);
TASK_PP(16'h186BB,4);
TASK_PP(16'h186BC,4);
TASK_PP(16'h186BD,4);
TASK_PP(16'h186BE,4);
TASK_PP(16'h186BF,4);
TASK_PP(16'h186C0,4);
TASK_PP(16'h186C1,4);
TASK_PP(16'h186C2,4);
TASK_PP(16'h186C3,4);
TASK_PP(16'h186C4,4);
TASK_PP(16'h186C5,4);
TASK_PP(16'h186C6,4);
TASK_PP(16'h186C7,4);
TASK_PP(16'h186C8,4);
TASK_PP(16'h186C9,4);
TASK_PP(16'h186CA,4);
TASK_PP(16'h186CB,4);
TASK_PP(16'h186CC,4);
TASK_PP(16'h186CD,4);
TASK_PP(16'h186CE,4);
TASK_PP(16'h186CF,4);
TASK_PP(16'h186D0,4);
TASK_PP(16'h186D1,4);
TASK_PP(16'h186D2,4);
TASK_PP(16'h186D3,4);
TASK_PP(16'h186D4,4);
TASK_PP(16'h186D5,4);
TASK_PP(16'h186D6,4);
TASK_PP(16'h186D7,4);
TASK_PP(16'h186D8,4);
TASK_PP(16'h186D9,4);
TASK_PP(16'h186DA,4);
TASK_PP(16'h186DB,4);
TASK_PP(16'h186DC,4);
TASK_PP(16'h186DD,4);
TASK_PP(16'h186DE,4);
TASK_PP(16'h186DF,4);
TASK_PP(16'h186E0,4);
TASK_PP(16'h186E1,4);
TASK_PP(16'h186E2,4);
TASK_PP(16'h186E3,4);
TASK_PP(16'h186E4,4);
TASK_PP(16'h186E5,4);
TASK_PP(16'h186E6,4);
TASK_PP(16'h186E7,4);
TASK_PP(16'h186E8,4);
TASK_PP(16'h186E9,4);
TASK_PP(16'h186EA,4);
TASK_PP(16'h186EB,4);
TASK_PP(16'h186EC,4);
TASK_PP(16'h186ED,4);
TASK_PP(16'h186EE,4);
TASK_PP(16'h186EF,4);
TASK_PP(16'h186F0,4);
TASK_PP(16'h186F1,4);
TASK_PP(16'h186F2,4);
TASK_PP(16'h186F3,4);
TASK_PP(16'h186F4,4);
TASK_PP(16'h186F5,4);
TASK_PP(16'h186F6,4);
TASK_PP(16'h186F7,4);
TASK_PP(16'h186F8,4);
TASK_PP(16'h186F9,4);
TASK_PP(16'h186FA,4);
TASK_PP(16'h186FB,4);
TASK_PP(16'h186FC,4);
TASK_PP(16'h186FD,4);
TASK_PP(16'h186FE,4);
TASK_PP(16'h186FF,4);
TASK_PP(16'h18700,4);
TASK_PP(16'h18701,4);
TASK_PP(16'h18702,4);
TASK_PP(16'h18703,4);
TASK_PP(16'h18704,4);
TASK_PP(16'h18705,4);
TASK_PP(16'h18706,4);
TASK_PP(16'h18707,4);
TASK_PP(16'h18708,4);
TASK_PP(16'h18709,4);
TASK_PP(16'h1870A,4);
TASK_PP(16'h1870B,4);
TASK_PP(16'h1870C,4);
TASK_PP(16'h1870D,4);
TASK_PP(16'h1870E,4);
TASK_PP(16'h1870F,4);
TASK_PP(16'h18710,4);
TASK_PP(16'h18711,4);
TASK_PP(16'h18712,4);
TASK_PP(16'h18713,4);
TASK_PP(16'h18714,4);
TASK_PP(16'h18715,4);
TASK_PP(16'h18716,4);
TASK_PP(16'h18717,4);
TASK_PP(16'h18718,4);
TASK_PP(16'h18719,4);
TASK_PP(16'h1871A,4);
TASK_PP(16'h1871B,4);
TASK_PP(16'h1871C,4);
TASK_PP(16'h1871D,4);
TASK_PP(16'h1871E,4);
TASK_PP(16'h1871F,4);
TASK_PP(16'h18720,4);
TASK_PP(16'h18721,4);
TASK_PP(16'h18722,4);
TASK_PP(16'h18723,4);
TASK_PP(16'h18724,4);
TASK_PP(16'h18725,4);
TASK_PP(16'h18726,4);
TASK_PP(16'h18727,4);
TASK_PP(16'h18728,4);
TASK_PP(16'h18729,4);
TASK_PP(16'h1872A,4);
TASK_PP(16'h1872B,4);
TASK_PP(16'h1872C,4);
TASK_PP(16'h1872D,4);
TASK_PP(16'h1872E,4);
TASK_PP(16'h1872F,4);
TASK_PP(16'h18730,4);
TASK_PP(16'h18731,4);
TASK_PP(16'h18732,4);
TASK_PP(16'h18733,4);
TASK_PP(16'h18734,4);
TASK_PP(16'h18735,4);
TASK_PP(16'h18736,4);
TASK_PP(16'h18737,4);
TASK_PP(16'h18738,4);
TASK_PP(16'h18739,4);
TASK_PP(16'h1873A,4);
TASK_PP(16'h1873B,4);
TASK_PP(16'h1873C,4);
TASK_PP(16'h1873D,4);
TASK_PP(16'h1873E,4);
TASK_PP(16'h1873F,4);
TASK_PP(16'h18740,4);
TASK_PP(16'h18741,4);
TASK_PP(16'h18742,4);
TASK_PP(16'h18743,4);
TASK_PP(16'h18744,4);
TASK_PP(16'h18745,4);
TASK_PP(16'h18746,4);
TASK_PP(16'h18747,4);
TASK_PP(16'h18748,4);
TASK_PP(16'h18749,4);
TASK_PP(16'h1874A,4);
TASK_PP(16'h1874B,4);
TASK_PP(16'h1874C,4);
TASK_PP(16'h1874D,4);
TASK_PP(16'h1874E,4);
TASK_PP(16'h1874F,4);
TASK_PP(16'h18750,4);
TASK_PP(16'h18751,4);
TASK_PP(16'h18752,4);
TASK_PP(16'h18753,4);
TASK_PP(16'h18754,4);
TASK_PP(16'h18755,4);
TASK_PP(16'h18756,4);
TASK_PP(16'h18757,4);
TASK_PP(16'h18758,4);
TASK_PP(16'h18759,4);
TASK_PP(16'h1875A,4);
TASK_PP(16'h1875B,4);
TASK_PP(16'h1875C,4);
TASK_PP(16'h1875D,4);
TASK_PP(16'h1875E,4);
TASK_PP(16'h1875F,4);
TASK_PP(16'h18760,4);
TASK_PP(16'h18761,4);
TASK_PP(16'h18762,4);
TASK_PP(16'h18763,4);
TASK_PP(16'h18764,4);
TASK_PP(16'h18765,4);
TASK_PP(16'h18766,4);
TASK_PP(16'h18767,4);
TASK_PP(16'h18768,4);
TASK_PP(16'h18769,4);
TASK_PP(16'h1876A,4);
TASK_PP(16'h1876B,4);
TASK_PP(16'h1876C,4);
TASK_PP(16'h1876D,4);
TASK_PP(16'h1876E,4);
TASK_PP(16'h1876F,4);
TASK_PP(16'h18770,4);
TASK_PP(16'h18771,4);
TASK_PP(16'h18772,4);
TASK_PP(16'h18773,4);
TASK_PP(16'h18774,4);
TASK_PP(16'h18775,4);
TASK_PP(16'h18776,4);
TASK_PP(16'h18777,4);
TASK_PP(16'h18778,4);
TASK_PP(16'h18779,4);
TASK_PP(16'h1877A,4);
TASK_PP(16'h1877B,4);
TASK_PP(16'h1877C,4);
TASK_PP(16'h1877D,4);
TASK_PP(16'h1877E,4);
TASK_PP(16'h1877F,4);
TASK_PP(16'h18780,4);
TASK_PP(16'h18781,4);
TASK_PP(16'h18782,4);
TASK_PP(16'h18783,4);
TASK_PP(16'h18784,4);
TASK_PP(16'h18785,4);
TASK_PP(16'h18786,4);
TASK_PP(16'h18787,4);
TASK_PP(16'h18788,4);
TASK_PP(16'h18789,4);
TASK_PP(16'h1878A,4);
TASK_PP(16'h1878B,4);
TASK_PP(16'h1878C,4);
TASK_PP(16'h1878D,4);
TASK_PP(16'h1878E,4);
TASK_PP(16'h1878F,4);
TASK_PP(16'h18790,4);
TASK_PP(16'h18791,4);
TASK_PP(16'h18792,4);
TASK_PP(16'h18793,4);
TASK_PP(16'h18794,4);
TASK_PP(16'h18795,4);
TASK_PP(16'h18796,4);
TASK_PP(16'h18797,4);
TASK_PP(16'h18798,4);
TASK_PP(16'h18799,4);
TASK_PP(16'h1879A,4);
TASK_PP(16'h1879B,4);
TASK_PP(16'h1879C,4);
TASK_PP(16'h1879D,4);
TASK_PP(16'h1879E,4);
TASK_PP(16'h1879F,4);
TASK_PP(16'h187A0,4);
TASK_PP(16'h187A1,4);
TASK_PP(16'h187A2,4);
TASK_PP(16'h187A3,4);
TASK_PP(16'h187A4,4);
TASK_PP(16'h187A5,4);
TASK_PP(16'h187A6,4);
TASK_PP(16'h187A7,4);
TASK_PP(16'h187A8,4);
TASK_PP(16'h187A9,4);
TASK_PP(16'h187AA,4);
TASK_PP(16'h187AB,4);
TASK_PP(16'h187AC,4);
TASK_PP(16'h187AD,4);
TASK_PP(16'h187AE,4);
TASK_PP(16'h187AF,4);
TASK_PP(16'h187B0,4);
TASK_PP(16'h187B1,4);
TASK_PP(16'h187B2,4);
TASK_PP(16'h187B3,4);
TASK_PP(16'h187B4,4);
TASK_PP(16'h187B5,4);
TASK_PP(16'h187B6,4);
TASK_PP(16'h187B7,4);
TASK_PP(16'h187B8,4);
TASK_PP(16'h187B9,4);
TASK_PP(16'h187BA,4);
TASK_PP(16'h187BB,4);
TASK_PP(16'h187BC,4);
TASK_PP(16'h187BD,4);
TASK_PP(16'h187BE,4);
TASK_PP(16'h187BF,4);
TASK_PP(16'h187C0,4);
TASK_PP(16'h187C1,4);
TASK_PP(16'h187C2,4);
TASK_PP(16'h187C3,4);
TASK_PP(16'h187C4,4);
TASK_PP(16'h187C5,4);
TASK_PP(16'h187C6,4);
TASK_PP(16'h187C7,4);
TASK_PP(16'h187C8,4);
TASK_PP(16'h187C9,4);
TASK_PP(16'h187CA,4);
TASK_PP(16'h187CB,4);
TASK_PP(16'h187CC,4);
TASK_PP(16'h187CD,4);
TASK_PP(16'h187CE,4);
TASK_PP(16'h187CF,4);
TASK_PP(16'h187D0,4);
TASK_PP(16'h187D1,4);
TASK_PP(16'h187D2,4);
TASK_PP(16'h187D3,4);
TASK_PP(16'h187D4,4);
TASK_PP(16'h187D5,4);
TASK_PP(16'h187D6,4);
TASK_PP(16'h187D7,4);
TASK_PP(16'h187D8,4);
TASK_PP(16'h187D9,4);
TASK_PP(16'h187DA,4);
TASK_PP(16'h187DB,4);
TASK_PP(16'h187DC,4);
TASK_PP(16'h187DD,4);
TASK_PP(16'h187DE,4);
TASK_PP(16'h187DF,4);
TASK_PP(16'h187E0,4);
TASK_PP(16'h187E1,4);
TASK_PP(16'h187E2,4);
TASK_PP(16'h187E3,4);
TASK_PP(16'h187E4,4);
TASK_PP(16'h187E5,4);
TASK_PP(16'h187E6,4);
TASK_PP(16'h187E7,4);
TASK_PP(16'h187E8,4);
TASK_PP(16'h187E9,4);
TASK_PP(16'h187EA,4);
TASK_PP(16'h187EB,4);
TASK_PP(16'h187EC,4);
TASK_PP(16'h187ED,4);
TASK_PP(16'h187EE,4);
TASK_PP(16'h187EF,4);
TASK_PP(16'h187F0,4);
TASK_PP(16'h187F1,4);
TASK_PP(16'h187F2,4);
TASK_PP(16'h187F3,4);
TASK_PP(16'h187F4,4);
TASK_PP(16'h187F5,4);
TASK_PP(16'h187F6,4);
TASK_PP(16'h187F7,4);
TASK_PP(16'h187F8,4);
TASK_PP(16'h187F9,4);
TASK_PP(16'h187FA,4);
TASK_PP(16'h187FB,4);
TASK_PP(16'h187FC,4);
TASK_PP(16'h187FD,4);
TASK_PP(16'h187FE,4);
TASK_PP(16'h187FF,4);
TASK_PP(16'h18800,4);
TASK_PP(16'h18801,4);
TASK_PP(16'h18802,4);
TASK_PP(16'h18803,4);
TASK_PP(16'h18804,4);
TASK_PP(16'h18805,4);
TASK_PP(16'h18806,4);
TASK_PP(16'h18807,4);
TASK_PP(16'h18808,4);
TASK_PP(16'h18809,4);
TASK_PP(16'h1880A,4);
TASK_PP(16'h1880B,4);
TASK_PP(16'h1880C,4);
TASK_PP(16'h1880D,4);
TASK_PP(16'h1880E,4);
TASK_PP(16'h1880F,4);
TASK_PP(16'h18810,4);
TASK_PP(16'h18811,4);
TASK_PP(16'h18812,4);
TASK_PP(16'h18813,4);
TASK_PP(16'h18814,4);
TASK_PP(16'h18815,4);
TASK_PP(16'h18816,4);
TASK_PP(16'h18817,4);
TASK_PP(16'h18818,4);
TASK_PP(16'h18819,4);
TASK_PP(16'h1881A,4);
TASK_PP(16'h1881B,4);
TASK_PP(16'h1881C,4);
TASK_PP(16'h1881D,4);
TASK_PP(16'h1881E,4);
TASK_PP(16'h1881F,4);
TASK_PP(16'h18820,4);
TASK_PP(16'h18821,4);
TASK_PP(16'h18822,4);
TASK_PP(16'h18823,4);
TASK_PP(16'h18824,4);
TASK_PP(16'h18825,4);
TASK_PP(16'h18826,4);
TASK_PP(16'h18827,4);
TASK_PP(16'h18828,4);
TASK_PP(16'h18829,4);
TASK_PP(16'h1882A,4);
TASK_PP(16'h1882B,4);
TASK_PP(16'h1882C,4);
TASK_PP(16'h1882D,4);
TASK_PP(16'h1882E,4);
TASK_PP(16'h1882F,4);
TASK_PP(16'h18830,4);
TASK_PP(16'h18831,4);
TASK_PP(16'h18832,4);
TASK_PP(16'h18833,4);
TASK_PP(16'h18834,4);
TASK_PP(16'h18835,4);
TASK_PP(16'h18836,4);
TASK_PP(16'h18837,4);
TASK_PP(16'h18838,4);
TASK_PP(16'h18839,4);
TASK_PP(16'h1883A,4);
TASK_PP(16'h1883B,4);
TASK_PP(16'h1883C,4);
TASK_PP(16'h1883D,4);
TASK_PP(16'h1883E,4);
TASK_PP(16'h1883F,4);
TASK_PP(16'h18840,4);
TASK_PP(16'h18841,4);
TASK_PP(16'h18842,4);
TASK_PP(16'h18843,4);
TASK_PP(16'h18844,4);
TASK_PP(16'h18845,4);
TASK_PP(16'h18846,4);
TASK_PP(16'h18847,4);
TASK_PP(16'h18848,4);
TASK_PP(16'h18849,4);
TASK_PP(16'h1884A,4);
TASK_PP(16'h1884B,4);
TASK_PP(16'h1884C,4);
TASK_PP(16'h1884D,4);
TASK_PP(16'h1884E,4);
TASK_PP(16'h1884F,4);
TASK_PP(16'h18850,4);
TASK_PP(16'h18851,4);
TASK_PP(16'h18852,4);
TASK_PP(16'h18853,4);
TASK_PP(16'h18854,4);
TASK_PP(16'h18855,4);
TASK_PP(16'h18856,4);
TASK_PP(16'h18857,4);
TASK_PP(16'h18858,4);
TASK_PP(16'h18859,4);
TASK_PP(16'h1885A,4);
TASK_PP(16'h1885B,4);
TASK_PP(16'h1885C,4);
TASK_PP(16'h1885D,4);
TASK_PP(16'h1885E,4);
TASK_PP(16'h1885F,4);
TASK_PP(16'h18860,4);
TASK_PP(16'h18861,4);
TASK_PP(16'h18862,4);
TASK_PP(16'h18863,4);
TASK_PP(16'h18864,4);
TASK_PP(16'h18865,4);
TASK_PP(16'h18866,4);
TASK_PP(16'h18867,4);
TASK_PP(16'h18868,4);
TASK_PP(16'h18869,4);
TASK_PP(16'h1886A,4);
TASK_PP(16'h1886B,4);
TASK_PP(16'h1886C,4);
TASK_PP(16'h1886D,4);
TASK_PP(16'h1886E,4);
TASK_PP(16'h1886F,4);
TASK_PP(16'h18870,4);
TASK_PP(16'h18871,4);
TASK_PP(16'h18872,4);
TASK_PP(16'h18873,4);
TASK_PP(16'h18874,4);
TASK_PP(16'h18875,4);
TASK_PP(16'h18876,4);
TASK_PP(16'h18877,4);
TASK_PP(16'h18878,4);
TASK_PP(16'h18879,4);
TASK_PP(16'h1887A,4);
TASK_PP(16'h1887B,4);
TASK_PP(16'h1887C,4);
TASK_PP(16'h1887D,4);
TASK_PP(16'h1887E,4);
TASK_PP(16'h1887F,4);
TASK_PP(16'h18880,4);
TASK_PP(16'h18881,4);
TASK_PP(16'h18882,4);
TASK_PP(16'h18883,4);
TASK_PP(16'h18884,4);
TASK_PP(16'h18885,4);
TASK_PP(16'h18886,4);
TASK_PP(16'h18887,4);
TASK_PP(16'h18888,4);
TASK_PP(16'h18889,4);
TASK_PP(16'h1888A,4);
TASK_PP(16'h1888B,4);
TASK_PP(16'h1888C,4);
TASK_PP(16'h1888D,4);
TASK_PP(16'h1888E,4);
TASK_PP(16'h1888F,4);
TASK_PP(16'h18890,4);
TASK_PP(16'h18891,4);
TASK_PP(16'h18892,4);
TASK_PP(16'h18893,4);
TASK_PP(16'h18894,4);
TASK_PP(16'h18895,4);
TASK_PP(16'h18896,4);
TASK_PP(16'h18897,4);
TASK_PP(16'h18898,4);
TASK_PP(16'h18899,4);
TASK_PP(16'h1889A,4);
TASK_PP(16'h1889B,4);
TASK_PP(16'h1889C,4);
TASK_PP(16'h1889D,4);
TASK_PP(16'h1889E,4);
TASK_PP(16'h1889F,4);
TASK_PP(16'h188A0,4);
TASK_PP(16'h188A1,4);
TASK_PP(16'h188A2,4);
TASK_PP(16'h188A3,4);
TASK_PP(16'h188A4,4);
TASK_PP(16'h188A5,4);
TASK_PP(16'h188A6,4);
TASK_PP(16'h188A7,4);
TASK_PP(16'h188A8,4);
TASK_PP(16'h188A9,4);
TASK_PP(16'h188AA,4);
TASK_PP(16'h188AB,4);
TASK_PP(16'h188AC,4);
TASK_PP(16'h188AD,4);
TASK_PP(16'h188AE,4);
TASK_PP(16'h188AF,4);
TASK_PP(16'h188B0,4);
TASK_PP(16'h188B1,4);
TASK_PP(16'h188B2,4);
TASK_PP(16'h188B3,4);
TASK_PP(16'h188B4,4);
TASK_PP(16'h188B5,4);
TASK_PP(16'h188B6,4);
TASK_PP(16'h188B7,4);
TASK_PP(16'h188B8,4);
TASK_PP(16'h188B9,4);
TASK_PP(16'h188BA,4);
TASK_PP(16'h188BB,4);
TASK_PP(16'h188BC,4);
TASK_PP(16'h188BD,4);
TASK_PP(16'h188BE,4);
TASK_PP(16'h188BF,4);
TASK_PP(16'h188C0,4);
TASK_PP(16'h188C1,4);
TASK_PP(16'h188C2,4);
TASK_PP(16'h188C3,4);
TASK_PP(16'h188C4,4);
TASK_PP(16'h188C5,4);
TASK_PP(16'h188C6,4);
TASK_PP(16'h188C7,4);
TASK_PP(16'h188C8,4);
TASK_PP(16'h188C9,4);
TASK_PP(16'h188CA,4);
TASK_PP(16'h188CB,4);
TASK_PP(16'h188CC,4);
TASK_PP(16'h188CD,4);
TASK_PP(16'h188CE,4);
TASK_PP(16'h188CF,4);
TASK_PP(16'h188D0,4);
TASK_PP(16'h188D1,4);
TASK_PP(16'h188D2,4);
TASK_PP(16'h188D3,4);
TASK_PP(16'h188D4,4);
TASK_PP(16'h188D5,4);
TASK_PP(16'h188D6,4);
TASK_PP(16'h188D7,4);
TASK_PP(16'h188D8,4);
TASK_PP(16'h188D9,4);
TASK_PP(16'h188DA,4);
TASK_PP(16'h188DB,4);
TASK_PP(16'h188DC,4);
TASK_PP(16'h188DD,4);
TASK_PP(16'h188DE,4);
TASK_PP(16'h188DF,4);
TASK_PP(16'h188E0,4);
TASK_PP(16'h188E1,4);
TASK_PP(16'h188E2,4);
TASK_PP(16'h188E3,4);
TASK_PP(16'h188E4,4);
TASK_PP(16'h188E5,4);
TASK_PP(16'h188E6,4);
TASK_PP(16'h188E7,4);
TASK_PP(16'h188E8,4);
TASK_PP(16'h188E9,4);
TASK_PP(16'h188EA,4);
TASK_PP(16'h188EB,4);
TASK_PP(16'h188EC,4);
TASK_PP(16'h188ED,4);
TASK_PP(16'h188EE,4);
TASK_PP(16'h188EF,4);
TASK_PP(16'h188F0,4);
TASK_PP(16'h188F1,4);
TASK_PP(16'h188F2,4);
TASK_PP(16'h188F3,4);
TASK_PP(16'h188F4,4);
TASK_PP(16'h188F5,4);
TASK_PP(16'h188F6,4);
TASK_PP(16'h188F7,4);
TASK_PP(16'h188F8,4);
TASK_PP(16'h188F9,4);
TASK_PP(16'h188FA,4);
TASK_PP(16'h188FB,4);
TASK_PP(16'h188FC,4);
TASK_PP(16'h188FD,4);
TASK_PP(16'h188FE,4);
TASK_PP(16'h188FF,4);
TASK_PP(16'h18900,4);
TASK_PP(16'h18901,4);
TASK_PP(16'h18902,4);
TASK_PP(16'h18903,4);
TASK_PP(16'h18904,4);
TASK_PP(16'h18905,4);
TASK_PP(16'h18906,4);
TASK_PP(16'h18907,4);
TASK_PP(16'h18908,4);
TASK_PP(16'h18909,4);
TASK_PP(16'h1890A,4);
TASK_PP(16'h1890B,4);
TASK_PP(16'h1890C,4);
TASK_PP(16'h1890D,4);
TASK_PP(16'h1890E,4);
TASK_PP(16'h1890F,4);
TASK_PP(16'h18910,4);
TASK_PP(16'h18911,4);
TASK_PP(16'h18912,4);
TASK_PP(16'h18913,4);
TASK_PP(16'h18914,4);
TASK_PP(16'h18915,4);
TASK_PP(16'h18916,4);
TASK_PP(16'h18917,4);
TASK_PP(16'h18918,4);
TASK_PP(16'h18919,4);
TASK_PP(16'h1891A,4);
TASK_PP(16'h1891B,4);
TASK_PP(16'h1891C,4);
TASK_PP(16'h1891D,4);
TASK_PP(16'h1891E,4);
TASK_PP(16'h1891F,4);
TASK_PP(16'h18920,4);
TASK_PP(16'h18921,4);
TASK_PP(16'h18922,4);
TASK_PP(16'h18923,4);
TASK_PP(16'h18924,4);
TASK_PP(16'h18925,4);
TASK_PP(16'h18926,4);
TASK_PP(16'h18927,4);
TASK_PP(16'h18928,4);
TASK_PP(16'h18929,4);
TASK_PP(16'h1892A,4);
TASK_PP(16'h1892B,4);
TASK_PP(16'h1892C,4);
TASK_PP(16'h1892D,4);
TASK_PP(16'h1892E,4);
TASK_PP(16'h1892F,4);
TASK_PP(16'h18930,4);
TASK_PP(16'h18931,4);
TASK_PP(16'h18932,4);
TASK_PP(16'h18933,4);
TASK_PP(16'h18934,4);
TASK_PP(16'h18935,4);
TASK_PP(16'h18936,4);
TASK_PP(16'h18937,4);
TASK_PP(16'h18938,4);
TASK_PP(16'h18939,4);
TASK_PP(16'h1893A,4);
TASK_PP(16'h1893B,4);
TASK_PP(16'h1893C,4);
TASK_PP(16'h1893D,4);
TASK_PP(16'h1893E,4);
TASK_PP(16'h1893F,4);
TASK_PP(16'h18940,4);
TASK_PP(16'h18941,4);
TASK_PP(16'h18942,4);
TASK_PP(16'h18943,4);
TASK_PP(16'h18944,4);
TASK_PP(16'h18945,4);
TASK_PP(16'h18946,4);
TASK_PP(16'h18947,4);
TASK_PP(16'h18948,4);
TASK_PP(16'h18949,4);
TASK_PP(16'h1894A,4);
TASK_PP(16'h1894B,4);
TASK_PP(16'h1894C,4);
TASK_PP(16'h1894D,4);
TASK_PP(16'h1894E,4);
TASK_PP(16'h1894F,4);
TASK_PP(16'h18950,4);
TASK_PP(16'h18951,4);
TASK_PP(16'h18952,4);
TASK_PP(16'h18953,4);
TASK_PP(16'h18954,4);
TASK_PP(16'h18955,4);
TASK_PP(16'h18956,4);
TASK_PP(16'h18957,4);
TASK_PP(16'h18958,4);
TASK_PP(16'h18959,4);
TASK_PP(16'h1895A,4);
TASK_PP(16'h1895B,4);
TASK_PP(16'h1895C,4);
TASK_PP(16'h1895D,4);
TASK_PP(16'h1895E,4);
TASK_PP(16'h1895F,4);
TASK_PP(16'h18960,4);
TASK_PP(16'h18961,4);
TASK_PP(16'h18962,4);
TASK_PP(16'h18963,4);
TASK_PP(16'h18964,4);
TASK_PP(16'h18965,4);
TASK_PP(16'h18966,4);
TASK_PP(16'h18967,4);
TASK_PP(16'h18968,4);
TASK_PP(16'h18969,4);
TASK_PP(16'h1896A,4);
TASK_PP(16'h1896B,4);
TASK_PP(16'h1896C,4);
TASK_PP(16'h1896D,4);
TASK_PP(16'h1896E,4);
TASK_PP(16'h1896F,4);
TASK_PP(16'h18970,4);
TASK_PP(16'h18971,4);
TASK_PP(16'h18972,4);
TASK_PP(16'h18973,4);
TASK_PP(16'h18974,4);
TASK_PP(16'h18975,4);
TASK_PP(16'h18976,4);
TASK_PP(16'h18977,4);
TASK_PP(16'h18978,4);
TASK_PP(16'h18979,4);
TASK_PP(16'h1897A,4);
TASK_PP(16'h1897B,4);
TASK_PP(16'h1897C,4);
TASK_PP(16'h1897D,4);
TASK_PP(16'h1897E,4);
TASK_PP(16'h1897F,4);
TASK_PP(16'h18980,4);
TASK_PP(16'h18981,4);
TASK_PP(16'h18982,4);
TASK_PP(16'h18983,4);
TASK_PP(16'h18984,4);
TASK_PP(16'h18985,4);
TASK_PP(16'h18986,4);
TASK_PP(16'h18987,4);
TASK_PP(16'h18988,4);
TASK_PP(16'h18989,4);
TASK_PP(16'h1898A,4);
TASK_PP(16'h1898B,4);
TASK_PP(16'h1898C,4);
TASK_PP(16'h1898D,4);
TASK_PP(16'h1898E,4);
TASK_PP(16'h1898F,4);
TASK_PP(16'h18990,4);
TASK_PP(16'h18991,4);
TASK_PP(16'h18992,4);
TASK_PP(16'h18993,4);
TASK_PP(16'h18994,4);
TASK_PP(16'h18995,4);
TASK_PP(16'h18996,4);
TASK_PP(16'h18997,4);
TASK_PP(16'h18998,4);
TASK_PP(16'h18999,4);
TASK_PP(16'h1899A,4);
TASK_PP(16'h1899B,4);
TASK_PP(16'h1899C,4);
TASK_PP(16'h1899D,4);
TASK_PP(16'h1899E,4);
TASK_PP(16'h1899F,4);
TASK_PP(16'h189A0,4);
TASK_PP(16'h189A1,4);
TASK_PP(16'h189A2,4);
TASK_PP(16'h189A3,4);
TASK_PP(16'h189A4,4);
TASK_PP(16'h189A5,4);
TASK_PP(16'h189A6,4);
TASK_PP(16'h189A7,4);
TASK_PP(16'h189A8,4);
TASK_PP(16'h189A9,4);
TASK_PP(16'h189AA,4);
TASK_PP(16'h189AB,4);
TASK_PP(16'h189AC,4);
TASK_PP(16'h189AD,4);
TASK_PP(16'h189AE,4);
TASK_PP(16'h189AF,4);
TASK_PP(16'h189B0,4);
TASK_PP(16'h189B1,4);
TASK_PP(16'h189B2,4);
TASK_PP(16'h189B3,4);
TASK_PP(16'h189B4,4);
TASK_PP(16'h189B5,4);
TASK_PP(16'h189B6,4);
TASK_PP(16'h189B7,4);
TASK_PP(16'h189B8,4);
TASK_PP(16'h189B9,4);
TASK_PP(16'h189BA,4);
TASK_PP(16'h189BB,4);
TASK_PP(16'h189BC,4);
TASK_PP(16'h189BD,4);
TASK_PP(16'h189BE,4);
TASK_PP(16'h189BF,4);
TASK_PP(16'h189C0,4);
TASK_PP(16'h189C1,4);
TASK_PP(16'h189C2,4);
TASK_PP(16'h189C3,4);
TASK_PP(16'h189C4,4);
TASK_PP(16'h189C5,4);
TASK_PP(16'h189C6,4);
TASK_PP(16'h189C7,4);
TASK_PP(16'h189C8,4);
TASK_PP(16'h189C9,4);
TASK_PP(16'h189CA,4);
TASK_PP(16'h189CB,4);
TASK_PP(16'h189CC,4);
TASK_PP(16'h189CD,4);
TASK_PP(16'h189CE,4);
TASK_PP(16'h189CF,4);
TASK_PP(16'h189D0,4);
TASK_PP(16'h189D1,4);
TASK_PP(16'h189D2,4);
TASK_PP(16'h189D3,4);
TASK_PP(16'h189D4,4);
TASK_PP(16'h189D5,4);
TASK_PP(16'h189D6,4);
TASK_PP(16'h189D7,4);
TASK_PP(16'h189D8,4);
TASK_PP(16'h189D9,4);
TASK_PP(16'h189DA,4);
TASK_PP(16'h189DB,4);
TASK_PP(16'h189DC,4);
TASK_PP(16'h189DD,4);
TASK_PP(16'h189DE,4);
TASK_PP(16'h189DF,4);
TASK_PP(16'h189E0,4);
TASK_PP(16'h189E1,4);
TASK_PP(16'h189E2,4);
TASK_PP(16'h189E3,4);
TASK_PP(16'h189E4,4);
TASK_PP(16'h189E5,4);
TASK_PP(16'h189E6,4);
TASK_PP(16'h189E7,4);
TASK_PP(16'h189E8,4);
TASK_PP(16'h189E9,4);
TASK_PP(16'h189EA,4);
TASK_PP(16'h189EB,4);
TASK_PP(16'h189EC,4);
TASK_PP(16'h189ED,4);
TASK_PP(16'h189EE,4);
TASK_PP(16'h189EF,4);
TASK_PP(16'h189F0,4);
TASK_PP(16'h189F1,4);
TASK_PP(16'h189F2,4);
TASK_PP(16'h189F3,4);
TASK_PP(16'h189F4,4);
TASK_PP(16'h189F5,4);
TASK_PP(16'h189F6,4);
TASK_PP(16'h189F7,4);
TASK_PP(16'h189F8,4);
TASK_PP(16'h189F9,4);
TASK_PP(16'h189FA,4);
TASK_PP(16'h189FB,4);
TASK_PP(16'h189FC,4);
TASK_PP(16'h189FD,4);
TASK_PP(16'h189FE,4);
TASK_PP(16'h189FF,4);
TASK_PP(16'h18A00,4);
TASK_PP(16'h18A01,4);
TASK_PP(16'h18A02,4);
TASK_PP(16'h18A03,4);
TASK_PP(16'h18A04,4);
TASK_PP(16'h18A05,4);
TASK_PP(16'h18A06,4);
TASK_PP(16'h18A07,4);
TASK_PP(16'h18A08,4);
TASK_PP(16'h18A09,4);
TASK_PP(16'h18A0A,4);
TASK_PP(16'h18A0B,4);
TASK_PP(16'h18A0C,4);
TASK_PP(16'h18A0D,4);
TASK_PP(16'h18A0E,4);
TASK_PP(16'h18A0F,4);
TASK_PP(16'h18A10,4);
TASK_PP(16'h18A11,4);
TASK_PP(16'h18A12,4);
TASK_PP(16'h18A13,4);
TASK_PP(16'h18A14,4);
TASK_PP(16'h18A15,4);
TASK_PP(16'h18A16,4);
TASK_PP(16'h18A17,4);
TASK_PP(16'h18A18,4);
TASK_PP(16'h18A19,4);
TASK_PP(16'h18A1A,4);
TASK_PP(16'h18A1B,4);
TASK_PP(16'h18A1C,4);
TASK_PP(16'h18A1D,4);
TASK_PP(16'h18A1E,4);
TASK_PP(16'h18A1F,4);
TASK_PP(16'h18A20,4);
TASK_PP(16'h18A21,4);
TASK_PP(16'h18A22,4);
TASK_PP(16'h18A23,4);
TASK_PP(16'h18A24,4);
TASK_PP(16'h18A25,4);
TASK_PP(16'h18A26,4);
TASK_PP(16'h18A27,4);
TASK_PP(16'h18A28,4);
TASK_PP(16'h18A29,4);
TASK_PP(16'h18A2A,4);
TASK_PP(16'h18A2B,4);
TASK_PP(16'h18A2C,4);
TASK_PP(16'h18A2D,4);
TASK_PP(16'h18A2E,4);
TASK_PP(16'h18A2F,4);
TASK_PP(16'h18A30,4);
TASK_PP(16'h18A31,4);
TASK_PP(16'h18A32,4);
TASK_PP(16'h18A33,4);
TASK_PP(16'h18A34,4);
TASK_PP(16'h18A35,4);
TASK_PP(16'h18A36,4);
TASK_PP(16'h18A37,4);
TASK_PP(16'h18A38,4);
TASK_PP(16'h18A39,4);
TASK_PP(16'h18A3A,4);
TASK_PP(16'h18A3B,4);
TASK_PP(16'h18A3C,4);
TASK_PP(16'h18A3D,4);
TASK_PP(16'h18A3E,4);
TASK_PP(16'h18A3F,4);
TASK_PP(16'h18A40,4);
TASK_PP(16'h18A41,4);
TASK_PP(16'h18A42,4);
TASK_PP(16'h18A43,4);
TASK_PP(16'h18A44,4);
TASK_PP(16'h18A45,4);
TASK_PP(16'h18A46,4);
TASK_PP(16'h18A47,4);
TASK_PP(16'h18A48,4);
TASK_PP(16'h18A49,4);
TASK_PP(16'h18A4A,4);
TASK_PP(16'h18A4B,4);
TASK_PP(16'h18A4C,4);
TASK_PP(16'h18A4D,4);
TASK_PP(16'h18A4E,4);
TASK_PP(16'h18A4F,4);
TASK_PP(16'h18A50,4);
TASK_PP(16'h18A51,4);
TASK_PP(16'h18A52,4);
TASK_PP(16'h18A53,4);
TASK_PP(16'h18A54,4);
TASK_PP(16'h18A55,4);
TASK_PP(16'h18A56,4);
TASK_PP(16'h18A57,4);
TASK_PP(16'h18A58,4);
TASK_PP(16'h18A59,4);
TASK_PP(16'h18A5A,4);
TASK_PP(16'h18A5B,4);
TASK_PP(16'h18A5C,4);
TASK_PP(16'h18A5D,4);
TASK_PP(16'h18A5E,4);
TASK_PP(16'h18A5F,4);
TASK_PP(16'h18A60,4);
TASK_PP(16'h18A61,4);
TASK_PP(16'h18A62,4);
TASK_PP(16'h18A63,4);
TASK_PP(16'h18A64,4);
TASK_PP(16'h18A65,4);
TASK_PP(16'h18A66,4);
TASK_PP(16'h18A67,4);
TASK_PP(16'h18A68,4);
TASK_PP(16'h18A69,4);
TASK_PP(16'h18A6A,4);
TASK_PP(16'h18A6B,4);
TASK_PP(16'h18A6C,4);
TASK_PP(16'h18A6D,4);
TASK_PP(16'h18A6E,4);
TASK_PP(16'h18A6F,4);
TASK_PP(16'h18A70,4);
TASK_PP(16'h18A71,4);
TASK_PP(16'h18A72,4);
TASK_PP(16'h18A73,4);
TASK_PP(16'h18A74,4);
TASK_PP(16'h18A75,4);
TASK_PP(16'h18A76,4);
TASK_PP(16'h18A77,4);
TASK_PP(16'h18A78,4);
TASK_PP(16'h18A79,4);
TASK_PP(16'h18A7A,4);
TASK_PP(16'h18A7B,4);
TASK_PP(16'h18A7C,4);
TASK_PP(16'h18A7D,4);
TASK_PP(16'h18A7E,4);
TASK_PP(16'h18A7F,4);
TASK_PP(16'h18A80,4);
TASK_PP(16'h18A81,4);
TASK_PP(16'h18A82,4);
TASK_PP(16'h18A83,4);
TASK_PP(16'h18A84,4);
TASK_PP(16'h18A85,4);
TASK_PP(16'h18A86,4);
TASK_PP(16'h18A87,4);
TASK_PP(16'h18A88,4);
TASK_PP(16'h18A89,4);
TASK_PP(16'h18A8A,4);
TASK_PP(16'h18A8B,4);
TASK_PP(16'h18A8C,4);
TASK_PP(16'h18A8D,4);
TASK_PP(16'h18A8E,4);
TASK_PP(16'h18A8F,4);
TASK_PP(16'h18A90,4);
TASK_PP(16'h18A91,4);
TASK_PP(16'h18A92,4);
TASK_PP(16'h18A93,4);
TASK_PP(16'h18A94,4);
TASK_PP(16'h18A95,4);
TASK_PP(16'h18A96,4);
TASK_PP(16'h18A97,4);
TASK_PP(16'h18A98,4);
TASK_PP(16'h18A99,4);
TASK_PP(16'h18A9A,4);
TASK_PP(16'h18A9B,4);
TASK_PP(16'h18A9C,4);
TASK_PP(16'h18A9D,4);
TASK_PP(16'h18A9E,4);
TASK_PP(16'h18A9F,4);
TASK_PP(16'h18AA0,4);
TASK_PP(16'h18AA1,4);
TASK_PP(16'h18AA2,4);
TASK_PP(16'h18AA3,4);
TASK_PP(16'h18AA4,4);
TASK_PP(16'h18AA5,4);
TASK_PP(16'h18AA6,4);
TASK_PP(16'h18AA7,4);
TASK_PP(16'h18AA8,4);
TASK_PP(16'h18AA9,4);
TASK_PP(16'h18AAA,4);
TASK_PP(16'h18AAB,4);
TASK_PP(16'h18AAC,4);
TASK_PP(16'h18AAD,4);
TASK_PP(16'h18AAE,4);
TASK_PP(16'h18AAF,4);
TASK_PP(16'h18AB0,4);
TASK_PP(16'h18AB1,4);
TASK_PP(16'h18AB2,4);
TASK_PP(16'h18AB3,4);
TASK_PP(16'h18AB4,4);
TASK_PP(16'h18AB5,4);
TASK_PP(16'h18AB6,4);
TASK_PP(16'h18AB7,4);
TASK_PP(16'h18AB8,4);
TASK_PP(16'h18AB9,4);
TASK_PP(16'h18ABA,4);
TASK_PP(16'h18ABB,4);
TASK_PP(16'h18ABC,4);
TASK_PP(16'h18ABD,4);
TASK_PP(16'h18ABE,4);
TASK_PP(16'h18ABF,4);
TASK_PP(16'h18AC0,4);
TASK_PP(16'h18AC1,4);
TASK_PP(16'h18AC2,4);
TASK_PP(16'h18AC3,4);
TASK_PP(16'h18AC4,4);
TASK_PP(16'h18AC5,4);
TASK_PP(16'h18AC6,4);
TASK_PP(16'h18AC7,4);
TASK_PP(16'h18AC8,4);
TASK_PP(16'h18AC9,4);
TASK_PP(16'h18ACA,4);
TASK_PP(16'h18ACB,4);
TASK_PP(16'h18ACC,4);
TASK_PP(16'h18ACD,4);
TASK_PP(16'h18ACE,4);
TASK_PP(16'h18ACF,4);
TASK_PP(16'h18AD0,4);
TASK_PP(16'h18AD1,4);
TASK_PP(16'h18AD2,4);
TASK_PP(16'h18AD3,4);
TASK_PP(16'h18AD4,4);
TASK_PP(16'h18AD5,4);
TASK_PP(16'h18AD6,4);
TASK_PP(16'h18AD7,4);
TASK_PP(16'h18AD8,4);
TASK_PP(16'h18AD9,4);
TASK_PP(16'h18ADA,4);
TASK_PP(16'h18ADB,4);
TASK_PP(16'h18ADC,4);
TASK_PP(16'h18ADD,4);
TASK_PP(16'h18ADE,4);
TASK_PP(16'h18ADF,4);
TASK_PP(16'h18AE0,4);
TASK_PP(16'h18AE1,4);
TASK_PP(16'h18AE2,4);
TASK_PP(16'h18AE3,4);
TASK_PP(16'h18AE4,4);
TASK_PP(16'h18AE5,4);
TASK_PP(16'h18AE6,4);
TASK_PP(16'h18AE7,4);
TASK_PP(16'h18AE8,4);
TASK_PP(16'h18AE9,4);
TASK_PP(16'h18AEA,4);
TASK_PP(16'h18AEB,4);
TASK_PP(16'h18AEC,4);
TASK_PP(16'h18AED,4);
TASK_PP(16'h18AEE,4);
TASK_PP(16'h18AEF,4);
TASK_PP(16'h18AF0,4);
TASK_PP(16'h18AF1,4);
TASK_PP(16'h18AF2,4);
TASK_PP(16'h18AF3,4);
TASK_PP(16'h18AF4,4);
TASK_PP(16'h18AF5,4);
TASK_PP(16'h18AF6,4);
TASK_PP(16'h18AF7,4);
TASK_PP(16'h18AF8,4);
TASK_PP(16'h18AF9,4);
TASK_PP(16'h18AFA,4);
TASK_PP(16'h18AFB,4);
TASK_PP(16'h18AFC,4);
TASK_PP(16'h18AFD,4);
TASK_PP(16'h18AFE,4);
TASK_PP(16'h18AFF,4);
TASK_PP(16'h18B00,4);
TASK_PP(16'h18B01,4);
TASK_PP(16'h18B02,4);
TASK_PP(16'h18B03,4);
TASK_PP(16'h18B04,4);
TASK_PP(16'h18B05,4);
TASK_PP(16'h18B06,4);
TASK_PP(16'h18B07,4);
TASK_PP(16'h18B08,4);
TASK_PP(16'h18B09,4);
TASK_PP(16'h18B0A,4);
TASK_PP(16'h18B0B,4);
TASK_PP(16'h18B0C,4);
TASK_PP(16'h18B0D,4);
TASK_PP(16'h18B0E,4);
TASK_PP(16'h18B0F,4);
TASK_PP(16'h18B10,4);
TASK_PP(16'h18B11,4);
TASK_PP(16'h18B12,4);
TASK_PP(16'h18B13,4);
TASK_PP(16'h18B14,4);
TASK_PP(16'h18B15,4);
TASK_PP(16'h18B16,4);
TASK_PP(16'h18B17,4);
TASK_PP(16'h18B18,4);
TASK_PP(16'h18B19,4);
TASK_PP(16'h18B1A,4);
TASK_PP(16'h18B1B,4);
TASK_PP(16'h18B1C,4);
TASK_PP(16'h18B1D,4);
TASK_PP(16'h18B1E,4);
TASK_PP(16'h18B1F,4);
TASK_PP(16'h18B20,4);
TASK_PP(16'h18B21,4);
TASK_PP(16'h18B22,4);
TASK_PP(16'h18B23,4);
TASK_PP(16'h18B24,4);
TASK_PP(16'h18B25,4);
TASK_PP(16'h18B26,4);
TASK_PP(16'h18B27,4);
TASK_PP(16'h18B28,4);
TASK_PP(16'h18B29,4);
TASK_PP(16'h18B2A,4);
TASK_PP(16'h18B2B,4);
TASK_PP(16'h18B2C,4);
TASK_PP(16'h18B2D,4);
TASK_PP(16'h18B2E,4);
TASK_PP(16'h18B2F,4);
TASK_PP(16'h18B30,4);
TASK_PP(16'h18B31,4);
TASK_PP(16'h18B32,4);
TASK_PP(16'h18B33,4);
TASK_PP(16'h18B34,4);
TASK_PP(16'h18B35,4);
TASK_PP(16'h18B36,4);
TASK_PP(16'h18B37,4);
TASK_PP(16'h18B38,4);
TASK_PP(16'h18B39,4);
TASK_PP(16'h18B3A,4);
TASK_PP(16'h18B3B,4);
TASK_PP(16'h18B3C,4);
TASK_PP(16'h18B3D,4);
TASK_PP(16'h18B3E,4);
TASK_PP(16'h18B3F,4);
TASK_PP(16'h18B40,4);
TASK_PP(16'h18B41,4);
TASK_PP(16'h18B42,4);
TASK_PP(16'h18B43,4);
TASK_PP(16'h18B44,4);
TASK_PP(16'h18B45,4);
TASK_PP(16'h18B46,4);
TASK_PP(16'h18B47,4);
TASK_PP(16'h18B48,4);
TASK_PP(16'h18B49,4);
TASK_PP(16'h18B4A,4);
TASK_PP(16'h18B4B,4);
TASK_PP(16'h18B4C,4);
TASK_PP(16'h18B4D,4);
TASK_PP(16'h18B4E,4);
TASK_PP(16'h18B4F,4);
TASK_PP(16'h18B50,4);
TASK_PP(16'h18B51,4);
TASK_PP(16'h18B52,4);
TASK_PP(16'h18B53,4);
TASK_PP(16'h18B54,4);
TASK_PP(16'h18B55,4);
TASK_PP(16'h18B56,4);
TASK_PP(16'h18B57,4);
TASK_PP(16'h18B58,4);
TASK_PP(16'h18B59,4);
TASK_PP(16'h18B5A,4);
TASK_PP(16'h18B5B,4);
TASK_PP(16'h18B5C,4);
TASK_PP(16'h18B5D,4);
TASK_PP(16'h18B5E,4);
TASK_PP(16'h18B5F,4);
TASK_PP(16'h18B60,4);
TASK_PP(16'h18B61,4);
TASK_PP(16'h18B62,4);
TASK_PP(16'h18B63,4);
TASK_PP(16'h18B64,4);
TASK_PP(16'h18B65,4);
TASK_PP(16'h18B66,4);
TASK_PP(16'h18B67,4);
TASK_PP(16'h18B68,4);
TASK_PP(16'h18B69,4);
TASK_PP(16'h18B6A,4);
TASK_PP(16'h18B6B,4);
TASK_PP(16'h18B6C,4);
TASK_PP(16'h18B6D,4);
TASK_PP(16'h18B6E,4);
TASK_PP(16'h18B6F,4);
TASK_PP(16'h18B70,4);
TASK_PP(16'h18B71,4);
TASK_PP(16'h18B72,4);
TASK_PP(16'h18B73,4);
TASK_PP(16'h18B74,4);
TASK_PP(16'h18B75,4);
TASK_PP(16'h18B76,4);
TASK_PP(16'h18B77,4);
TASK_PP(16'h18B78,4);
TASK_PP(16'h18B79,4);
TASK_PP(16'h18B7A,4);
TASK_PP(16'h18B7B,4);
TASK_PP(16'h18B7C,4);
TASK_PP(16'h18B7D,4);
TASK_PP(16'h18B7E,4);
TASK_PP(16'h18B7F,4);
TASK_PP(16'h18B80,4);
TASK_PP(16'h18B81,4);
TASK_PP(16'h18B82,4);
TASK_PP(16'h18B83,4);
TASK_PP(16'h18B84,4);
TASK_PP(16'h18B85,4);
TASK_PP(16'h18B86,4);
TASK_PP(16'h18B87,4);
TASK_PP(16'h18B88,4);
TASK_PP(16'h18B89,4);
TASK_PP(16'h18B8A,4);
TASK_PP(16'h18B8B,4);
TASK_PP(16'h18B8C,4);
TASK_PP(16'h18B8D,4);
TASK_PP(16'h18B8E,4);
TASK_PP(16'h18B8F,4);
TASK_PP(16'h18B90,4);
TASK_PP(16'h18B91,4);
TASK_PP(16'h18B92,4);
TASK_PP(16'h18B93,4);
TASK_PP(16'h18B94,4);
TASK_PP(16'h18B95,4);
TASK_PP(16'h18B96,4);
TASK_PP(16'h18B97,4);
TASK_PP(16'h18B98,4);
TASK_PP(16'h18B99,4);
TASK_PP(16'h18B9A,4);
TASK_PP(16'h18B9B,4);
TASK_PP(16'h18B9C,4);
TASK_PP(16'h18B9D,4);
TASK_PP(16'h18B9E,4);
TASK_PP(16'h18B9F,4);
TASK_PP(16'h18BA0,4);
TASK_PP(16'h18BA1,4);
TASK_PP(16'h18BA2,4);
TASK_PP(16'h18BA3,4);
TASK_PP(16'h18BA4,4);
TASK_PP(16'h18BA5,4);
TASK_PP(16'h18BA6,4);
TASK_PP(16'h18BA7,4);
TASK_PP(16'h18BA8,4);
TASK_PP(16'h18BA9,4);
TASK_PP(16'h18BAA,4);
TASK_PP(16'h18BAB,4);
TASK_PP(16'h18BAC,4);
TASK_PP(16'h18BAD,4);
TASK_PP(16'h18BAE,4);
TASK_PP(16'h18BAF,4);
TASK_PP(16'h18BB0,4);
TASK_PP(16'h18BB1,4);
TASK_PP(16'h18BB2,4);
TASK_PP(16'h18BB3,4);
TASK_PP(16'h18BB4,4);
TASK_PP(16'h18BB5,4);
TASK_PP(16'h18BB6,4);
TASK_PP(16'h18BB7,4);
TASK_PP(16'h18BB8,4);
TASK_PP(16'h18BB9,4);
TASK_PP(16'h18BBA,4);
TASK_PP(16'h18BBB,4);
TASK_PP(16'h18BBC,4);
TASK_PP(16'h18BBD,4);
TASK_PP(16'h18BBE,4);
TASK_PP(16'h18BBF,4);
TASK_PP(16'h18BC0,4);
TASK_PP(16'h18BC1,4);
TASK_PP(16'h18BC2,4);
TASK_PP(16'h18BC3,4);
TASK_PP(16'h18BC4,4);
TASK_PP(16'h18BC5,4);
TASK_PP(16'h18BC6,4);
TASK_PP(16'h18BC7,4);
TASK_PP(16'h18BC8,4);
TASK_PP(16'h18BC9,4);
TASK_PP(16'h18BCA,4);
TASK_PP(16'h18BCB,4);
TASK_PP(16'h18BCC,4);
TASK_PP(16'h18BCD,4);
TASK_PP(16'h18BCE,4);
TASK_PP(16'h18BCF,4);
TASK_PP(16'h18BD0,4);
TASK_PP(16'h18BD1,4);
TASK_PP(16'h18BD2,4);
TASK_PP(16'h18BD3,4);
TASK_PP(16'h18BD4,4);
TASK_PP(16'h18BD5,4);
TASK_PP(16'h18BD6,4);
TASK_PP(16'h18BD7,4);
TASK_PP(16'h18BD8,4);
TASK_PP(16'h18BD9,4);
TASK_PP(16'h18BDA,4);
TASK_PP(16'h18BDB,4);
TASK_PP(16'h18BDC,4);
TASK_PP(16'h18BDD,4);
TASK_PP(16'h18BDE,4);
TASK_PP(16'h18BDF,4);
TASK_PP(16'h18BE0,4);
TASK_PP(16'h18BE1,4);
TASK_PP(16'h18BE2,4);
TASK_PP(16'h18BE3,4);
TASK_PP(16'h18BE4,4);
TASK_PP(16'h18BE5,4);
TASK_PP(16'h18BE6,4);
TASK_PP(16'h18BE7,4);
TASK_PP(16'h18BE8,4);
TASK_PP(16'h18BE9,4);
TASK_PP(16'h18BEA,4);
TASK_PP(16'h18BEB,4);
TASK_PP(16'h18BEC,4);
TASK_PP(16'h18BED,4);
TASK_PP(16'h18BEE,4);
TASK_PP(16'h18BEF,4);
TASK_PP(16'h18BF0,4);
TASK_PP(16'h18BF1,4);
TASK_PP(16'h18BF2,4);
TASK_PP(16'h18BF3,4);
TASK_PP(16'h18BF4,4);
TASK_PP(16'h18BF5,4);
TASK_PP(16'h18BF6,4);
TASK_PP(16'h18BF7,4);
TASK_PP(16'h18BF8,4);
TASK_PP(16'h18BF9,4);
TASK_PP(16'h18BFA,4);
TASK_PP(16'h18BFB,4);
TASK_PP(16'h18BFC,4);
TASK_PP(16'h18BFD,4);
TASK_PP(16'h18BFE,4);
TASK_PP(16'h18BFF,4);
TASK_PP(16'h18C00,4);
TASK_PP(16'h18C01,4);
TASK_PP(16'h18C02,4);
TASK_PP(16'h18C03,4);
TASK_PP(16'h18C04,4);
TASK_PP(16'h18C05,4);
TASK_PP(16'h18C06,4);
TASK_PP(16'h18C07,4);
TASK_PP(16'h18C08,4);
TASK_PP(16'h18C09,4);
TASK_PP(16'h18C0A,4);
TASK_PP(16'h18C0B,4);
TASK_PP(16'h18C0C,4);
TASK_PP(16'h18C0D,4);
TASK_PP(16'h18C0E,4);
TASK_PP(16'h18C0F,4);
TASK_PP(16'h18C10,4);
TASK_PP(16'h18C11,4);
TASK_PP(16'h18C12,4);
TASK_PP(16'h18C13,4);
TASK_PP(16'h18C14,4);
TASK_PP(16'h18C15,4);
TASK_PP(16'h18C16,4);
TASK_PP(16'h18C17,4);
TASK_PP(16'h18C18,4);
TASK_PP(16'h18C19,4);
TASK_PP(16'h18C1A,4);
TASK_PP(16'h18C1B,4);
TASK_PP(16'h18C1C,4);
TASK_PP(16'h18C1D,4);
TASK_PP(16'h18C1E,4);
TASK_PP(16'h18C1F,4);
TASK_PP(16'h18C20,4);
TASK_PP(16'h18C21,4);
TASK_PP(16'h18C22,4);
TASK_PP(16'h18C23,4);
TASK_PP(16'h18C24,4);
TASK_PP(16'h18C25,4);
TASK_PP(16'h18C26,4);
TASK_PP(16'h18C27,4);
TASK_PP(16'h18C28,4);
TASK_PP(16'h18C29,4);
TASK_PP(16'h18C2A,4);
TASK_PP(16'h18C2B,4);
TASK_PP(16'h18C2C,4);
TASK_PP(16'h18C2D,4);
TASK_PP(16'h18C2E,4);
TASK_PP(16'h18C2F,4);
TASK_PP(16'h18C30,4);
TASK_PP(16'h18C31,4);
TASK_PP(16'h18C32,4);
TASK_PP(16'h18C33,4);
TASK_PP(16'h18C34,4);
TASK_PP(16'h18C35,4);
TASK_PP(16'h18C36,4);
TASK_PP(16'h18C37,4);
TASK_PP(16'h18C38,4);
TASK_PP(16'h18C39,4);
TASK_PP(16'h18C3A,4);
TASK_PP(16'h18C3B,4);
TASK_PP(16'h18C3C,4);
TASK_PP(16'h18C3D,4);
TASK_PP(16'h18C3E,4);
TASK_PP(16'h18C3F,4);
TASK_PP(16'h18C40,4);
TASK_PP(16'h18C41,4);
TASK_PP(16'h18C42,4);
TASK_PP(16'h18C43,4);
TASK_PP(16'h18C44,4);
TASK_PP(16'h18C45,4);
TASK_PP(16'h18C46,4);
TASK_PP(16'h18C47,4);
TASK_PP(16'h18C48,4);
TASK_PP(16'h18C49,4);
TASK_PP(16'h18C4A,4);
TASK_PP(16'h18C4B,4);
TASK_PP(16'h18C4C,4);
TASK_PP(16'h18C4D,4);
TASK_PP(16'h18C4E,4);
TASK_PP(16'h18C4F,4);
TASK_PP(16'h18C50,4);
TASK_PP(16'h18C51,4);
TASK_PP(16'h18C52,4);
TASK_PP(16'h18C53,4);
TASK_PP(16'h18C54,4);
TASK_PP(16'h18C55,4);
TASK_PP(16'h18C56,4);
TASK_PP(16'h18C57,4);
TASK_PP(16'h18C58,4);
TASK_PP(16'h18C59,4);
TASK_PP(16'h18C5A,4);
TASK_PP(16'h18C5B,4);
TASK_PP(16'h18C5C,4);
TASK_PP(16'h18C5D,4);
TASK_PP(16'h18C5E,4);
TASK_PP(16'h18C5F,4);
TASK_PP(16'h18C60,4);
TASK_PP(16'h18C61,4);
TASK_PP(16'h18C62,4);
TASK_PP(16'h18C63,4);
TASK_PP(16'h18C64,4);
TASK_PP(16'h18C65,4);
TASK_PP(16'h18C66,4);
TASK_PP(16'h18C67,4);
TASK_PP(16'h18C68,4);
TASK_PP(16'h18C69,4);
TASK_PP(16'h18C6A,4);
TASK_PP(16'h18C6B,4);
TASK_PP(16'h18C6C,4);
TASK_PP(16'h18C6D,4);
TASK_PP(16'h18C6E,4);
TASK_PP(16'h18C6F,4);
TASK_PP(16'h18C70,4);
TASK_PP(16'h18C71,4);
TASK_PP(16'h18C72,4);
TASK_PP(16'h18C73,4);
TASK_PP(16'h18C74,4);
TASK_PP(16'h18C75,4);
TASK_PP(16'h18C76,4);
TASK_PP(16'h18C77,4);
TASK_PP(16'h18C78,4);
TASK_PP(16'h18C79,4);
TASK_PP(16'h18C7A,4);
TASK_PP(16'h18C7B,4);
TASK_PP(16'h18C7C,4);
TASK_PP(16'h18C7D,4);
TASK_PP(16'h18C7E,4);
TASK_PP(16'h18C7F,4);
TASK_PP(16'h18C80,4);
TASK_PP(16'h18C81,4);
TASK_PP(16'h18C82,4);
TASK_PP(16'h18C83,4);
TASK_PP(16'h18C84,4);
TASK_PP(16'h18C85,4);
TASK_PP(16'h18C86,4);
TASK_PP(16'h18C87,4);
TASK_PP(16'h18C88,4);
TASK_PP(16'h18C89,4);
TASK_PP(16'h18C8A,4);
TASK_PP(16'h18C8B,4);
TASK_PP(16'h18C8C,4);
TASK_PP(16'h18C8D,4);
TASK_PP(16'h18C8E,4);
TASK_PP(16'h18C8F,4);
TASK_PP(16'h18C90,4);
TASK_PP(16'h18C91,4);
TASK_PP(16'h18C92,4);
TASK_PP(16'h18C93,4);
TASK_PP(16'h18C94,4);
TASK_PP(16'h18C95,4);
TASK_PP(16'h18C96,4);
TASK_PP(16'h18C97,4);
TASK_PP(16'h18C98,4);
TASK_PP(16'h18C99,4);
TASK_PP(16'h18C9A,4);
TASK_PP(16'h18C9B,4);
TASK_PP(16'h18C9C,4);
TASK_PP(16'h18C9D,4);
TASK_PP(16'h18C9E,4);
TASK_PP(16'h18C9F,4);
TASK_PP(16'h18CA0,4);
TASK_PP(16'h18CA1,4);
TASK_PP(16'h18CA2,4);
TASK_PP(16'h18CA3,4);
TASK_PP(16'h18CA4,4);
TASK_PP(16'h18CA5,4);
TASK_PP(16'h18CA6,4);
TASK_PP(16'h18CA7,4);
TASK_PP(16'h18CA8,4);
TASK_PP(16'h18CA9,4);
TASK_PP(16'h18CAA,4);
TASK_PP(16'h18CAB,4);
TASK_PP(16'h18CAC,4);
TASK_PP(16'h18CAD,4);
TASK_PP(16'h18CAE,4);
TASK_PP(16'h18CAF,4);
TASK_PP(16'h18CB0,4);
TASK_PP(16'h18CB1,4);
TASK_PP(16'h18CB2,4);
TASK_PP(16'h18CB3,4);
TASK_PP(16'h18CB4,4);
TASK_PP(16'h18CB5,4);
TASK_PP(16'h18CB6,4);
TASK_PP(16'h18CB7,4);
TASK_PP(16'h18CB8,4);
TASK_PP(16'h18CB9,4);
TASK_PP(16'h18CBA,4);
TASK_PP(16'h18CBB,4);
TASK_PP(16'h18CBC,4);
TASK_PP(16'h18CBD,4);
TASK_PP(16'h18CBE,4);
TASK_PP(16'h18CBF,4);
TASK_PP(16'h18CC0,4);
TASK_PP(16'h18CC1,4);
TASK_PP(16'h18CC2,4);
TASK_PP(16'h18CC3,4);
TASK_PP(16'h18CC4,4);
TASK_PP(16'h18CC5,4);
TASK_PP(16'h18CC6,4);
TASK_PP(16'h18CC7,4);
TASK_PP(16'h18CC8,4);
TASK_PP(16'h18CC9,4);
TASK_PP(16'h18CCA,4);
TASK_PP(16'h18CCB,4);
TASK_PP(16'h18CCC,4);
TASK_PP(16'h18CCD,4);
TASK_PP(16'h18CCE,4);
TASK_PP(16'h18CCF,4);
TASK_PP(16'h18CD0,4);
TASK_PP(16'h18CD1,4);
TASK_PP(16'h18CD2,4);
TASK_PP(16'h18CD3,4);
TASK_PP(16'h18CD4,4);
TASK_PP(16'h18CD5,4);
TASK_PP(16'h18CD6,4);
TASK_PP(16'h18CD7,4);
TASK_PP(16'h18CD8,4);
TASK_PP(16'h18CD9,4);
TASK_PP(16'h18CDA,4);
TASK_PP(16'h18CDB,4);
TASK_PP(16'h18CDC,4);
TASK_PP(16'h18CDD,4);
TASK_PP(16'h18CDE,4);
TASK_PP(16'h18CDF,4);
TASK_PP(16'h18CE0,4);
TASK_PP(16'h18CE1,4);
TASK_PP(16'h18CE2,4);
TASK_PP(16'h18CE3,4);
TASK_PP(16'h18CE4,4);
TASK_PP(16'h18CE5,4);
TASK_PP(16'h18CE6,4);
TASK_PP(16'h18CE7,4);
TASK_PP(16'h18CE8,4);
TASK_PP(16'h18CE9,4);
TASK_PP(16'h18CEA,4);
TASK_PP(16'h18CEB,4);
TASK_PP(16'h18CEC,4);
TASK_PP(16'h18CED,4);
TASK_PP(16'h18CEE,4);
TASK_PP(16'h18CEF,4);
TASK_PP(16'h18CF0,4);
TASK_PP(16'h18CF1,4);
TASK_PP(16'h18CF2,4);
TASK_PP(16'h18CF3,4);
TASK_PP(16'h18CF4,4);
TASK_PP(16'h18CF5,4);
TASK_PP(16'h18CF6,4);
TASK_PP(16'h18CF7,4);
TASK_PP(16'h18CF8,4);
TASK_PP(16'h18CF9,4);
TASK_PP(16'h18CFA,4);
TASK_PP(16'h18CFB,4);
TASK_PP(16'h18CFC,4);
TASK_PP(16'h18CFD,4);
TASK_PP(16'h18CFE,4);
TASK_PP(16'h18CFF,4);
TASK_PP(16'h18D00,4);
TASK_PP(16'h18D01,4);
TASK_PP(16'h18D02,4);
TASK_PP(16'h18D03,4);
TASK_PP(16'h18D04,4);
TASK_PP(16'h18D05,4);
TASK_PP(16'h18D06,4);
TASK_PP(16'h18D07,4);
TASK_PP(16'h18D08,4);
TASK_PP(16'h18D09,4);
TASK_PP(16'h18D0A,4);
TASK_PP(16'h18D0B,4);
TASK_PP(16'h18D0C,4);
TASK_PP(16'h18D0D,4);
TASK_PP(16'h18D0E,4);
TASK_PP(16'h18D0F,4);
TASK_PP(16'h18D10,4);
TASK_PP(16'h18D11,4);
TASK_PP(16'h18D12,4);
TASK_PP(16'h18D13,4);
TASK_PP(16'h18D14,4);
TASK_PP(16'h18D15,4);
TASK_PP(16'h18D16,4);
TASK_PP(16'h18D17,4);
TASK_PP(16'h18D18,4);
TASK_PP(16'h18D19,4);
TASK_PP(16'h18D1A,4);
TASK_PP(16'h18D1B,4);
TASK_PP(16'h18D1C,4);
TASK_PP(16'h18D1D,4);
TASK_PP(16'h18D1E,4);
TASK_PP(16'h18D1F,4);
TASK_PP(16'h18D20,4);
TASK_PP(16'h18D21,4);
TASK_PP(16'h18D22,4);
TASK_PP(16'h18D23,4);
TASK_PP(16'h18D24,4);
TASK_PP(16'h18D25,4);
TASK_PP(16'h18D26,4);
TASK_PP(16'h18D27,4);
TASK_PP(16'h18D28,4);
TASK_PP(16'h18D29,4);
TASK_PP(16'h18D2A,4);
TASK_PP(16'h18D2B,4);
TASK_PP(16'h18D2C,4);
TASK_PP(16'h18D2D,4);
TASK_PP(16'h18D2E,4);
TASK_PP(16'h18D2F,4);
TASK_PP(16'h18D30,4);
TASK_PP(16'h18D31,4);
TASK_PP(16'h18D32,4);
TASK_PP(16'h18D33,4);
TASK_PP(16'h18D34,4);
TASK_PP(16'h18D35,4);
TASK_PP(16'h18D36,4);
TASK_PP(16'h18D37,4);
TASK_PP(16'h18D38,4);
TASK_PP(16'h18D39,4);
TASK_PP(16'h18D3A,4);
TASK_PP(16'h18D3B,4);
TASK_PP(16'h18D3C,4);
TASK_PP(16'h18D3D,4);
TASK_PP(16'h18D3E,4);
TASK_PP(16'h18D3F,4);
TASK_PP(16'h18D40,4);
TASK_PP(16'h18D41,4);
TASK_PP(16'h18D42,4);
TASK_PP(16'h18D43,4);
TASK_PP(16'h18D44,4);
TASK_PP(16'h18D45,4);
TASK_PP(16'h18D46,4);
TASK_PP(16'h18D47,4);
TASK_PP(16'h18D48,4);
TASK_PP(16'h18D49,4);
TASK_PP(16'h18D4A,4);
TASK_PP(16'h18D4B,4);
TASK_PP(16'h18D4C,4);
TASK_PP(16'h18D4D,4);
TASK_PP(16'h18D4E,4);
TASK_PP(16'h18D4F,4);
TASK_PP(16'h18D50,4);
TASK_PP(16'h18D51,4);
TASK_PP(16'h18D52,4);
TASK_PP(16'h18D53,4);
TASK_PP(16'h18D54,4);
TASK_PP(16'h18D55,4);
TASK_PP(16'h18D56,4);
TASK_PP(16'h18D57,4);
TASK_PP(16'h18D58,4);
TASK_PP(16'h18D59,4);
TASK_PP(16'h18D5A,4);
TASK_PP(16'h18D5B,4);
TASK_PP(16'h18D5C,4);
TASK_PP(16'h18D5D,4);
TASK_PP(16'h18D5E,4);
TASK_PP(16'h18D5F,4);
TASK_PP(16'h18D60,4);
TASK_PP(16'h18D61,4);
TASK_PP(16'h18D62,4);
TASK_PP(16'h18D63,4);
TASK_PP(16'h18D64,4);
TASK_PP(16'h18D65,4);
TASK_PP(16'h18D66,4);
TASK_PP(16'h18D67,4);
TASK_PP(16'h18D68,4);
TASK_PP(16'h18D69,4);
TASK_PP(16'h18D6A,4);
TASK_PP(16'h18D6B,4);
TASK_PP(16'h18D6C,4);
TASK_PP(16'h18D6D,4);
TASK_PP(16'h18D6E,4);
TASK_PP(16'h18D6F,4);
TASK_PP(16'h18D70,4);
TASK_PP(16'h18D71,4);
TASK_PP(16'h18D72,4);
TASK_PP(16'h18D73,4);
TASK_PP(16'h18D74,4);
TASK_PP(16'h18D75,4);
TASK_PP(16'h18D76,4);
TASK_PP(16'h18D77,4);
TASK_PP(16'h18D78,4);
TASK_PP(16'h18D79,4);
TASK_PP(16'h18D7A,4);
TASK_PP(16'h18D7B,4);
TASK_PP(16'h18D7C,4);
TASK_PP(16'h18D7D,4);
TASK_PP(16'h18D7E,4);
TASK_PP(16'h18D7F,4);
TASK_PP(16'h18D80,4);
TASK_PP(16'h18D81,4);
TASK_PP(16'h18D82,4);
TASK_PP(16'h18D83,4);
TASK_PP(16'h18D84,4);
TASK_PP(16'h18D85,4);
TASK_PP(16'h18D86,4);
TASK_PP(16'h18D87,4);
TASK_PP(16'h18D88,4);
TASK_PP(16'h18D89,4);
TASK_PP(16'h18D8A,4);
TASK_PP(16'h18D8B,4);
TASK_PP(16'h18D8C,4);
TASK_PP(16'h18D8D,4);
TASK_PP(16'h18D8E,4);
TASK_PP(16'h18D8F,4);
TASK_PP(16'h18D90,4);
TASK_PP(16'h18D91,4);
TASK_PP(16'h18D92,4);
TASK_PP(16'h18D93,4);
TASK_PP(16'h18D94,4);
TASK_PP(16'h18D95,4);
TASK_PP(16'h18D96,4);
TASK_PP(16'h18D97,4);
TASK_PP(16'h18D98,4);
TASK_PP(16'h18D99,4);
TASK_PP(16'h18D9A,4);
TASK_PP(16'h18D9B,4);
TASK_PP(16'h18D9C,4);
TASK_PP(16'h18D9D,4);
TASK_PP(16'h18D9E,4);
TASK_PP(16'h18D9F,4);
TASK_PP(16'h18DA0,4);
TASK_PP(16'h18DA1,4);
TASK_PP(16'h18DA2,4);
TASK_PP(16'h18DA3,4);
TASK_PP(16'h18DA4,4);
TASK_PP(16'h18DA5,4);
TASK_PP(16'h18DA6,4);
TASK_PP(16'h18DA7,4);
TASK_PP(16'h18DA8,4);
TASK_PP(16'h18DA9,4);
TASK_PP(16'h18DAA,4);
TASK_PP(16'h18DAB,4);
TASK_PP(16'h18DAC,4);
TASK_PP(16'h18DAD,4);
TASK_PP(16'h18DAE,4);
TASK_PP(16'h18DAF,4);
TASK_PP(16'h18DB0,4);
TASK_PP(16'h18DB1,4);
TASK_PP(16'h18DB2,4);
TASK_PP(16'h18DB3,4);
TASK_PP(16'h18DB4,4);
TASK_PP(16'h18DB5,4);
TASK_PP(16'h18DB6,4);
TASK_PP(16'h18DB7,4);
TASK_PP(16'h18DB8,4);
TASK_PP(16'h18DB9,4);
TASK_PP(16'h18DBA,4);
TASK_PP(16'h18DBB,4);
TASK_PP(16'h18DBC,4);
TASK_PP(16'h18DBD,4);
TASK_PP(16'h18DBE,4);
TASK_PP(16'h18DBF,4);
TASK_PP(16'h18DC0,4);
TASK_PP(16'h18DC1,4);
TASK_PP(16'h18DC2,4);
TASK_PP(16'h18DC3,4);
TASK_PP(16'h18DC4,4);
TASK_PP(16'h18DC5,4);
TASK_PP(16'h18DC6,4);
TASK_PP(16'h18DC7,4);
TASK_PP(16'h18DC8,4);
TASK_PP(16'h18DC9,4);
TASK_PP(16'h18DCA,4);
TASK_PP(16'h18DCB,4);
TASK_PP(16'h18DCC,4);
TASK_PP(16'h18DCD,4);
TASK_PP(16'h18DCE,4);
TASK_PP(16'h18DCF,4);
TASK_PP(16'h18DD0,4);
TASK_PP(16'h18DD1,4);
TASK_PP(16'h18DD2,4);
TASK_PP(16'h18DD3,4);
TASK_PP(16'h18DD4,4);
TASK_PP(16'h18DD5,4);
TASK_PP(16'h18DD6,4);
TASK_PP(16'h18DD7,4);
TASK_PP(16'h18DD8,4);
TASK_PP(16'h18DD9,4);
TASK_PP(16'h18DDA,4);
TASK_PP(16'h18DDB,4);
TASK_PP(16'h18DDC,4);
TASK_PP(16'h18DDD,4);
TASK_PP(16'h18DDE,4);
TASK_PP(16'h18DDF,4);
TASK_PP(16'h18DE0,4);
TASK_PP(16'h18DE1,4);
TASK_PP(16'h18DE2,4);
TASK_PP(16'h18DE3,4);
TASK_PP(16'h18DE4,4);
TASK_PP(16'h18DE5,4);
TASK_PP(16'h18DE6,4);
TASK_PP(16'h18DE7,4);
TASK_PP(16'h18DE8,4);
TASK_PP(16'h18DE9,4);
TASK_PP(16'h18DEA,4);
TASK_PP(16'h18DEB,4);
TASK_PP(16'h18DEC,4);
TASK_PP(16'h18DED,4);
TASK_PP(16'h18DEE,4);
TASK_PP(16'h18DEF,4);
TASK_PP(16'h18DF0,4);
TASK_PP(16'h18DF1,4);
TASK_PP(16'h18DF2,4);
TASK_PP(16'h18DF3,4);
TASK_PP(16'h18DF4,4);
TASK_PP(16'h18DF5,4);
TASK_PP(16'h18DF6,4);
TASK_PP(16'h18DF7,4);
TASK_PP(16'h18DF8,4);
TASK_PP(16'h18DF9,4);
TASK_PP(16'h18DFA,4);
TASK_PP(16'h18DFB,4);
TASK_PP(16'h18DFC,4);
TASK_PP(16'h18DFD,4);
TASK_PP(16'h18DFE,4);
TASK_PP(16'h18DFF,4);
TASK_PP(16'h18E00,4);
TASK_PP(16'h18E01,4);
TASK_PP(16'h18E02,4);
TASK_PP(16'h18E03,4);
TASK_PP(16'h18E04,4);
TASK_PP(16'h18E05,4);
TASK_PP(16'h18E06,4);
TASK_PP(16'h18E07,4);
TASK_PP(16'h18E08,4);
TASK_PP(16'h18E09,4);
TASK_PP(16'h18E0A,4);
TASK_PP(16'h18E0B,4);
TASK_PP(16'h18E0C,4);
TASK_PP(16'h18E0D,4);
TASK_PP(16'h18E0E,4);
TASK_PP(16'h18E0F,4);
TASK_PP(16'h18E10,4);
TASK_PP(16'h18E11,4);
TASK_PP(16'h18E12,4);
TASK_PP(16'h18E13,4);
TASK_PP(16'h18E14,4);
TASK_PP(16'h18E15,4);
TASK_PP(16'h18E16,4);
TASK_PP(16'h18E17,4);
TASK_PP(16'h18E18,4);
TASK_PP(16'h18E19,4);
TASK_PP(16'h18E1A,4);
TASK_PP(16'h18E1B,4);
TASK_PP(16'h18E1C,4);
TASK_PP(16'h18E1D,4);
TASK_PP(16'h18E1E,4);
TASK_PP(16'h18E1F,4);
TASK_PP(16'h18E20,4);
TASK_PP(16'h18E21,4);
TASK_PP(16'h18E22,4);
TASK_PP(16'h18E23,4);
TASK_PP(16'h18E24,4);
TASK_PP(16'h18E25,4);
TASK_PP(16'h18E26,4);
TASK_PP(16'h18E27,4);
TASK_PP(16'h18E28,4);
TASK_PP(16'h18E29,4);
TASK_PP(16'h18E2A,4);
TASK_PP(16'h18E2B,4);
TASK_PP(16'h18E2C,4);
TASK_PP(16'h18E2D,4);
TASK_PP(16'h18E2E,4);
TASK_PP(16'h18E2F,4);
TASK_PP(16'h18E30,4);
TASK_PP(16'h18E31,4);
TASK_PP(16'h18E32,4);
TASK_PP(16'h18E33,4);
TASK_PP(16'h18E34,4);
TASK_PP(16'h18E35,4);
TASK_PP(16'h18E36,4);
TASK_PP(16'h18E37,4);
TASK_PP(16'h18E38,4);
TASK_PP(16'h18E39,4);
TASK_PP(16'h18E3A,4);
TASK_PP(16'h18E3B,4);
TASK_PP(16'h18E3C,4);
TASK_PP(16'h18E3D,4);
TASK_PP(16'h18E3E,4);
TASK_PP(16'h18E3F,4);
TASK_PP(16'h18E40,4);
TASK_PP(16'h18E41,4);
TASK_PP(16'h18E42,4);
TASK_PP(16'h18E43,4);
TASK_PP(16'h18E44,4);
TASK_PP(16'h18E45,4);
TASK_PP(16'h18E46,4);
TASK_PP(16'h18E47,4);
TASK_PP(16'h18E48,4);
TASK_PP(16'h18E49,4);
TASK_PP(16'h18E4A,4);
TASK_PP(16'h18E4B,4);
TASK_PP(16'h18E4C,4);
TASK_PP(16'h18E4D,4);
TASK_PP(16'h18E4E,4);
TASK_PP(16'h18E4F,4);
TASK_PP(16'h18E50,4);
TASK_PP(16'h18E51,4);
TASK_PP(16'h18E52,4);
TASK_PP(16'h18E53,4);
TASK_PP(16'h18E54,4);
TASK_PP(16'h18E55,4);
TASK_PP(16'h18E56,4);
TASK_PP(16'h18E57,4);
TASK_PP(16'h18E58,4);
TASK_PP(16'h18E59,4);
TASK_PP(16'h18E5A,4);
TASK_PP(16'h18E5B,4);
TASK_PP(16'h18E5C,4);
TASK_PP(16'h18E5D,4);
TASK_PP(16'h18E5E,4);
TASK_PP(16'h18E5F,4);
TASK_PP(16'h18E60,4);
TASK_PP(16'h18E61,4);
TASK_PP(16'h18E62,4);
TASK_PP(16'h18E63,4);
TASK_PP(16'h18E64,4);
TASK_PP(16'h18E65,4);
TASK_PP(16'h18E66,4);
TASK_PP(16'h18E67,4);
TASK_PP(16'h18E68,4);
TASK_PP(16'h18E69,4);
TASK_PP(16'h18E6A,4);
TASK_PP(16'h18E6B,4);
TASK_PP(16'h18E6C,4);
TASK_PP(16'h18E6D,4);
TASK_PP(16'h18E6E,4);
TASK_PP(16'h18E6F,4);
TASK_PP(16'h18E70,4);
TASK_PP(16'h18E71,4);
TASK_PP(16'h18E72,4);
TASK_PP(16'h18E73,4);
TASK_PP(16'h18E74,4);
TASK_PP(16'h18E75,4);
TASK_PP(16'h18E76,4);
TASK_PP(16'h18E77,4);
TASK_PP(16'h18E78,4);
TASK_PP(16'h18E79,4);
TASK_PP(16'h18E7A,4);
TASK_PP(16'h18E7B,4);
TASK_PP(16'h18E7C,4);
TASK_PP(16'h18E7D,4);
TASK_PP(16'h18E7E,4);
TASK_PP(16'h18E7F,4);
TASK_PP(16'h18E80,4);
TASK_PP(16'h18E81,4);
TASK_PP(16'h18E82,4);
TASK_PP(16'h18E83,4);
TASK_PP(16'h18E84,4);
TASK_PP(16'h18E85,4);
TASK_PP(16'h18E86,4);
TASK_PP(16'h18E87,4);
TASK_PP(16'h18E88,4);
TASK_PP(16'h18E89,4);
TASK_PP(16'h18E8A,4);
TASK_PP(16'h18E8B,4);
TASK_PP(16'h18E8C,4);
TASK_PP(16'h18E8D,4);
TASK_PP(16'h18E8E,4);
TASK_PP(16'h18E8F,4);
TASK_PP(16'h18E90,4);
TASK_PP(16'h18E91,4);
TASK_PP(16'h18E92,4);
TASK_PP(16'h18E93,4);
TASK_PP(16'h18E94,4);
TASK_PP(16'h18E95,4);
TASK_PP(16'h18E96,4);
TASK_PP(16'h18E97,4);
TASK_PP(16'h18E98,4);
TASK_PP(16'h18E99,4);
TASK_PP(16'h18E9A,4);
TASK_PP(16'h18E9B,4);
TASK_PP(16'h18E9C,4);
TASK_PP(16'h18E9D,4);
TASK_PP(16'h18E9E,4);
TASK_PP(16'h18E9F,4);
TASK_PP(16'h18EA0,4);
TASK_PP(16'h18EA1,4);
TASK_PP(16'h18EA2,4);
TASK_PP(16'h18EA3,4);
TASK_PP(16'h18EA4,4);
TASK_PP(16'h18EA5,4);
TASK_PP(16'h18EA6,4);
TASK_PP(16'h18EA7,4);
TASK_PP(16'h18EA8,4);
TASK_PP(16'h18EA9,4);
TASK_PP(16'h18EAA,4);
TASK_PP(16'h18EAB,4);
TASK_PP(16'h18EAC,4);
TASK_PP(16'h18EAD,4);
TASK_PP(16'h18EAE,4);
TASK_PP(16'h18EAF,4);
TASK_PP(16'h18EB0,4);
TASK_PP(16'h18EB1,4);
TASK_PP(16'h18EB2,4);
TASK_PP(16'h18EB3,4);
TASK_PP(16'h18EB4,4);
TASK_PP(16'h18EB5,4);
TASK_PP(16'h18EB6,4);
TASK_PP(16'h18EB7,4);
TASK_PP(16'h18EB8,4);
TASK_PP(16'h18EB9,4);
TASK_PP(16'h18EBA,4);
TASK_PP(16'h18EBB,4);
TASK_PP(16'h18EBC,4);
TASK_PP(16'h18EBD,4);
TASK_PP(16'h18EBE,4);
TASK_PP(16'h18EBF,4);
TASK_PP(16'h18EC0,4);
TASK_PP(16'h18EC1,4);
TASK_PP(16'h18EC2,4);
TASK_PP(16'h18EC3,4);
TASK_PP(16'h18EC4,4);
TASK_PP(16'h18EC5,4);
TASK_PP(16'h18EC6,4);
TASK_PP(16'h18EC7,4);
TASK_PP(16'h18EC8,4);
TASK_PP(16'h18EC9,4);
TASK_PP(16'h18ECA,4);
TASK_PP(16'h18ECB,4);
TASK_PP(16'h18ECC,4);
TASK_PP(16'h18ECD,4);
TASK_PP(16'h18ECE,4);
TASK_PP(16'h18ECF,4);
TASK_PP(16'h18ED0,4);
TASK_PP(16'h18ED1,4);
TASK_PP(16'h18ED2,4);
TASK_PP(16'h18ED3,4);
TASK_PP(16'h18ED4,4);
TASK_PP(16'h18ED5,4);
TASK_PP(16'h18ED6,4);
TASK_PP(16'h18ED7,4);
TASK_PP(16'h18ED8,4);
TASK_PP(16'h18ED9,4);
TASK_PP(16'h18EDA,4);
TASK_PP(16'h18EDB,4);
TASK_PP(16'h18EDC,4);
TASK_PP(16'h18EDD,4);
TASK_PP(16'h18EDE,4);
TASK_PP(16'h18EDF,4);
TASK_PP(16'h18EE0,4);
TASK_PP(16'h18EE1,4);
TASK_PP(16'h18EE2,4);
TASK_PP(16'h18EE3,4);
TASK_PP(16'h18EE4,4);
TASK_PP(16'h18EE5,4);
TASK_PP(16'h18EE6,4);
TASK_PP(16'h18EE7,4);
TASK_PP(16'h18EE8,4);
TASK_PP(16'h18EE9,4);
TASK_PP(16'h18EEA,4);
TASK_PP(16'h18EEB,4);
TASK_PP(16'h18EEC,4);
TASK_PP(16'h18EED,4);
TASK_PP(16'h18EEE,4);
TASK_PP(16'h18EEF,4);
TASK_PP(16'h18EF0,4);
TASK_PP(16'h18EF1,4);
TASK_PP(16'h18EF2,4);
TASK_PP(16'h18EF3,4);
TASK_PP(16'h18EF4,4);
TASK_PP(16'h18EF5,4);
TASK_PP(16'h18EF6,4);
TASK_PP(16'h18EF7,4);
TASK_PP(16'h18EF8,4);
TASK_PP(16'h18EF9,4);
TASK_PP(16'h18EFA,4);
TASK_PP(16'h18EFB,4);
TASK_PP(16'h18EFC,4);
TASK_PP(16'h18EFD,4);
TASK_PP(16'h18EFE,4);
TASK_PP(16'h18EFF,4);
TASK_PP(16'h18F00,4);
TASK_PP(16'h18F01,4);
TASK_PP(16'h18F02,4);
TASK_PP(16'h18F03,4);
TASK_PP(16'h18F04,4);
TASK_PP(16'h18F05,4);
TASK_PP(16'h18F06,4);
TASK_PP(16'h18F07,4);
TASK_PP(16'h18F08,4);
TASK_PP(16'h18F09,4);
TASK_PP(16'h18F0A,4);
TASK_PP(16'h18F0B,4);
TASK_PP(16'h18F0C,4);
TASK_PP(16'h18F0D,4);
TASK_PP(16'h18F0E,4);
TASK_PP(16'h18F0F,4);
TASK_PP(16'h18F10,4);
TASK_PP(16'h18F11,4);
TASK_PP(16'h18F12,4);
TASK_PP(16'h18F13,4);
TASK_PP(16'h18F14,4);
TASK_PP(16'h18F15,4);
TASK_PP(16'h18F16,4);
TASK_PP(16'h18F17,4);
TASK_PP(16'h18F18,4);
TASK_PP(16'h18F19,4);
TASK_PP(16'h18F1A,4);
TASK_PP(16'h18F1B,4);
TASK_PP(16'h18F1C,4);
TASK_PP(16'h18F1D,4);
TASK_PP(16'h18F1E,4);
TASK_PP(16'h18F1F,4);
TASK_PP(16'h18F20,4);
TASK_PP(16'h18F21,4);
TASK_PP(16'h18F22,4);
TASK_PP(16'h18F23,4);
TASK_PP(16'h18F24,4);
TASK_PP(16'h18F25,4);
TASK_PP(16'h18F26,4);
TASK_PP(16'h18F27,4);
TASK_PP(16'h18F28,4);
TASK_PP(16'h18F29,4);
TASK_PP(16'h18F2A,4);
TASK_PP(16'h18F2B,4);
TASK_PP(16'h18F2C,4);
TASK_PP(16'h18F2D,4);
TASK_PP(16'h18F2E,4);
TASK_PP(16'h18F2F,4);
TASK_PP(16'h18F30,4);
TASK_PP(16'h18F31,4);
TASK_PP(16'h18F32,4);
TASK_PP(16'h18F33,4);
TASK_PP(16'h18F34,4);
TASK_PP(16'h18F35,4);
TASK_PP(16'h18F36,4);
TASK_PP(16'h18F37,4);
TASK_PP(16'h18F38,4);
TASK_PP(16'h18F39,4);
TASK_PP(16'h18F3A,4);
TASK_PP(16'h18F3B,4);
TASK_PP(16'h18F3C,4);
TASK_PP(16'h18F3D,4);
TASK_PP(16'h18F3E,4);
TASK_PP(16'h18F3F,4);
TASK_PP(16'h18F40,4);
TASK_PP(16'h18F41,4);
TASK_PP(16'h18F42,4);
TASK_PP(16'h18F43,4);
TASK_PP(16'h18F44,4);
TASK_PP(16'h18F45,4);
TASK_PP(16'h18F46,4);
TASK_PP(16'h18F47,4);
TASK_PP(16'h18F48,4);
TASK_PP(16'h18F49,4);
TASK_PP(16'h18F4A,4);
TASK_PP(16'h18F4B,4);
TASK_PP(16'h18F4C,4);
TASK_PP(16'h18F4D,4);
TASK_PP(16'h18F4E,4);
TASK_PP(16'h18F4F,4);
TASK_PP(16'h18F50,4);
TASK_PP(16'h18F51,4);
TASK_PP(16'h18F52,4);
TASK_PP(16'h18F53,4);
TASK_PP(16'h18F54,4);
TASK_PP(16'h18F55,4);
TASK_PP(16'h18F56,4);
TASK_PP(16'h18F57,4);
TASK_PP(16'h18F58,4);
TASK_PP(16'h18F59,4);
TASK_PP(16'h18F5A,4);
TASK_PP(16'h18F5B,4);
TASK_PP(16'h18F5C,4);
TASK_PP(16'h18F5D,4);
TASK_PP(16'h18F5E,4);
TASK_PP(16'h18F5F,4);
TASK_PP(16'h18F60,4);
TASK_PP(16'h18F61,4);
TASK_PP(16'h18F62,4);
TASK_PP(16'h18F63,4);
TASK_PP(16'h18F64,4);
TASK_PP(16'h18F65,4);
TASK_PP(16'h18F66,4);
TASK_PP(16'h18F67,4);
TASK_PP(16'h18F68,4);
TASK_PP(16'h18F69,4);
TASK_PP(16'h18F6A,4);
TASK_PP(16'h18F6B,4);
TASK_PP(16'h18F6C,4);
TASK_PP(16'h18F6D,4);
TASK_PP(16'h18F6E,4);
TASK_PP(16'h18F6F,4);
TASK_PP(16'h18F70,4);
TASK_PP(16'h18F71,4);
TASK_PP(16'h18F72,4);
TASK_PP(16'h18F73,4);
TASK_PP(16'h18F74,4);
TASK_PP(16'h18F75,4);
TASK_PP(16'h18F76,4);
TASK_PP(16'h18F77,4);
TASK_PP(16'h18F78,4);
TASK_PP(16'h18F79,4);
TASK_PP(16'h18F7A,4);
TASK_PP(16'h18F7B,4);
TASK_PP(16'h18F7C,4);
TASK_PP(16'h18F7D,4);
TASK_PP(16'h18F7E,4);
TASK_PP(16'h18F7F,4);
TASK_PP(16'h18F80,4);
TASK_PP(16'h18F81,4);
TASK_PP(16'h18F82,4);
TASK_PP(16'h18F83,4);
TASK_PP(16'h18F84,4);
TASK_PP(16'h18F85,4);
TASK_PP(16'h18F86,4);
TASK_PP(16'h18F87,4);
TASK_PP(16'h18F88,4);
TASK_PP(16'h18F89,4);
TASK_PP(16'h18F8A,4);
TASK_PP(16'h18F8B,4);
TASK_PP(16'h18F8C,4);
TASK_PP(16'h18F8D,4);
TASK_PP(16'h18F8E,4);
TASK_PP(16'h18F8F,4);
TASK_PP(16'h18F90,4);
TASK_PP(16'h18F91,4);
TASK_PP(16'h18F92,4);
TASK_PP(16'h18F93,4);
TASK_PP(16'h18F94,4);
TASK_PP(16'h18F95,4);
TASK_PP(16'h18F96,4);
TASK_PP(16'h18F97,4);
TASK_PP(16'h18F98,4);
TASK_PP(16'h18F99,4);
TASK_PP(16'h18F9A,4);
TASK_PP(16'h18F9B,4);
TASK_PP(16'h18F9C,4);
TASK_PP(16'h18F9D,4);
TASK_PP(16'h18F9E,4);
TASK_PP(16'h18F9F,4);
TASK_PP(16'h18FA0,4);
TASK_PP(16'h18FA1,4);
TASK_PP(16'h18FA2,4);
TASK_PP(16'h18FA3,4);
TASK_PP(16'h18FA4,4);
TASK_PP(16'h18FA5,4);
TASK_PP(16'h18FA6,4);
TASK_PP(16'h18FA7,4);
TASK_PP(16'h18FA8,4);
TASK_PP(16'h18FA9,4);
TASK_PP(16'h18FAA,4);
TASK_PP(16'h18FAB,4);
TASK_PP(16'h18FAC,4);
TASK_PP(16'h18FAD,4);
TASK_PP(16'h18FAE,4);
TASK_PP(16'h18FAF,4);
TASK_PP(16'h18FB0,4);
TASK_PP(16'h18FB1,4);
TASK_PP(16'h18FB2,4);
TASK_PP(16'h18FB3,4);
TASK_PP(16'h18FB4,4);
TASK_PP(16'h18FB5,4);
TASK_PP(16'h18FB6,4);
TASK_PP(16'h18FB7,4);
TASK_PP(16'h18FB8,4);
TASK_PP(16'h18FB9,4);
TASK_PP(16'h18FBA,4);
TASK_PP(16'h18FBB,4);
TASK_PP(16'h18FBC,4);
TASK_PP(16'h18FBD,4);
TASK_PP(16'h18FBE,4);
TASK_PP(16'h18FBF,4);
TASK_PP(16'h18FC0,4);
TASK_PP(16'h18FC1,4);
TASK_PP(16'h18FC2,4);
TASK_PP(16'h18FC3,4);
TASK_PP(16'h18FC4,4);
TASK_PP(16'h18FC5,4);
TASK_PP(16'h18FC6,4);
TASK_PP(16'h18FC7,4);
TASK_PP(16'h18FC8,4);
TASK_PP(16'h18FC9,4);
TASK_PP(16'h18FCA,4);
TASK_PP(16'h18FCB,4);
TASK_PP(16'h18FCC,4);
TASK_PP(16'h18FCD,4);
TASK_PP(16'h18FCE,4);
TASK_PP(16'h18FCF,4);
TASK_PP(16'h18FD0,4);
TASK_PP(16'h18FD1,4);
TASK_PP(16'h18FD2,4);
TASK_PP(16'h18FD3,4);
TASK_PP(16'h18FD4,4);
TASK_PP(16'h18FD5,4);
TASK_PP(16'h18FD6,4);
TASK_PP(16'h18FD7,4);
TASK_PP(16'h18FD8,4);
TASK_PP(16'h18FD9,4);
TASK_PP(16'h18FDA,4);
TASK_PP(16'h18FDB,4);
TASK_PP(16'h18FDC,4);
TASK_PP(16'h18FDD,4);
TASK_PP(16'h18FDE,4);
TASK_PP(16'h18FDF,4);
TASK_PP(16'h18FE0,4);
TASK_PP(16'h18FE1,4);
TASK_PP(16'h18FE2,4);
TASK_PP(16'h18FE3,4);
TASK_PP(16'h18FE4,4);
TASK_PP(16'h18FE5,4);
TASK_PP(16'h18FE6,4);
TASK_PP(16'h18FE7,4);
TASK_PP(16'h18FE8,4);
TASK_PP(16'h18FE9,4);
TASK_PP(16'h18FEA,4);
TASK_PP(16'h18FEB,4);
TASK_PP(16'h18FEC,4);
TASK_PP(16'h18FED,4);
TASK_PP(16'h18FEE,4);
TASK_PP(16'h18FEF,4);
TASK_PP(16'h18FF0,4);
TASK_PP(16'h18FF1,4);
TASK_PP(16'h18FF2,4);
TASK_PP(16'h18FF3,4);
TASK_PP(16'h18FF4,4);
TASK_PP(16'h18FF5,4);
TASK_PP(16'h18FF6,4);
TASK_PP(16'h18FF7,4);
TASK_PP(16'h18FF8,4);
TASK_PP(16'h18FF9,4);
TASK_PP(16'h18FFA,4);
TASK_PP(16'h18FFB,4);
TASK_PP(16'h18FFC,4);
TASK_PP(16'h18FFD,4);
TASK_PP(16'h18FFE,4);
TASK_PP(16'h18FFF,4);
TASK_PP(16'h19000,4);
TASK_PP(16'h19001,4);
TASK_PP(16'h19002,4);
TASK_PP(16'h19003,4);
TASK_PP(16'h19004,4);
TASK_PP(16'h19005,4);
TASK_PP(16'h19006,4);
TASK_PP(16'h19007,4);
TASK_PP(16'h19008,4);
TASK_PP(16'h19009,4);
TASK_PP(16'h1900A,4);
TASK_PP(16'h1900B,4);
TASK_PP(16'h1900C,4);
TASK_PP(16'h1900D,4);
TASK_PP(16'h1900E,4);
TASK_PP(16'h1900F,4);
TASK_PP(16'h19010,4);
TASK_PP(16'h19011,4);
TASK_PP(16'h19012,4);
TASK_PP(16'h19013,4);
TASK_PP(16'h19014,4);
TASK_PP(16'h19015,4);
TASK_PP(16'h19016,4);
TASK_PP(16'h19017,4);
TASK_PP(16'h19018,4);
TASK_PP(16'h19019,4);
TASK_PP(16'h1901A,4);
TASK_PP(16'h1901B,4);
TASK_PP(16'h1901C,4);
TASK_PP(16'h1901D,4);
TASK_PP(16'h1901E,4);
TASK_PP(16'h1901F,4);
TASK_PP(16'h19020,4);
TASK_PP(16'h19021,4);
TASK_PP(16'h19022,4);
TASK_PP(16'h19023,4);
TASK_PP(16'h19024,4);
TASK_PP(16'h19025,4);
TASK_PP(16'h19026,4);
TASK_PP(16'h19027,4);
TASK_PP(16'h19028,4);
TASK_PP(16'h19029,4);
TASK_PP(16'h1902A,4);
TASK_PP(16'h1902B,4);
TASK_PP(16'h1902C,4);
TASK_PP(16'h1902D,4);
TASK_PP(16'h1902E,4);
TASK_PP(16'h1902F,4);
TASK_PP(16'h19030,4);
TASK_PP(16'h19031,4);
TASK_PP(16'h19032,4);
TASK_PP(16'h19033,4);
TASK_PP(16'h19034,4);
TASK_PP(16'h19035,4);
TASK_PP(16'h19036,4);
TASK_PP(16'h19037,4);
TASK_PP(16'h19038,4);
TASK_PP(16'h19039,4);
TASK_PP(16'h1903A,4);
TASK_PP(16'h1903B,4);
TASK_PP(16'h1903C,4);
TASK_PP(16'h1903D,4);
TASK_PP(16'h1903E,4);
TASK_PP(16'h1903F,4);
TASK_PP(16'h19040,4);
TASK_PP(16'h19041,4);
TASK_PP(16'h19042,4);
TASK_PP(16'h19043,4);
TASK_PP(16'h19044,4);
TASK_PP(16'h19045,4);
TASK_PP(16'h19046,4);
TASK_PP(16'h19047,4);
TASK_PP(16'h19048,4);
TASK_PP(16'h19049,4);
TASK_PP(16'h1904A,4);
TASK_PP(16'h1904B,4);
TASK_PP(16'h1904C,4);
TASK_PP(16'h1904D,4);
TASK_PP(16'h1904E,4);
TASK_PP(16'h1904F,4);
TASK_PP(16'h19050,4);
TASK_PP(16'h19051,4);
TASK_PP(16'h19052,4);
TASK_PP(16'h19053,4);
TASK_PP(16'h19054,4);
TASK_PP(16'h19055,4);
TASK_PP(16'h19056,4);
TASK_PP(16'h19057,4);
TASK_PP(16'h19058,4);
TASK_PP(16'h19059,4);
TASK_PP(16'h1905A,4);
TASK_PP(16'h1905B,4);
TASK_PP(16'h1905C,4);
TASK_PP(16'h1905D,4);
TASK_PP(16'h1905E,4);
TASK_PP(16'h1905F,4);
TASK_PP(16'h19060,4);
TASK_PP(16'h19061,4);
TASK_PP(16'h19062,4);
TASK_PP(16'h19063,4);
TASK_PP(16'h19064,4);
TASK_PP(16'h19065,4);
TASK_PP(16'h19066,4);
TASK_PP(16'h19067,4);
TASK_PP(16'h19068,4);
TASK_PP(16'h19069,4);
TASK_PP(16'h1906A,4);
TASK_PP(16'h1906B,4);
TASK_PP(16'h1906C,4);
TASK_PP(16'h1906D,4);
TASK_PP(16'h1906E,4);
TASK_PP(16'h1906F,4);
TASK_PP(16'h19070,4);
TASK_PP(16'h19071,4);
TASK_PP(16'h19072,4);
TASK_PP(16'h19073,4);
TASK_PP(16'h19074,4);
TASK_PP(16'h19075,4);
TASK_PP(16'h19076,4);
TASK_PP(16'h19077,4);
TASK_PP(16'h19078,4);
TASK_PP(16'h19079,4);
TASK_PP(16'h1907A,4);
TASK_PP(16'h1907B,4);
TASK_PP(16'h1907C,4);
TASK_PP(16'h1907D,4);
TASK_PP(16'h1907E,4);
TASK_PP(16'h1907F,4);
TASK_PP(16'h19080,4);
TASK_PP(16'h19081,4);
TASK_PP(16'h19082,4);
TASK_PP(16'h19083,4);
TASK_PP(16'h19084,4);
TASK_PP(16'h19085,4);
TASK_PP(16'h19086,4);
TASK_PP(16'h19087,4);
TASK_PP(16'h19088,4);
TASK_PP(16'h19089,4);
TASK_PP(16'h1908A,4);
TASK_PP(16'h1908B,4);
TASK_PP(16'h1908C,4);
TASK_PP(16'h1908D,4);
TASK_PP(16'h1908E,4);
TASK_PP(16'h1908F,4);
TASK_PP(16'h19090,4);
TASK_PP(16'h19091,4);
TASK_PP(16'h19092,4);
TASK_PP(16'h19093,4);
TASK_PP(16'h19094,4);
TASK_PP(16'h19095,4);
TASK_PP(16'h19096,4);
TASK_PP(16'h19097,4);
TASK_PP(16'h19098,4);
TASK_PP(16'h19099,4);
TASK_PP(16'h1909A,4);
TASK_PP(16'h1909B,4);
TASK_PP(16'h1909C,4);
TASK_PP(16'h1909D,4);
TASK_PP(16'h1909E,4);
TASK_PP(16'h1909F,4);
TASK_PP(16'h190A0,4);
TASK_PP(16'h190A1,4);
TASK_PP(16'h190A2,4);
TASK_PP(16'h190A3,4);
TASK_PP(16'h190A4,4);
TASK_PP(16'h190A5,4);
TASK_PP(16'h190A6,4);
TASK_PP(16'h190A7,4);
TASK_PP(16'h190A8,4);
TASK_PP(16'h190A9,4);
TASK_PP(16'h190AA,4);
TASK_PP(16'h190AB,4);
TASK_PP(16'h190AC,4);
TASK_PP(16'h190AD,4);
TASK_PP(16'h190AE,4);
TASK_PP(16'h190AF,4);
TASK_PP(16'h190B0,4);
TASK_PP(16'h190B1,4);
TASK_PP(16'h190B2,4);
TASK_PP(16'h190B3,4);
TASK_PP(16'h190B4,4);
TASK_PP(16'h190B5,4);
TASK_PP(16'h190B6,4);
TASK_PP(16'h190B7,4);
TASK_PP(16'h190B8,4);
TASK_PP(16'h190B9,4);
TASK_PP(16'h190BA,4);
TASK_PP(16'h190BB,4);
TASK_PP(16'h190BC,4);
TASK_PP(16'h190BD,4);
TASK_PP(16'h190BE,4);
TASK_PP(16'h190BF,4);
TASK_PP(16'h190C0,4);
TASK_PP(16'h190C1,4);
TASK_PP(16'h190C2,4);
TASK_PP(16'h190C3,4);
TASK_PP(16'h190C4,4);
TASK_PP(16'h190C5,4);
TASK_PP(16'h190C6,4);
TASK_PP(16'h190C7,4);
TASK_PP(16'h190C8,4);
TASK_PP(16'h190C9,4);
TASK_PP(16'h190CA,4);
TASK_PP(16'h190CB,4);
TASK_PP(16'h190CC,4);
TASK_PP(16'h190CD,4);
TASK_PP(16'h190CE,4);
TASK_PP(16'h190CF,4);
TASK_PP(16'h190D0,4);
TASK_PP(16'h190D1,4);
TASK_PP(16'h190D2,4);
TASK_PP(16'h190D3,4);
TASK_PP(16'h190D4,4);
TASK_PP(16'h190D5,4);
TASK_PP(16'h190D6,4);
TASK_PP(16'h190D7,4);
TASK_PP(16'h190D8,4);
TASK_PP(16'h190D9,4);
TASK_PP(16'h190DA,4);
TASK_PP(16'h190DB,4);
TASK_PP(16'h190DC,4);
TASK_PP(16'h190DD,4);
TASK_PP(16'h190DE,4);
TASK_PP(16'h190DF,4);
TASK_PP(16'h190E0,4);
TASK_PP(16'h190E1,4);
TASK_PP(16'h190E2,4);
TASK_PP(16'h190E3,4);
TASK_PP(16'h190E4,4);
TASK_PP(16'h190E5,4);
TASK_PP(16'h190E6,4);
TASK_PP(16'h190E7,4);
TASK_PP(16'h190E8,4);
TASK_PP(16'h190E9,4);
TASK_PP(16'h190EA,4);
TASK_PP(16'h190EB,4);
TASK_PP(16'h190EC,4);
TASK_PP(16'h190ED,4);
TASK_PP(16'h190EE,4);
TASK_PP(16'h190EF,4);
TASK_PP(16'h190F0,4);
TASK_PP(16'h190F1,4);
TASK_PP(16'h190F2,4);
TASK_PP(16'h190F3,4);
TASK_PP(16'h190F4,4);
TASK_PP(16'h190F5,4);
TASK_PP(16'h190F6,4);
TASK_PP(16'h190F7,4);
TASK_PP(16'h190F8,4);
TASK_PP(16'h190F9,4);
TASK_PP(16'h190FA,4);
TASK_PP(16'h190FB,4);
TASK_PP(16'h190FC,4);
TASK_PP(16'h190FD,4);
TASK_PP(16'h190FE,4);
TASK_PP(16'h190FF,4);
TASK_PP(16'h19100,4);
TASK_PP(16'h19101,4);
TASK_PP(16'h19102,4);
TASK_PP(16'h19103,4);
TASK_PP(16'h19104,4);
TASK_PP(16'h19105,4);
TASK_PP(16'h19106,4);
TASK_PP(16'h19107,4);
TASK_PP(16'h19108,4);
TASK_PP(16'h19109,4);
TASK_PP(16'h1910A,4);
TASK_PP(16'h1910B,4);
TASK_PP(16'h1910C,4);
TASK_PP(16'h1910D,4);
TASK_PP(16'h1910E,4);
TASK_PP(16'h1910F,4);
TASK_PP(16'h19110,4);
TASK_PP(16'h19111,4);
TASK_PP(16'h19112,4);
TASK_PP(16'h19113,4);
TASK_PP(16'h19114,4);
TASK_PP(16'h19115,4);
TASK_PP(16'h19116,4);
TASK_PP(16'h19117,4);
TASK_PP(16'h19118,4);
TASK_PP(16'h19119,4);
TASK_PP(16'h1911A,4);
TASK_PP(16'h1911B,4);
TASK_PP(16'h1911C,4);
TASK_PP(16'h1911D,4);
TASK_PP(16'h1911E,4);
TASK_PP(16'h1911F,4);
TASK_PP(16'h19120,4);
TASK_PP(16'h19121,4);
TASK_PP(16'h19122,4);
TASK_PP(16'h19123,4);
TASK_PP(16'h19124,4);
TASK_PP(16'h19125,4);
TASK_PP(16'h19126,4);
TASK_PP(16'h19127,4);
TASK_PP(16'h19128,4);
TASK_PP(16'h19129,4);
TASK_PP(16'h1912A,4);
TASK_PP(16'h1912B,4);
TASK_PP(16'h1912C,4);
TASK_PP(16'h1912D,4);
TASK_PP(16'h1912E,4);
TASK_PP(16'h1912F,4);
TASK_PP(16'h19130,4);
TASK_PP(16'h19131,4);
TASK_PP(16'h19132,4);
TASK_PP(16'h19133,4);
TASK_PP(16'h19134,4);
TASK_PP(16'h19135,4);
TASK_PP(16'h19136,4);
TASK_PP(16'h19137,4);
TASK_PP(16'h19138,4);
TASK_PP(16'h19139,4);
TASK_PP(16'h1913A,4);
TASK_PP(16'h1913B,4);
TASK_PP(16'h1913C,4);
TASK_PP(16'h1913D,4);
TASK_PP(16'h1913E,4);
TASK_PP(16'h1913F,4);
TASK_PP(16'h19140,4);
TASK_PP(16'h19141,4);
TASK_PP(16'h19142,4);
TASK_PP(16'h19143,4);
TASK_PP(16'h19144,4);
TASK_PP(16'h19145,4);
TASK_PP(16'h19146,4);
TASK_PP(16'h19147,4);
TASK_PP(16'h19148,4);
TASK_PP(16'h19149,4);
TASK_PP(16'h1914A,4);
TASK_PP(16'h1914B,4);
TASK_PP(16'h1914C,4);
TASK_PP(16'h1914D,4);
TASK_PP(16'h1914E,4);
TASK_PP(16'h1914F,4);
TASK_PP(16'h19150,4);
TASK_PP(16'h19151,4);
TASK_PP(16'h19152,4);
TASK_PP(16'h19153,4);
TASK_PP(16'h19154,4);
TASK_PP(16'h19155,4);
TASK_PP(16'h19156,4);
TASK_PP(16'h19157,4);
TASK_PP(16'h19158,4);
TASK_PP(16'h19159,4);
TASK_PP(16'h1915A,4);
TASK_PP(16'h1915B,4);
TASK_PP(16'h1915C,4);
TASK_PP(16'h1915D,4);
TASK_PP(16'h1915E,4);
TASK_PP(16'h1915F,4);
TASK_PP(16'h19160,4);
TASK_PP(16'h19161,4);
TASK_PP(16'h19162,4);
TASK_PP(16'h19163,4);
TASK_PP(16'h19164,4);
TASK_PP(16'h19165,4);
TASK_PP(16'h19166,4);
TASK_PP(16'h19167,4);
TASK_PP(16'h19168,4);
TASK_PP(16'h19169,4);
TASK_PP(16'h1916A,4);
TASK_PP(16'h1916B,4);
TASK_PP(16'h1916C,4);
TASK_PP(16'h1916D,4);
TASK_PP(16'h1916E,4);
TASK_PP(16'h1916F,4);
TASK_PP(16'h19170,4);
TASK_PP(16'h19171,4);
TASK_PP(16'h19172,4);
TASK_PP(16'h19173,4);
TASK_PP(16'h19174,4);
TASK_PP(16'h19175,4);
TASK_PP(16'h19176,4);
TASK_PP(16'h19177,4);
TASK_PP(16'h19178,4);
TASK_PP(16'h19179,4);
TASK_PP(16'h1917A,4);
TASK_PP(16'h1917B,4);
TASK_PP(16'h1917C,4);
TASK_PP(16'h1917D,4);
TASK_PP(16'h1917E,4);
TASK_PP(16'h1917F,4);
TASK_PP(16'h19180,4);
TASK_PP(16'h19181,4);
TASK_PP(16'h19182,4);
TASK_PP(16'h19183,4);
TASK_PP(16'h19184,4);
TASK_PP(16'h19185,4);
TASK_PP(16'h19186,4);
TASK_PP(16'h19187,4);
TASK_PP(16'h19188,4);
TASK_PP(16'h19189,4);
TASK_PP(16'h1918A,4);
TASK_PP(16'h1918B,4);
TASK_PP(16'h1918C,4);
TASK_PP(16'h1918D,4);
TASK_PP(16'h1918E,4);
TASK_PP(16'h1918F,4);
TASK_PP(16'h19190,4);
TASK_PP(16'h19191,4);
TASK_PP(16'h19192,4);
TASK_PP(16'h19193,4);
TASK_PP(16'h19194,4);
TASK_PP(16'h19195,4);
TASK_PP(16'h19196,4);
TASK_PP(16'h19197,4);
TASK_PP(16'h19198,4);
TASK_PP(16'h19199,4);
TASK_PP(16'h1919A,4);
TASK_PP(16'h1919B,4);
TASK_PP(16'h1919C,4);
TASK_PP(16'h1919D,4);
TASK_PP(16'h1919E,4);
TASK_PP(16'h1919F,4);
TASK_PP(16'h191A0,4);
TASK_PP(16'h191A1,4);
TASK_PP(16'h191A2,4);
TASK_PP(16'h191A3,4);
TASK_PP(16'h191A4,4);
TASK_PP(16'h191A5,4);
TASK_PP(16'h191A6,4);
TASK_PP(16'h191A7,4);
TASK_PP(16'h191A8,4);
TASK_PP(16'h191A9,4);
TASK_PP(16'h191AA,4);
TASK_PP(16'h191AB,4);
TASK_PP(16'h191AC,4);
TASK_PP(16'h191AD,4);
TASK_PP(16'h191AE,4);
TASK_PP(16'h191AF,4);
TASK_PP(16'h191B0,4);
TASK_PP(16'h191B1,4);
TASK_PP(16'h191B2,4);
TASK_PP(16'h191B3,4);
TASK_PP(16'h191B4,4);
TASK_PP(16'h191B5,4);
TASK_PP(16'h191B6,4);
TASK_PP(16'h191B7,4);
TASK_PP(16'h191B8,4);
TASK_PP(16'h191B9,4);
TASK_PP(16'h191BA,4);
TASK_PP(16'h191BB,4);
TASK_PP(16'h191BC,4);
TASK_PP(16'h191BD,4);
TASK_PP(16'h191BE,4);
TASK_PP(16'h191BF,4);
TASK_PP(16'h191C0,4);
TASK_PP(16'h191C1,4);
TASK_PP(16'h191C2,4);
TASK_PP(16'h191C3,4);
TASK_PP(16'h191C4,4);
TASK_PP(16'h191C5,4);
TASK_PP(16'h191C6,4);
TASK_PP(16'h191C7,4);
TASK_PP(16'h191C8,4);
TASK_PP(16'h191C9,4);
TASK_PP(16'h191CA,4);
TASK_PP(16'h191CB,4);
TASK_PP(16'h191CC,4);
TASK_PP(16'h191CD,4);
TASK_PP(16'h191CE,4);
TASK_PP(16'h191CF,4);
TASK_PP(16'h191D0,4);
TASK_PP(16'h191D1,4);
TASK_PP(16'h191D2,4);
TASK_PP(16'h191D3,4);
TASK_PP(16'h191D4,4);
TASK_PP(16'h191D5,4);
TASK_PP(16'h191D6,4);
TASK_PP(16'h191D7,4);
TASK_PP(16'h191D8,4);
TASK_PP(16'h191D9,4);
TASK_PP(16'h191DA,4);
TASK_PP(16'h191DB,4);
TASK_PP(16'h191DC,4);
TASK_PP(16'h191DD,4);
TASK_PP(16'h191DE,4);
TASK_PP(16'h191DF,4);
TASK_PP(16'h191E0,4);
TASK_PP(16'h191E1,4);
TASK_PP(16'h191E2,4);
TASK_PP(16'h191E3,4);
TASK_PP(16'h191E4,4);
TASK_PP(16'h191E5,4);
TASK_PP(16'h191E6,4);
TASK_PP(16'h191E7,4);
TASK_PP(16'h191E8,4);
TASK_PP(16'h191E9,4);
TASK_PP(16'h191EA,4);
TASK_PP(16'h191EB,4);
TASK_PP(16'h191EC,4);
TASK_PP(16'h191ED,4);
TASK_PP(16'h191EE,4);
TASK_PP(16'h191EF,4);
TASK_PP(16'h191F0,4);
TASK_PP(16'h191F1,4);
TASK_PP(16'h191F2,4);
TASK_PP(16'h191F3,4);
TASK_PP(16'h191F4,4);
TASK_PP(16'h191F5,4);
TASK_PP(16'h191F6,4);
TASK_PP(16'h191F7,4);
TASK_PP(16'h191F8,4);
TASK_PP(16'h191F9,4);
TASK_PP(16'h191FA,4);
TASK_PP(16'h191FB,4);
TASK_PP(16'h191FC,4);
TASK_PP(16'h191FD,4);
TASK_PP(16'h191FE,4);
TASK_PP(16'h191FF,4);
TASK_PP(16'h19200,4);
TASK_PP(16'h19201,4);
TASK_PP(16'h19202,4);
TASK_PP(16'h19203,4);
TASK_PP(16'h19204,4);
TASK_PP(16'h19205,4);
TASK_PP(16'h19206,4);
TASK_PP(16'h19207,4);
TASK_PP(16'h19208,4);
TASK_PP(16'h19209,4);
TASK_PP(16'h1920A,4);
TASK_PP(16'h1920B,4);
TASK_PP(16'h1920C,4);
TASK_PP(16'h1920D,4);
TASK_PP(16'h1920E,4);
TASK_PP(16'h1920F,4);
TASK_PP(16'h19210,4);
TASK_PP(16'h19211,4);
TASK_PP(16'h19212,4);
TASK_PP(16'h19213,4);
TASK_PP(16'h19214,4);
TASK_PP(16'h19215,4);
TASK_PP(16'h19216,4);
TASK_PP(16'h19217,4);
TASK_PP(16'h19218,4);
TASK_PP(16'h19219,4);
TASK_PP(16'h1921A,4);
TASK_PP(16'h1921B,4);
TASK_PP(16'h1921C,4);
TASK_PP(16'h1921D,4);
TASK_PP(16'h1921E,4);
TASK_PP(16'h1921F,4);
TASK_PP(16'h19220,4);
TASK_PP(16'h19221,4);
TASK_PP(16'h19222,4);
TASK_PP(16'h19223,4);
TASK_PP(16'h19224,4);
TASK_PP(16'h19225,4);
TASK_PP(16'h19226,4);
TASK_PP(16'h19227,4);
TASK_PP(16'h19228,4);
TASK_PP(16'h19229,4);
TASK_PP(16'h1922A,4);
TASK_PP(16'h1922B,4);
TASK_PP(16'h1922C,4);
TASK_PP(16'h1922D,4);
TASK_PP(16'h1922E,4);
TASK_PP(16'h1922F,4);
TASK_PP(16'h19230,4);
TASK_PP(16'h19231,4);
TASK_PP(16'h19232,4);
TASK_PP(16'h19233,4);
TASK_PP(16'h19234,4);
TASK_PP(16'h19235,4);
TASK_PP(16'h19236,4);
TASK_PP(16'h19237,4);
TASK_PP(16'h19238,4);
TASK_PP(16'h19239,4);
TASK_PP(16'h1923A,4);
TASK_PP(16'h1923B,4);
TASK_PP(16'h1923C,4);
TASK_PP(16'h1923D,4);
TASK_PP(16'h1923E,4);
TASK_PP(16'h1923F,4);
TASK_PP(16'h19240,4);
TASK_PP(16'h19241,4);
TASK_PP(16'h19242,4);
TASK_PP(16'h19243,4);
TASK_PP(16'h19244,4);
TASK_PP(16'h19245,4);
TASK_PP(16'h19246,4);
TASK_PP(16'h19247,4);
TASK_PP(16'h19248,4);
TASK_PP(16'h19249,4);
TASK_PP(16'h1924A,4);
TASK_PP(16'h1924B,4);
TASK_PP(16'h1924C,4);
TASK_PP(16'h1924D,4);
TASK_PP(16'h1924E,4);
TASK_PP(16'h1924F,4);
TASK_PP(16'h19250,4);
TASK_PP(16'h19251,4);
TASK_PP(16'h19252,4);
TASK_PP(16'h19253,4);
TASK_PP(16'h19254,4);
TASK_PP(16'h19255,4);
TASK_PP(16'h19256,4);
TASK_PP(16'h19257,4);
TASK_PP(16'h19258,4);
TASK_PP(16'h19259,4);
TASK_PP(16'h1925A,4);
TASK_PP(16'h1925B,4);
TASK_PP(16'h1925C,4);
TASK_PP(16'h1925D,4);
TASK_PP(16'h1925E,4);
TASK_PP(16'h1925F,4);
TASK_PP(16'h19260,4);
TASK_PP(16'h19261,4);
TASK_PP(16'h19262,4);
TASK_PP(16'h19263,4);
TASK_PP(16'h19264,4);
TASK_PP(16'h19265,4);
TASK_PP(16'h19266,4);
TASK_PP(16'h19267,4);
TASK_PP(16'h19268,4);
TASK_PP(16'h19269,4);
TASK_PP(16'h1926A,4);
TASK_PP(16'h1926B,4);
TASK_PP(16'h1926C,4);
TASK_PP(16'h1926D,4);
TASK_PP(16'h1926E,4);
TASK_PP(16'h1926F,4);
TASK_PP(16'h19270,4);
TASK_PP(16'h19271,4);
TASK_PP(16'h19272,4);
TASK_PP(16'h19273,4);
TASK_PP(16'h19274,4);
TASK_PP(16'h19275,4);
TASK_PP(16'h19276,4);
TASK_PP(16'h19277,4);
TASK_PP(16'h19278,4);
TASK_PP(16'h19279,4);
TASK_PP(16'h1927A,4);
TASK_PP(16'h1927B,4);
TASK_PP(16'h1927C,4);
TASK_PP(16'h1927D,4);
TASK_PP(16'h1927E,4);
TASK_PP(16'h1927F,4);
TASK_PP(16'h19280,4);
TASK_PP(16'h19281,4);
TASK_PP(16'h19282,4);
TASK_PP(16'h19283,4);
TASK_PP(16'h19284,4);
TASK_PP(16'h19285,4);
TASK_PP(16'h19286,4);
TASK_PP(16'h19287,4);
TASK_PP(16'h19288,4);
TASK_PP(16'h19289,4);
TASK_PP(16'h1928A,4);
TASK_PP(16'h1928B,4);
TASK_PP(16'h1928C,4);
TASK_PP(16'h1928D,4);
TASK_PP(16'h1928E,4);
TASK_PP(16'h1928F,4);
TASK_PP(16'h19290,4);
TASK_PP(16'h19291,4);
TASK_PP(16'h19292,4);
TASK_PP(16'h19293,4);
TASK_PP(16'h19294,4);
TASK_PP(16'h19295,4);
TASK_PP(16'h19296,4);
TASK_PP(16'h19297,4);
TASK_PP(16'h19298,4);
TASK_PP(16'h19299,4);
TASK_PP(16'h1929A,4);
TASK_PP(16'h1929B,4);
TASK_PP(16'h1929C,4);
TASK_PP(16'h1929D,4);
TASK_PP(16'h1929E,4);
TASK_PP(16'h1929F,4);
TASK_PP(16'h192A0,4);
TASK_PP(16'h192A1,4);
TASK_PP(16'h192A2,4);
TASK_PP(16'h192A3,4);
TASK_PP(16'h192A4,4);
TASK_PP(16'h192A5,4);
TASK_PP(16'h192A6,4);
TASK_PP(16'h192A7,4);
TASK_PP(16'h192A8,4);
TASK_PP(16'h192A9,4);
TASK_PP(16'h192AA,4);
TASK_PP(16'h192AB,4);
TASK_PP(16'h192AC,4);
TASK_PP(16'h192AD,4);
TASK_PP(16'h192AE,4);
TASK_PP(16'h192AF,4);
TASK_PP(16'h192B0,4);
TASK_PP(16'h192B1,4);
TASK_PP(16'h192B2,4);
TASK_PP(16'h192B3,4);
TASK_PP(16'h192B4,4);
TASK_PP(16'h192B5,4);
TASK_PP(16'h192B6,4);
TASK_PP(16'h192B7,4);
TASK_PP(16'h192B8,4);
TASK_PP(16'h192B9,4);
TASK_PP(16'h192BA,4);
TASK_PP(16'h192BB,4);
TASK_PP(16'h192BC,4);
TASK_PP(16'h192BD,4);
TASK_PP(16'h192BE,4);
TASK_PP(16'h192BF,4);
TASK_PP(16'h192C0,4);
TASK_PP(16'h192C1,4);
TASK_PP(16'h192C2,4);
TASK_PP(16'h192C3,4);
TASK_PP(16'h192C4,4);
TASK_PP(16'h192C5,4);
TASK_PP(16'h192C6,4);
TASK_PP(16'h192C7,4);
TASK_PP(16'h192C8,4);
TASK_PP(16'h192C9,4);
TASK_PP(16'h192CA,4);
TASK_PP(16'h192CB,4);
TASK_PP(16'h192CC,4);
TASK_PP(16'h192CD,4);
TASK_PP(16'h192CE,4);
TASK_PP(16'h192CF,4);
TASK_PP(16'h192D0,4);
TASK_PP(16'h192D1,4);
TASK_PP(16'h192D2,4);
TASK_PP(16'h192D3,4);
TASK_PP(16'h192D4,4);
TASK_PP(16'h192D5,4);
TASK_PP(16'h192D6,4);
TASK_PP(16'h192D7,4);
TASK_PP(16'h192D8,4);
TASK_PP(16'h192D9,4);
TASK_PP(16'h192DA,4);
TASK_PP(16'h192DB,4);
TASK_PP(16'h192DC,4);
TASK_PP(16'h192DD,4);
TASK_PP(16'h192DE,4);
TASK_PP(16'h192DF,4);
TASK_PP(16'h192E0,4);
TASK_PP(16'h192E1,4);
TASK_PP(16'h192E2,4);
TASK_PP(16'h192E3,4);
TASK_PP(16'h192E4,4);
TASK_PP(16'h192E5,4);
TASK_PP(16'h192E6,4);
TASK_PP(16'h192E7,4);
TASK_PP(16'h192E8,4);
TASK_PP(16'h192E9,4);
TASK_PP(16'h192EA,4);
TASK_PP(16'h192EB,4);
TASK_PP(16'h192EC,4);
TASK_PP(16'h192ED,4);
TASK_PP(16'h192EE,4);
TASK_PP(16'h192EF,4);
TASK_PP(16'h192F0,4);
TASK_PP(16'h192F1,4);
TASK_PP(16'h192F2,4);
TASK_PP(16'h192F3,4);
TASK_PP(16'h192F4,4);
TASK_PP(16'h192F5,4);
TASK_PP(16'h192F6,4);
TASK_PP(16'h192F7,4);
TASK_PP(16'h192F8,4);
TASK_PP(16'h192F9,4);
TASK_PP(16'h192FA,4);
TASK_PP(16'h192FB,4);
TASK_PP(16'h192FC,4);
TASK_PP(16'h192FD,4);
TASK_PP(16'h192FE,4);
TASK_PP(16'h192FF,4);
TASK_PP(16'h19300,4);
TASK_PP(16'h19301,4);
TASK_PP(16'h19302,4);
TASK_PP(16'h19303,4);
TASK_PP(16'h19304,4);
TASK_PP(16'h19305,4);
TASK_PP(16'h19306,4);
TASK_PP(16'h19307,4);
TASK_PP(16'h19308,4);
TASK_PP(16'h19309,4);
TASK_PP(16'h1930A,4);
TASK_PP(16'h1930B,4);
TASK_PP(16'h1930C,4);
TASK_PP(16'h1930D,4);
TASK_PP(16'h1930E,4);
TASK_PP(16'h1930F,4);
TASK_PP(16'h19310,4);
TASK_PP(16'h19311,4);
TASK_PP(16'h19312,4);
TASK_PP(16'h19313,4);
TASK_PP(16'h19314,4);
TASK_PP(16'h19315,4);
TASK_PP(16'h19316,4);
TASK_PP(16'h19317,4);
TASK_PP(16'h19318,4);
TASK_PP(16'h19319,4);
TASK_PP(16'h1931A,4);
TASK_PP(16'h1931B,4);
TASK_PP(16'h1931C,4);
TASK_PP(16'h1931D,4);
TASK_PP(16'h1931E,4);
TASK_PP(16'h1931F,4);
TASK_PP(16'h19320,4);
TASK_PP(16'h19321,4);
TASK_PP(16'h19322,4);
TASK_PP(16'h19323,4);
TASK_PP(16'h19324,4);
TASK_PP(16'h19325,4);
TASK_PP(16'h19326,4);
TASK_PP(16'h19327,4);
TASK_PP(16'h19328,4);
TASK_PP(16'h19329,4);
TASK_PP(16'h1932A,4);
TASK_PP(16'h1932B,4);
TASK_PP(16'h1932C,4);
TASK_PP(16'h1932D,4);
TASK_PP(16'h1932E,4);
TASK_PP(16'h1932F,4);
TASK_PP(16'h19330,4);
TASK_PP(16'h19331,4);
TASK_PP(16'h19332,4);
TASK_PP(16'h19333,4);
TASK_PP(16'h19334,4);
TASK_PP(16'h19335,4);
TASK_PP(16'h19336,4);
TASK_PP(16'h19337,4);
TASK_PP(16'h19338,4);
TASK_PP(16'h19339,4);
TASK_PP(16'h1933A,4);
TASK_PP(16'h1933B,4);
TASK_PP(16'h1933C,4);
TASK_PP(16'h1933D,4);
TASK_PP(16'h1933E,4);
TASK_PP(16'h1933F,4);
TASK_PP(16'h19340,4);
TASK_PP(16'h19341,4);
TASK_PP(16'h19342,4);
TASK_PP(16'h19343,4);
TASK_PP(16'h19344,4);
TASK_PP(16'h19345,4);
TASK_PP(16'h19346,4);
TASK_PP(16'h19347,4);
TASK_PP(16'h19348,4);
TASK_PP(16'h19349,4);
TASK_PP(16'h1934A,4);
TASK_PP(16'h1934B,4);
TASK_PP(16'h1934C,4);
TASK_PP(16'h1934D,4);
TASK_PP(16'h1934E,4);
TASK_PP(16'h1934F,4);
TASK_PP(16'h19350,4);
TASK_PP(16'h19351,4);
TASK_PP(16'h19352,4);
TASK_PP(16'h19353,4);
TASK_PP(16'h19354,4);
TASK_PP(16'h19355,4);
TASK_PP(16'h19356,4);
TASK_PP(16'h19357,4);
TASK_PP(16'h19358,4);
TASK_PP(16'h19359,4);
TASK_PP(16'h1935A,4);
TASK_PP(16'h1935B,4);
TASK_PP(16'h1935C,4);
TASK_PP(16'h1935D,4);
TASK_PP(16'h1935E,4);
TASK_PP(16'h1935F,4);
TASK_PP(16'h19360,4);
TASK_PP(16'h19361,4);
TASK_PP(16'h19362,4);
TASK_PP(16'h19363,4);
TASK_PP(16'h19364,4);
TASK_PP(16'h19365,4);
TASK_PP(16'h19366,4);
TASK_PP(16'h19367,4);
TASK_PP(16'h19368,4);
TASK_PP(16'h19369,4);
TASK_PP(16'h1936A,4);
TASK_PP(16'h1936B,4);
TASK_PP(16'h1936C,4);
TASK_PP(16'h1936D,4);
TASK_PP(16'h1936E,4);
TASK_PP(16'h1936F,4);
TASK_PP(16'h19370,4);
TASK_PP(16'h19371,4);
TASK_PP(16'h19372,4);
TASK_PP(16'h19373,4);
TASK_PP(16'h19374,4);
TASK_PP(16'h19375,4);
TASK_PP(16'h19376,4);
TASK_PP(16'h19377,4);
TASK_PP(16'h19378,4);
TASK_PP(16'h19379,4);
TASK_PP(16'h1937A,4);
TASK_PP(16'h1937B,4);
TASK_PP(16'h1937C,4);
TASK_PP(16'h1937D,4);
TASK_PP(16'h1937E,4);
TASK_PP(16'h1937F,4);
TASK_PP(16'h19380,4);
TASK_PP(16'h19381,4);
TASK_PP(16'h19382,4);
TASK_PP(16'h19383,4);
TASK_PP(16'h19384,4);
TASK_PP(16'h19385,4);
TASK_PP(16'h19386,4);
TASK_PP(16'h19387,4);
TASK_PP(16'h19388,4);
TASK_PP(16'h19389,4);
TASK_PP(16'h1938A,4);
TASK_PP(16'h1938B,4);
TASK_PP(16'h1938C,4);
TASK_PP(16'h1938D,4);
TASK_PP(16'h1938E,4);
TASK_PP(16'h1938F,4);
TASK_PP(16'h19390,4);
TASK_PP(16'h19391,4);
TASK_PP(16'h19392,4);
TASK_PP(16'h19393,4);
TASK_PP(16'h19394,4);
TASK_PP(16'h19395,4);
TASK_PP(16'h19396,4);
TASK_PP(16'h19397,4);
TASK_PP(16'h19398,4);
TASK_PP(16'h19399,4);
TASK_PP(16'h1939A,4);
TASK_PP(16'h1939B,4);
TASK_PP(16'h1939C,4);
TASK_PP(16'h1939D,4);
TASK_PP(16'h1939E,4);
TASK_PP(16'h1939F,4);
TASK_PP(16'h193A0,4);
TASK_PP(16'h193A1,4);
TASK_PP(16'h193A2,4);
TASK_PP(16'h193A3,4);
TASK_PP(16'h193A4,4);
TASK_PP(16'h193A5,4);
TASK_PP(16'h193A6,4);
TASK_PP(16'h193A7,4);
TASK_PP(16'h193A8,4);
TASK_PP(16'h193A9,4);
TASK_PP(16'h193AA,4);
TASK_PP(16'h193AB,4);
TASK_PP(16'h193AC,4);
TASK_PP(16'h193AD,4);
TASK_PP(16'h193AE,4);
TASK_PP(16'h193AF,4);
TASK_PP(16'h193B0,4);
TASK_PP(16'h193B1,4);
TASK_PP(16'h193B2,4);
TASK_PP(16'h193B3,4);
TASK_PP(16'h193B4,4);
TASK_PP(16'h193B5,4);
TASK_PP(16'h193B6,4);
TASK_PP(16'h193B7,4);
TASK_PP(16'h193B8,4);
TASK_PP(16'h193B9,4);
TASK_PP(16'h193BA,4);
TASK_PP(16'h193BB,4);
TASK_PP(16'h193BC,4);
TASK_PP(16'h193BD,4);
TASK_PP(16'h193BE,4);
TASK_PP(16'h193BF,4);
TASK_PP(16'h193C0,4);
TASK_PP(16'h193C1,4);
TASK_PP(16'h193C2,4);
TASK_PP(16'h193C3,4);
TASK_PP(16'h193C4,4);
TASK_PP(16'h193C5,4);
TASK_PP(16'h193C6,4);
TASK_PP(16'h193C7,4);
TASK_PP(16'h193C8,4);
TASK_PP(16'h193C9,4);
TASK_PP(16'h193CA,4);
TASK_PP(16'h193CB,4);
TASK_PP(16'h193CC,4);
TASK_PP(16'h193CD,4);
TASK_PP(16'h193CE,4);
TASK_PP(16'h193CF,4);
TASK_PP(16'h193D0,4);
TASK_PP(16'h193D1,4);
TASK_PP(16'h193D2,4);
TASK_PP(16'h193D3,4);
TASK_PP(16'h193D4,4);
TASK_PP(16'h193D5,4);
TASK_PP(16'h193D6,4);
TASK_PP(16'h193D7,4);
TASK_PP(16'h193D8,4);
TASK_PP(16'h193D9,4);
TASK_PP(16'h193DA,4);
TASK_PP(16'h193DB,4);
TASK_PP(16'h193DC,4);
TASK_PP(16'h193DD,4);
TASK_PP(16'h193DE,4);
TASK_PP(16'h193DF,4);
TASK_PP(16'h193E0,4);
TASK_PP(16'h193E1,4);
TASK_PP(16'h193E2,4);
TASK_PP(16'h193E3,4);
TASK_PP(16'h193E4,4);
TASK_PP(16'h193E5,4);
TASK_PP(16'h193E6,4);
TASK_PP(16'h193E7,4);
TASK_PP(16'h193E8,4);
TASK_PP(16'h193E9,4);
TASK_PP(16'h193EA,4);
TASK_PP(16'h193EB,4);
TASK_PP(16'h193EC,4);
TASK_PP(16'h193ED,4);
TASK_PP(16'h193EE,4);
TASK_PP(16'h193EF,4);
TASK_PP(16'h193F0,4);
TASK_PP(16'h193F1,4);
TASK_PP(16'h193F2,4);
TASK_PP(16'h193F3,4);
TASK_PP(16'h193F4,4);
TASK_PP(16'h193F5,4);
TASK_PP(16'h193F6,4);
TASK_PP(16'h193F7,4);
TASK_PP(16'h193F8,4);
TASK_PP(16'h193F9,4);
TASK_PP(16'h193FA,4);
TASK_PP(16'h193FB,4);
TASK_PP(16'h193FC,4);
TASK_PP(16'h193FD,4);
TASK_PP(16'h193FE,4);
TASK_PP(16'h193FF,4);
TASK_PP(16'h19400,4);
TASK_PP(16'h19401,4);
TASK_PP(16'h19402,4);
TASK_PP(16'h19403,4);
TASK_PP(16'h19404,4);
TASK_PP(16'h19405,4);
TASK_PP(16'h19406,4);
TASK_PP(16'h19407,4);
TASK_PP(16'h19408,4);
TASK_PP(16'h19409,4);
TASK_PP(16'h1940A,4);
TASK_PP(16'h1940B,4);
TASK_PP(16'h1940C,4);
TASK_PP(16'h1940D,4);
TASK_PP(16'h1940E,4);
TASK_PP(16'h1940F,4);
TASK_PP(16'h19410,4);
TASK_PP(16'h19411,4);
TASK_PP(16'h19412,4);
TASK_PP(16'h19413,4);
TASK_PP(16'h19414,4);
TASK_PP(16'h19415,4);
TASK_PP(16'h19416,4);
TASK_PP(16'h19417,4);
TASK_PP(16'h19418,4);
TASK_PP(16'h19419,4);
TASK_PP(16'h1941A,4);
TASK_PP(16'h1941B,4);
TASK_PP(16'h1941C,4);
TASK_PP(16'h1941D,4);
TASK_PP(16'h1941E,4);
TASK_PP(16'h1941F,4);
TASK_PP(16'h19420,4);
TASK_PP(16'h19421,4);
TASK_PP(16'h19422,4);
TASK_PP(16'h19423,4);
TASK_PP(16'h19424,4);
TASK_PP(16'h19425,4);
TASK_PP(16'h19426,4);
TASK_PP(16'h19427,4);
TASK_PP(16'h19428,4);
TASK_PP(16'h19429,4);
TASK_PP(16'h1942A,4);
TASK_PP(16'h1942B,4);
TASK_PP(16'h1942C,4);
TASK_PP(16'h1942D,4);
TASK_PP(16'h1942E,4);
TASK_PP(16'h1942F,4);
TASK_PP(16'h19430,4);
TASK_PP(16'h19431,4);
TASK_PP(16'h19432,4);
TASK_PP(16'h19433,4);
TASK_PP(16'h19434,4);
TASK_PP(16'h19435,4);
TASK_PP(16'h19436,4);
TASK_PP(16'h19437,4);
TASK_PP(16'h19438,4);
TASK_PP(16'h19439,4);
TASK_PP(16'h1943A,4);
TASK_PP(16'h1943B,4);
TASK_PP(16'h1943C,4);
TASK_PP(16'h1943D,4);
TASK_PP(16'h1943E,4);
TASK_PP(16'h1943F,4);
TASK_PP(16'h19440,4);
TASK_PP(16'h19441,4);
TASK_PP(16'h19442,4);
TASK_PP(16'h19443,4);
TASK_PP(16'h19444,4);
TASK_PP(16'h19445,4);
TASK_PP(16'h19446,4);
TASK_PP(16'h19447,4);
TASK_PP(16'h19448,4);
TASK_PP(16'h19449,4);
TASK_PP(16'h1944A,4);
TASK_PP(16'h1944B,4);
TASK_PP(16'h1944C,4);
TASK_PP(16'h1944D,4);
TASK_PP(16'h1944E,4);
TASK_PP(16'h1944F,4);
TASK_PP(16'h19450,4);
TASK_PP(16'h19451,4);
TASK_PP(16'h19452,4);
TASK_PP(16'h19453,4);
TASK_PP(16'h19454,4);
TASK_PP(16'h19455,4);
TASK_PP(16'h19456,4);
TASK_PP(16'h19457,4);
TASK_PP(16'h19458,4);
TASK_PP(16'h19459,4);
TASK_PP(16'h1945A,4);
TASK_PP(16'h1945B,4);
TASK_PP(16'h1945C,4);
TASK_PP(16'h1945D,4);
TASK_PP(16'h1945E,4);
TASK_PP(16'h1945F,4);
TASK_PP(16'h19460,4);
TASK_PP(16'h19461,4);
TASK_PP(16'h19462,4);
TASK_PP(16'h19463,4);
TASK_PP(16'h19464,4);
TASK_PP(16'h19465,4);
TASK_PP(16'h19466,4);
TASK_PP(16'h19467,4);
TASK_PP(16'h19468,4);
TASK_PP(16'h19469,4);
TASK_PP(16'h1946A,4);
TASK_PP(16'h1946B,4);
TASK_PP(16'h1946C,4);
TASK_PP(16'h1946D,4);
TASK_PP(16'h1946E,4);
TASK_PP(16'h1946F,4);
TASK_PP(16'h19470,4);
TASK_PP(16'h19471,4);
TASK_PP(16'h19472,4);
TASK_PP(16'h19473,4);
TASK_PP(16'h19474,4);
TASK_PP(16'h19475,4);
TASK_PP(16'h19476,4);
TASK_PP(16'h19477,4);
TASK_PP(16'h19478,4);
TASK_PP(16'h19479,4);
TASK_PP(16'h1947A,4);
TASK_PP(16'h1947B,4);
TASK_PP(16'h1947C,4);
TASK_PP(16'h1947D,4);
TASK_PP(16'h1947E,4);
TASK_PP(16'h1947F,4);
TASK_PP(16'h19480,4);
TASK_PP(16'h19481,4);
TASK_PP(16'h19482,4);
TASK_PP(16'h19483,4);
TASK_PP(16'h19484,4);
TASK_PP(16'h19485,4);
TASK_PP(16'h19486,4);
TASK_PP(16'h19487,4);
TASK_PP(16'h19488,4);
TASK_PP(16'h19489,4);
TASK_PP(16'h1948A,4);
TASK_PP(16'h1948B,4);
TASK_PP(16'h1948C,4);
TASK_PP(16'h1948D,4);
TASK_PP(16'h1948E,4);
TASK_PP(16'h1948F,4);
TASK_PP(16'h19490,4);
TASK_PP(16'h19491,4);
TASK_PP(16'h19492,4);
TASK_PP(16'h19493,4);
TASK_PP(16'h19494,4);
TASK_PP(16'h19495,4);
TASK_PP(16'h19496,4);
TASK_PP(16'h19497,4);
TASK_PP(16'h19498,4);
TASK_PP(16'h19499,4);
TASK_PP(16'h1949A,4);
TASK_PP(16'h1949B,4);
TASK_PP(16'h1949C,4);
TASK_PP(16'h1949D,4);
TASK_PP(16'h1949E,4);
TASK_PP(16'h1949F,4);
TASK_PP(16'h194A0,4);
TASK_PP(16'h194A1,4);
TASK_PP(16'h194A2,4);
TASK_PP(16'h194A3,4);
TASK_PP(16'h194A4,4);
TASK_PP(16'h194A5,4);
TASK_PP(16'h194A6,4);
TASK_PP(16'h194A7,4);
TASK_PP(16'h194A8,4);
TASK_PP(16'h194A9,4);
TASK_PP(16'h194AA,4);
TASK_PP(16'h194AB,4);
TASK_PP(16'h194AC,4);
TASK_PP(16'h194AD,4);
TASK_PP(16'h194AE,4);
TASK_PP(16'h194AF,4);
TASK_PP(16'h194B0,4);
TASK_PP(16'h194B1,4);
TASK_PP(16'h194B2,4);
TASK_PP(16'h194B3,4);
TASK_PP(16'h194B4,4);
TASK_PP(16'h194B5,4);
TASK_PP(16'h194B6,4);
TASK_PP(16'h194B7,4);
TASK_PP(16'h194B8,4);
TASK_PP(16'h194B9,4);
TASK_PP(16'h194BA,4);
TASK_PP(16'h194BB,4);
TASK_PP(16'h194BC,4);
TASK_PP(16'h194BD,4);
TASK_PP(16'h194BE,4);
TASK_PP(16'h194BF,4);
TASK_PP(16'h194C0,4);
TASK_PP(16'h194C1,4);
TASK_PP(16'h194C2,4);
TASK_PP(16'h194C3,4);
TASK_PP(16'h194C4,4);
TASK_PP(16'h194C5,4);
TASK_PP(16'h194C6,4);
TASK_PP(16'h194C7,4);
TASK_PP(16'h194C8,4);
TASK_PP(16'h194C9,4);
TASK_PP(16'h194CA,4);
TASK_PP(16'h194CB,4);
TASK_PP(16'h194CC,4);
TASK_PP(16'h194CD,4);
TASK_PP(16'h194CE,4);
TASK_PP(16'h194CF,4);
TASK_PP(16'h194D0,4);
TASK_PP(16'h194D1,4);
TASK_PP(16'h194D2,4);
TASK_PP(16'h194D3,4);
TASK_PP(16'h194D4,4);
TASK_PP(16'h194D5,4);
TASK_PP(16'h194D6,4);
TASK_PP(16'h194D7,4);
TASK_PP(16'h194D8,4);
TASK_PP(16'h194D9,4);
TASK_PP(16'h194DA,4);
TASK_PP(16'h194DB,4);
TASK_PP(16'h194DC,4);
TASK_PP(16'h194DD,4);
TASK_PP(16'h194DE,4);
TASK_PP(16'h194DF,4);
TASK_PP(16'h194E0,4);
TASK_PP(16'h194E1,4);
TASK_PP(16'h194E2,4);
TASK_PP(16'h194E3,4);
TASK_PP(16'h194E4,4);
TASK_PP(16'h194E5,4);
TASK_PP(16'h194E6,4);
TASK_PP(16'h194E7,4);
TASK_PP(16'h194E8,4);
TASK_PP(16'h194E9,4);
TASK_PP(16'h194EA,4);
TASK_PP(16'h194EB,4);
TASK_PP(16'h194EC,4);
TASK_PP(16'h194ED,4);
TASK_PP(16'h194EE,4);
TASK_PP(16'h194EF,4);
TASK_PP(16'h194F0,4);
TASK_PP(16'h194F1,4);
TASK_PP(16'h194F2,4);
TASK_PP(16'h194F3,4);
TASK_PP(16'h194F4,4);
TASK_PP(16'h194F5,4);
TASK_PP(16'h194F6,4);
TASK_PP(16'h194F7,4);
TASK_PP(16'h194F8,4);
TASK_PP(16'h194F9,4);
TASK_PP(16'h194FA,4);
TASK_PP(16'h194FB,4);
TASK_PP(16'h194FC,4);
TASK_PP(16'h194FD,4);
TASK_PP(16'h194FE,4);
TASK_PP(16'h194FF,4);
TASK_PP(16'h19500,4);
TASK_PP(16'h19501,4);
TASK_PP(16'h19502,4);
TASK_PP(16'h19503,4);
TASK_PP(16'h19504,4);
TASK_PP(16'h19505,4);
TASK_PP(16'h19506,4);
TASK_PP(16'h19507,4);
TASK_PP(16'h19508,4);
TASK_PP(16'h19509,4);
TASK_PP(16'h1950A,4);
TASK_PP(16'h1950B,4);
TASK_PP(16'h1950C,4);
TASK_PP(16'h1950D,4);
TASK_PP(16'h1950E,4);
TASK_PP(16'h1950F,4);
TASK_PP(16'h19510,4);
TASK_PP(16'h19511,4);
TASK_PP(16'h19512,4);
TASK_PP(16'h19513,4);
TASK_PP(16'h19514,4);
TASK_PP(16'h19515,4);
TASK_PP(16'h19516,4);
TASK_PP(16'h19517,4);
TASK_PP(16'h19518,4);
TASK_PP(16'h19519,4);
TASK_PP(16'h1951A,4);
TASK_PP(16'h1951B,4);
TASK_PP(16'h1951C,4);
TASK_PP(16'h1951D,4);
TASK_PP(16'h1951E,4);
TASK_PP(16'h1951F,4);
TASK_PP(16'h19520,4);
TASK_PP(16'h19521,4);
TASK_PP(16'h19522,4);
TASK_PP(16'h19523,4);
TASK_PP(16'h19524,4);
TASK_PP(16'h19525,4);
TASK_PP(16'h19526,4);
TASK_PP(16'h19527,4);
TASK_PP(16'h19528,4);
TASK_PP(16'h19529,4);
TASK_PP(16'h1952A,4);
TASK_PP(16'h1952B,4);
TASK_PP(16'h1952C,4);
TASK_PP(16'h1952D,4);
TASK_PP(16'h1952E,4);
TASK_PP(16'h1952F,4);
TASK_PP(16'h19530,4);
TASK_PP(16'h19531,4);
TASK_PP(16'h19532,4);
TASK_PP(16'h19533,4);
TASK_PP(16'h19534,4);
TASK_PP(16'h19535,4);
TASK_PP(16'h19536,4);
TASK_PP(16'h19537,4);
TASK_PP(16'h19538,4);
TASK_PP(16'h19539,4);
TASK_PP(16'h1953A,4);
TASK_PP(16'h1953B,4);
TASK_PP(16'h1953C,4);
TASK_PP(16'h1953D,4);
TASK_PP(16'h1953E,4);
TASK_PP(16'h1953F,4);
TASK_PP(16'h19540,4);
TASK_PP(16'h19541,4);
TASK_PP(16'h19542,4);
TASK_PP(16'h19543,4);
TASK_PP(16'h19544,4);
TASK_PP(16'h19545,4);
TASK_PP(16'h19546,4);
TASK_PP(16'h19547,4);
TASK_PP(16'h19548,4);
TASK_PP(16'h19549,4);
TASK_PP(16'h1954A,4);
TASK_PP(16'h1954B,4);
TASK_PP(16'h1954C,4);
TASK_PP(16'h1954D,4);
TASK_PP(16'h1954E,4);
TASK_PP(16'h1954F,4);
TASK_PP(16'h19550,4);
TASK_PP(16'h19551,4);
TASK_PP(16'h19552,4);
TASK_PP(16'h19553,4);
TASK_PP(16'h19554,4);
TASK_PP(16'h19555,4);
TASK_PP(16'h19556,4);
TASK_PP(16'h19557,4);
TASK_PP(16'h19558,4);
TASK_PP(16'h19559,4);
TASK_PP(16'h1955A,4);
TASK_PP(16'h1955B,4);
TASK_PP(16'h1955C,4);
TASK_PP(16'h1955D,4);
TASK_PP(16'h1955E,4);
TASK_PP(16'h1955F,4);
TASK_PP(16'h19560,4);
TASK_PP(16'h19561,4);
TASK_PP(16'h19562,4);
TASK_PP(16'h19563,4);
TASK_PP(16'h19564,4);
TASK_PP(16'h19565,4);
TASK_PP(16'h19566,4);
TASK_PP(16'h19567,4);
TASK_PP(16'h19568,4);
TASK_PP(16'h19569,4);
TASK_PP(16'h1956A,4);
TASK_PP(16'h1956B,4);
TASK_PP(16'h1956C,4);
TASK_PP(16'h1956D,4);
TASK_PP(16'h1956E,4);
TASK_PP(16'h1956F,4);
TASK_PP(16'h19570,4);
TASK_PP(16'h19571,4);
TASK_PP(16'h19572,4);
TASK_PP(16'h19573,4);
TASK_PP(16'h19574,4);
TASK_PP(16'h19575,4);
TASK_PP(16'h19576,4);
TASK_PP(16'h19577,4);
TASK_PP(16'h19578,4);
TASK_PP(16'h19579,4);
TASK_PP(16'h1957A,4);
TASK_PP(16'h1957B,4);
TASK_PP(16'h1957C,4);
TASK_PP(16'h1957D,4);
TASK_PP(16'h1957E,4);
TASK_PP(16'h1957F,4);
TASK_PP(16'h19580,4);
TASK_PP(16'h19581,4);
TASK_PP(16'h19582,4);
TASK_PP(16'h19583,4);
TASK_PP(16'h19584,4);
TASK_PP(16'h19585,4);
TASK_PP(16'h19586,4);
TASK_PP(16'h19587,4);
TASK_PP(16'h19588,4);
TASK_PP(16'h19589,4);
TASK_PP(16'h1958A,4);
TASK_PP(16'h1958B,4);
TASK_PP(16'h1958C,4);
TASK_PP(16'h1958D,4);
TASK_PP(16'h1958E,4);
TASK_PP(16'h1958F,4);
TASK_PP(16'h19590,4);
TASK_PP(16'h19591,4);
TASK_PP(16'h19592,4);
TASK_PP(16'h19593,4);
TASK_PP(16'h19594,4);
TASK_PP(16'h19595,4);
TASK_PP(16'h19596,4);
TASK_PP(16'h19597,4);
TASK_PP(16'h19598,4);
TASK_PP(16'h19599,4);
TASK_PP(16'h1959A,4);
TASK_PP(16'h1959B,4);
TASK_PP(16'h1959C,4);
TASK_PP(16'h1959D,4);
TASK_PP(16'h1959E,4);
TASK_PP(16'h1959F,4);
TASK_PP(16'h195A0,4);
TASK_PP(16'h195A1,4);
TASK_PP(16'h195A2,4);
TASK_PP(16'h195A3,4);
TASK_PP(16'h195A4,4);
TASK_PP(16'h195A5,4);
TASK_PP(16'h195A6,4);
TASK_PP(16'h195A7,4);
TASK_PP(16'h195A8,4);
TASK_PP(16'h195A9,4);
TASK_PP(16'h195AA,4);
TASK_PP(16'h195AB,4);
TASK_PP(16'h195AC,4);
TASK_PP(16'h195AD,4);
TASK_PP(16'h195AE,4);
TASK_PP(16'h195AF,4);
TASK_PP(16'h195B0,4);
TASK_PP(16'h195B1,4);
TASK_PP(16'h195B2,4);
TASK_PP(16'h195B3,4);
TASK_PP(16'h195B4,4);
TASK_PP(16'h195B5,4);
TASK_PP(16'h195B6,4);
TASK_PP(16'h195B7,4);
TASK_PP(16'h195B8,4);
TASK_PP(16'h195B9,4);
TASK_PP(16'h195BA,4);
TASK_PP(16'h195BB,4);
TASK_PP(16'h195BC,4);
TASK_PP(16'h195BD,4);
TASK_PP(16'h195BE,4);
TASK_PP(16'h195BF,4);
TASK_PP(16'h195C0,4);
TASK_PP(16'h195C1,4);
TASK_PP(16'h195C2,4);
TASK_PP(16'h195C3,4);
TASK_PP(16'h195C4,4);
TASK_PP(16'h195C5,4);
TASK_PP(16'h195C6,4);
TASK_PP(16'h195C7,4);
TASK_PP(16'h195C8,4);
TASK_PP(16'h195C9,4);
TASK_PP(16'h195CA,4);
TASK_PP(16'h195CB,4);
TASK_PP(16'h195CC,4);
TASK_PP(16'h195CD,4);
TASK_PP(16'h195CE,4);
TASK_PP(16'h195CF,4);
TASK_PP(16'h195D0,4);
TASK_PP(16'h195D1,4);
TASK_PP(16'h195D2,4);
TASK_PP(16'h195D3,4);
TASK_PP(16'h195D4,4);
TASK_PP(16'h195D5,4);
TASK_PP(16'h195D6,4);
TASK_PP(16'h195D7,4);
TASK_PP(16'h195D8,4);
TASK_PP(16'h195D9,4);
TASK_PP(16'h195DA,4);
TASK_PP(16'h195DB,4);
TASK_PP(16'h195DC,4);
TASK_PP(16'h195DD,4);
TASK_PP(16'h195DE,4);
TASK_PP(16'h195DF,4);
TASK_PP(16'h195E0,4);
TASK_PP(16'h195E1,4);
TASK_PP(16'h195E2,4);
TASK_PP(16'h195E3,4);
TASK_PP(16'h195E4,4);
TASK_PP(16'h195E5,4);
TASK_PP(16'h195E6,4);
TASK_PP(16'h195E7,4);
TASK_PP(16'h195E8,4);
TASK_PP(16'h195E9,4);
TASK_PP(16'h195EA,4);
TASK_PP(16'h195EB,4);
TASK_PP(16'h195EC,4);
TASK_PP(16'h195ED,4);
TASK_PP(16'h195EE,4);
TASK_PP(16'h195EF,4);
TASK_PP(16'h195F0,4);
TASK_PP(16'h195F1,4);
TASK_PP(16'h195F2,4);
TASK_PP(16'h195F3,4);
TASK_PP(16'h195F4,4);
TASK_PP(16'h195F5,4);
TASK_PP(16'h195F6,4);
TASK_PP(16'h195F7,4);
TASK_PP(16'h195F8,4);
TASK_PP(16'h195F9,4);
TASK_PP(16'h195FA,4);
TASK_PP(16'h195FB,4);
TASK_PP(16'h195FC,4);
TASK_PP(16'h195FD,4);
TASK_PP(16'h195FE,4);
TASK_PP(16'h195FF,4);
TASK_PP(16'h19600,4);
TASK_PP(16'h19601,4);
TASK_PP(16'h19602,4);
TASK_PP(16'h19603,4);
TASK_PP(16'h19604,4);
TASK_PP(16'h19605,4);
TASK_PP(16'h19606,4);
TASK_PP(16'h19607,4);
TASK_PP(16'h19608,4);
TASK_PP(16'h19609,4);
TASK_PP(16'h1960A,4);
TASK_PP(16'h1960B,4);
TASK_PP(16'h1960C,4);
TASK_PP(16'h1960D,4);
TASK_PP(16'h1960E,4);
TASK_PP(16'h1960F,4);
TASK_PP(16'h19610,4);
TASK_PP(16'h19611,4);
TASK_PP(16'h19612,4);
TASK_PP(16'h19613,4);
TASK_PP(16'h19614,4);
TASK_PP(16'h19615,4);
TASK_PP(16'h19616,4);
TASK_PP(16'h19617,4);
TASK_PP(16'h19618,4);
TASK_PP(16'h19619,4);
TASK_PP(16'h1961A,4);
TASK_PP(16'h1961B,4);
TASK_PP(16'h1961C,4);
TASK_PP(16'h1961D,4);
TASK_PP(16'h1961E,4);
TASK_PP(16'h1961F,4);
TASK_PP(16'h19620,4);
TASK_PP(16'h19621,4);
TASK_PP(16'h19622,4);
TASK_PP(16'h19623,4);
TASK_PP(16'h19624,4);
TASK_PP(16'h19625,4);
TASK_PP(16'h19626,4);
TASK_PP(16'h19627,4);
TASK_PP(16'h19628,4);
TASK_PP(16'h19629,4);
TASK_PP(16'h1962A,4);
TASK_PP(16'h1962B,4);
TASK_PP(16'h1962C,4);
TASK_PP(16'h1962D,4);
TASK_PP(16'h1962E,4);
TASK_PP(16'h1962F,4);
TASK_PP(16'h19630,4);
TASK_PP(16'h19631,4);
TASK_PP(16'h19632,4);
TASK_PP(16'h19633,4);
TASK_PP(16'h19634,4);
TASK_PP(16'h19635,4);
TASK_PP(16'h19636,4);
TASK_PP(16'h19637,4);
TASK_PP(16'h19638,4);
TASK_PP(16'h19639,4);
TASK_PP(16'h1963A,4);
TASK_PP(16'h1963B,4);
TASK_PP(16'h1963C,4);
TASK_PP(16'h1963D,4);
TASK_PP(16'h1963E,4);
TASK_PP(16'h1963F,4);
TASK_PP(16'h19640,4);
TASK_PP(16'h19641,4);
TASK_PP(16'h19642,4);
TASK_PP(16'h19643,4);
TASK_PP(16'h19644,4);
TASK_PP(16'h19645,4);
TASK_PP(16'h19646,4);
TASK_PP(16'h19647,4);
TASK_PP(16'h19648,4);
TASK_PP(16'h19649,4);
TASK_PP(16'h1964A,4);
TASK_PP(16'h1964B,4);
TASK_PP(16'h1964C,4);
TASK_PP(16'h1964D,4);
TASK_PP(16'h1964E,4);
TASK_PP(16'h1964F,4);
TASK_PP(16'h19650,4);
TASK_PP(16'h19651,4);
TASK_PP(16'h19652,4);
TASK_PP(16'h19653,4);
TASK_PP(16'h19654,4);
TASK_PP(16'h19655,4);
TASK_PP(16'h19656,4);
TASK_PP(16'h19657,4);
TASK_PP(16'h19658,4);
TASK_PP(16'h19659,4);
TASK_PP(16'h1965A,4);
TASK_PP(16'h1965B,4);
TASK_PP(16'h1965C,4);
TASK_PP(16'h1965D,4);
TASK_PP(16'h1965E,4);
TASK_PP(16'h1965F,4);
TASK_PP(16'h19660,4);
TASK_PP(16'h19661,4);
TASK_PP(16'h19662,4);
TASK_PP(16'h19663,4);
TASK_PP(16'h19664,4);
TASK_PP(16'h19665,4);
TASK_PP(16'h19666,4);
TASK_PP(16'h19667,4);
TASK_PP(16'h19668,4);
TASK_PP(16'h19669,4);
TASK_PP(16'h1966A,4);
TASK_PP(16'h1966B,4);
TASK_PP(16'h1966C,4);
TASK_PP(16'h1966D,4);
TASK_PP(16'h1966E,4);
TASK_PP(16'h1966F,4);
TASK_PP(16'h19670,4);
TASK_PP(16'h19671,4);
TASK_PP(16'h19672,4);
TASK_PP(16'h19673,4);
TASK_PP(16'h19674,4);
TASK_PP(16'h19675,4);
TASK_PP(16'h19676,4);
TASK_PP(16'h19677,4);
TASK_PP(16'h19678,4);
TASK_PP(16'h19679,4);
TASK_PP(16'h1967A,4);
TASK_PP(16'h1967B,4);
TASK_PP(16'h1967C,4);
TASK_PP(16'h1967D,4);
TASK_PP(16'h1967E,4);
TASK_PP(16'h1967F,4);
TASK_PP(16'h19680,4);
TASK_PP(16'h19681,4);
TASK_PP(16'h19682,4);
TASK_PP(16'h19683,4);
TASK_PP(16'h19684,4);
TASK_PP(16'h19685,4);
TASK_PP(16'h19686,4);
TASK_PP(16'h19687,4);
TASK_PP(16'h19688,4);
TASK_PP(16'h19689,4);
TASK_PP(16'h1968A,4);
TASK_PP(16'h1968B,4);
TASK_PP(16'h1968C,4);
TASK_PP(16'h1968D,4);
TASK_PP(16'h1968E,4);
TASK_PP(16'h1968F,4);
TASK_PP(16'h19690,4);
TASK_PP(16'h19691,4);
TASK_PP(16'h19692,4);
TASK_PP(16'h19693,4);
TASK_PP(16'h19694,4);
TASK_PP(16'h19695,4);
TASK_PP(16'h19696,4);
TASK_PP(16'h19697,4);
TASK_PP(16'h19698,4);
TASK_PP(16'h19699,4);
TASK_PP(16'h1969A,4);
TASK_PP(16'h1969B,4);
TASK_PP(16'h1969C,4);
TASK_PP(16'h1969D,4);
TASK_PP(16'h1969E,4);
TASK_PP(16'h1969F,4);
TASK_PP(16'h196A0,4);
TASK_PP(16'h196A1,4);
TASK_PP(16'h196A2,4);
TASK_PP(16'h196A3,4);
TASK_PP(16'h196A4,4);
TASK_PP(16'h196A5,4);
TASK_PP(16'h196A6,4);
TASK_PP(16'h196A7,4);
TASK_PP(16'h196A8,4);
TASK_PP(16'h196A9,4);
TASK_PP(16'h196AA,4);
TASK_PP(16'h196AB,4);
TASK_PP(16'h196AC,4);
TASK_PP(16'h196AD,4);
TASK_PP(16'h196AE,4);
TASK_PP(16'h196AF,4);
TASK_PP(16'h196B0,4);
TASK_PP(16'h196B1,4);
TASK_PP(16'h196B2,4);
TASK_PP(16'h196B3,4);
TASK_PP(16'h196B4,4);
TASK_PP(16'h196B5,4);
TASK_PP(16'h196B6,4);
TASK_PP(16'h196B7,4);
TASK_PP(16'h196B8,4);
TASK_PP(16'h196B9,4);
TASK_PP(16'h196BA,4);
TASK_PP(16'h196BB,4);
TASK_PP(16'h196BC,4);
TASK_PP(16'h196BD,4);
TASK_PP(16'h196BE,4);
TASK_PP(16'h196BF,4);
TASK_PP(16'h196C0,4);
TASK_PP(16'h196C1,4);
TASK_PP(16'h196C2,4);
TASK_PP(16'h196C3,4);
TASK_PP(16'h196C4,4);
TASK_PP(16'h196C5,4);
TASK_PP(16'h196C6,4);
TASK_PP(16'h196C7,4);
TASK_PP(16'h196C8,4);
TASK_PP(16'h196C9,4);
TASK_PP(16'h196CA,4);
TASK_PP(16'h196CB,4);
TASK_PP(16'h196CC,4);
TASK_PP(16'h196CD,4);
TASK_PP(16'h196CE,4);
TASK_PP(16'h196CF,4);
TASK_PP(16'h196D0,4);
TASK_PP(16'h196D1,4);
TASK_PP(16'h196D2,4);
TASK_PP(16'h196D3,4);
TASK_PP(16'h196D4,4);
TASK_PP(16'h196D5,4);
TASK_PP(16'h196D6,4);
TASK_PP(16'h196D7,4);
TASK_PP(16'h196D8,4);
TASK_PP(16'h196D9,4);
TASK_PP(16'h196DA,4);
TASK_PP(16'h196DB,4);
TASK_PP(16'h196DC,4);
TASK_PP(16'h196DD,4);
TASK_PP(16'h196DE,4);
TASK_PP(16'h196DF,4);
TASK_PP(16'h196E0,4);
TASK_PP(16'h196E1,4);
TASK_PP(16'h196E2,4);
TASK_PP(16'h196E3,4);
TASK_PP(16'h196E4,4);
TASK_PP(16'h196E5,4);
TASK_PP(16'h196E6,4);
TASK_PP(16'h196E7,4);
TASK_PP(16'h196E8,4);
TASK_PP(16'h196E9,4);
TASK_PP(16'h196EA,4);
TASK_PP(16'h196EB,4);
TASK_PP(16'h196EC,4);
TASK_PP(16'h196ED,4);
TASK_PP(16'h196EE,4);
TASK_PP(16'h196EF,4);
TASK_PP(16'h196F0,4);
TASK_PP(16'h196F1,4);
TASK_PP(16'h196F2,4);
TASK_PP(16'h196F3,4);
TASK_PP(16'h196F4,4);
TASK_PP(16'h196F5,4);
TASK_PP(16'h196F6,4);
TASK_PP(16'h196F7,4);
TASK_PP(16'h196F8,4);
TASK_PP(16'h196F9,4);
TASK_PP(16'h196FA,4);
TASK_PP(16'h196FB,4);
TASK_PP(16'h196FC,4);
TASK_PP(16'h196FD,4);
TASK_PP(16'h196FE,4);
TASK_PP(16'h196FF,4);
TASK_PP(16'h19700,4);
TASK_PP(16'h19701,4);
TASK_PP(16'h19702,4);
TASK_PP(16'h19703,4);
TASK_PP(16'h19704,4);
TASK_PP(16'h19705,4);
TASK_PP(16'h19706,4);
TASK_PP(16'h19707,4);
TASK_PP(16'h19708,4);
TASK_PP(16'h19709,4);
TASK_PP(16'h1970A,4);
TASK_PP(16'h1970B,4);
TASK_PP(16'h1970C,4);
TASK_PP(16'h1970D,4);
TASK_PP(16'h1970E,4);
TASK_PP(16'h1970F,4);
TASK_PP(16'h19710,4);
TASK_PP(16'h19711,4);
TASK_PP(16'h19712,4);
TASK_PP(16'h19713,4);
TASK_PP(16'h19714,4);
TASK_PP(16'h19715,4);
TASK_PP(16'h19716,4);
TASK_PP(16'h19717,4);
TASK_PP(16'h19718,4);
TASK_PP(16'h19719,4);
TASK_PP(16'h1971A,4);
TASK_PP(16'h1971B,4);
TASK_PP(16'h1971C,4);
TASK_PP(16'h1971D,4);
TASK_PP(16'h1971E,4);
TASK_PP(16'h1971F,4);
TASK_PP(16'h19720,4);
TASK_PP(16'h19721,4);
TASK_PP(16'h19722,4);
TASK_PP(16'h19723,4);
TASK_PP(16'h19724,4);
TASK_PP(16'h19725,4);
TASK_PP(16'h19726,4);
TASK_PP(16'h19727,4);
TASK_PP(16'h19728,4);
TASK_PP(16'h19729,4);
TASK_PP(16'h1972A,4);
TASK_PP(16'h1972B,4);
TASK_PP(16'h1972C,4);
TASK_PP(16'h1972D,4);
TASK_PP(16'h1972E,4);
TASK_PP(16'h1972F,4);
TASK_PP(16'h19730,4);
TASK_PP(16'h19731,4);
TASK_PP(16'h19732,4);
TASK_PP(16'h19733,4);
TASK_PP(16'h19734,4);
TASK_PP(16'h19735,4);
TASK_PP(16'h19736,4);
TASK_PP(16'h19737,4);
TASK_PP(16'h19738,4);
TASK_PP(16'h19739,4);
TASK_PP(16'h1973A,4);
TASK_PP(16'h1973B,4);
TASK_PP(16'h1973C,4);
TASK_PP(16'h1973D,4);
TASK_PP(16'h1973E,4);
TASK_PP(16'h1973F,4);
TASK_PP(16'h19740,4);
TASK_PP(16'h19741,4);
TASK_PP(16'h19742,4);
TASK_PP(16'h19743,4);
TASK_PP(16'h19744,4);
TASK_PP(16'h19745,4);
TASK_PP(16'h19746,4);
TASK_PP(16'h19747,4);
TASK_PP(16'h19748,4);
TASK_PP(16'h19749,4);
TASK_PP(16'h1974A,4);
TASK_PP(16'h1974B,4);
TASK_PP(16'h1974C,4);
TASK_PP(16'h1974D,4);
TASK_PP(16'h1974E,4);
TASK_PP(16'h1974F,4);
TASK_PP(16'h19750,4);
TASK_PP(16'h19751,4);
TASK_PP(16'h19752,4);
TASK_PP(16'h19753,4);
TASK_PP(16'h19754,4);
TASK_PP(16'h19755,4);
TASK_PP(16'h19756,4);
TASK_PP(16'h19757,4);
TASK_PP(16'h19758,4);
TASK_PP(16'h19759,4);
TASK_PP(16'h1975A,4);
TASK_PP(16'h1975B,4);
TASK_PP(16'h1975C,4);
TASK_PP(16'h1975D,4);
TASK_PP(16'h1975E,4);
TASK_PP(16'h1975F,4);
TASK_PP(16'h19760,4);
TASK_PP(16'h19761,4);
TASK_PP(16'h19762,4);
TASK_PP(16'h19763,4);
TASK_PP(16'h19764,4);
TASK_PP(16'h19765,4);
TASK_PP(16'h19766,4);
TASK_PP(16'h19767,4);
TASK_PP(16'h19768,4);
TASK_PP(16'h19769,4);
TASK_PP(16'h1976A,4);
TASK_PP(16'h1976B,4);
TASK_PP(16'h1976C,4);
TASK_PP(16'h1976D,4);
TASK_PP(16'h1976E,4);
TASK_PP(16'h1976F,4);
TASK_PP(16'h19770,4);
TASK_PP(16'h19771,4);
TASK_PP(16'h19772,4);
TASK_PP(16'h19773,4);
TASK_PP(16'h19774,4);
TASK_PP(16'h19775,4);
TASK_PP(16'h19776,4);
TASK_PP(16'h19777,4);
TASK_PP(16'h19778,4);
TASK_PP(16'h19779,4);
TASK_PP(16'h1977A,4);
TASK_PP(16'h1977B,4);
TASK_PP(16'h1977C,4);
TASK_PP(16'h1977D,4);
TASK_PP(16'h1977E,4);
TASK_PP(16'h1977F,4);
TASK_PP(16'h19780,4);
TASK_PP(16'h19781,4);
TASK_PP(16'h19782,4);
TASK_PP(16'h19783,4);
TASK_PP(16'h19784,4);
TASK_PP(16'h19785,4);
TASK_PP(16'h19786,4);
TASK_PP(16'h19787,4);
TASK_PP(16'h19788,4);
TASK_PP(16'h19789,4);
TASK_PP(16'h1978A,4);
TASK_PP(16'h1978B,4);
TASK_PP(16'h1978C,4);
TASK_PP(16'h1978D,4);
TASK_PP(16'h1978E,4);
TASK_PP(16'h1978F,4);
TASK_PP(16'h19790,4);
TASK_PP(16'h19791,4);
TASK_PP(16'h19792,4);
TASK_PP(16'h19793,4);
TASK_PP(16'h19794,4);
TASK_PP(16'h19795,4);
TASK_PP(16'h19796,4);
TASK_PP(16'h19797,4);
TASK_PP(16'h19798,4);
TASK_PP(16'h19799,4);
TASK_PP(16'h1979A,4);
TASK_PP(16'h1979B,4);
TASK_PP(16'h1979C,4);
TASK_PP(16'h1979D,4);
TASK_PP(16'h1979E,4);
TASK_PP(16'h1979F,4);
TASK_PP(16'h197A0,4);
TASK_PP(16'h197A1,4);
TASK_PP(16'h197A2,4);
TASK_PP(16'h197A3,4);
TASK_PP(16'h197A4,4);
TASK_PP(16'h197A5,4);
TASK_PP(16'h197A6,4);
TASK_PP(16'h197A7,4);
TASK_PP(16'h197A8,4);
TASK_PP(16'h197A9,4);
TASK_PP(16'h197AA,4);
TASK_PP(16'h197AB,4);
TASK_PP(16'h197AC,4);
TASK_PP(16'h197AD,4);
TASK_PP(16'h197AE,4);
TASK_PP(16'h197AF,4);
TASK_PP(16'h197B0,4);
TASK_PP(16'h197B1,4);
TASK_PP(16'h197B2,4);
TASK_PP(16'h197B3,4);
TASK_PP(16'h197B4,4);
TASK_PP(16'h197B5,4);
TASK_PP(16'h197B6,4);
TASK_PP(16'h197B7,4);
TASK_PP(16'h197B8,4);
TASK_PP(16'h197B9,4);
TASK_PP(16'h197BA,4);
TASK_PP(16'h197BB,4);
TASK_PP(16'h197BC,4);
TASK_PP(16'h197BD,4);
TASK_PP(16'h197BE,4);
TASK_PP(16'h197BF,4);
TASK_PP(16'h197C0,4);
TASK_PP(16'h197C1,4);
TASK_PP(16'h197C2,4);
TASK_PP(16'h197C3,4);
TASK_PP(16'h197C4,4);
TASK_PP(16'h197C5,4);
TASK_PP(16'h197C6,4);
TASK_PP(16'h197C7,4);
TASK_PP(16'h197C8,4);
TASK_PP(16'h197C9,4);
TASK_PP(16'h197CA,4);
TASK_PP(16'h197CB,4);
TASK_PP(16'h197CC,4);
TASK_PP(16'h197CD,4);
TASK_PP(16'h197CE,4);
TASK_PP(16'h197CF,4);
TASK_PP(16'h197D0,4);
TASK_PP(16'h197D1,4);
TASK_PP(16'h197D2,4);
TASK_PP(16'h197D3,4);
TASK_PP(16'h197D4,4);
TASK_PP(16'h197D5,4);
TASK_PP(16'h197D6,4);
TASK_PP(16'h197D7,4);
TASK_PP(16'h197D8,4);
TASK_PP(16'h197D9,4);
TASK_PP(16'h197DA,4);
TASK_PP(16'h197DB,4);
TASK_PP(16'h197DC,4);
TASK_PP(16'h197DD,4);
TASK_PP(16'h197DE,4);
TASK_PP(16'h197DF,4);
TASK_PP(16'h197E0,4);
TASK_PP(16'h197E1,4);
TASK_PP(16'h197E2,4);
TASK_PP(16'h197E3,4);
TASK_PP(16'h197E4,4);
TASK_PP(16'h197E5,4);
TASK_PP(16'h197E6,4);
TASK_PP(16'h197E7,4);
TASK_PP(16'h197E8,4);
TASK_PP(16'h197E9,4);
TASK_PP(16'h197EA,4);
TASK_PP(16'h197EB,4);
TASK_PP(16'h197EC,4);
TASK_PP(16'h197ED,4);
TASK_PP(16'h197EE,4);
TASK_PP(16'h197EF,4);
TASK_PP(16'h197F0,4);
TASK_PP(16'h197F1,4);
TASK_PP(16'h197F2,4);
TASK_PP(16'h197F3,4);
TASK_PP(16'h197F4,4);
TASK_PP(16'h197F5,4);
TASK_PP(16'h197F6,4);
TASK_PP(16'h197F7,4);
TASK_PP(16'h197F8,4);
TASK_PP(16'h197F9,4);
TASK_PP(16'h197FA,4);
TASK_PP(16'h197FB,4);
TASK_PP(16'h197FC,4);
TASK_PP(16'h197FD,4);
TASK_PP(16'h197FE,4);
TASK_PP(16'h197FF,4);
TASK_PP(16'h19800,4);
TASK_PP(16'h19801,4);
TASK_PP(16'h19802,4);
TASK_PP(16'h19803,4);
TASK_PP(16'h19804,4);
TASK_PP(16'h19805,4);
TASK_PP(16'h19806,4);
TASK_PP(16'h19807,4);
TASK_PP(16'h19808,4);
TASK_PP(16'h19809,4);
TASK_PP(16'h1980A,4);
TASK_PP(16'h1980B,4);
TASK_PP(16'h1980C,4);
TASK_PP(16'h1980D,4);
TASK_PP(16'h1980E,4);
TASK_PP(16'h1980F,4);
TASK_PP(16'h19810,4);
TASK_PP(16'h19811,4);
TASK_PP(16'h19812,4);
TASK_PP(16'h19813,4);
TASK_PP(16'h19814,4);
TASK_PP(16'h19815,4);
TASK_PP(16'h19816,4);
TASK_PP(16'h19817,4);
TASK_PP(16'h19818,4);
TASK_PP(16'h19819,4);
TASK_PP(16'h1981A,4);
TASK_PP(16'h1981B,4);
TASK_PP(16'h1981C,4);
TASK_PP(16'h1981D,4);
TASK_PP(16'h1981E,4);
TASK_PP(16'h1981F,4);
TASK_PP(16'h19820,4);
TASK_PP(16'h19821,4);
TASK_PP(16'h19822,4);
TASK_PP(16'h19823,4);
TASK_PP(16'h19824,4);
TASK_PP(16'h19825,4);
TASK_PP(16'h19826,4);
TASK_PP(16'h19827,4);
TASK_PP(16'h19828,4);
TASK_PP(16'h19829,4);
TASK_PP(16'h1982A,4);
TASK_PP(16'h1982B,4);
TASK_PP(16'h1982C,4);
TASK_PP(16'h1982D,4);
TASK_PP(16'h1982E,4);
TASK_PP(16'h1982F,4);
TASK_PP(16'h19830,4);
TASK_PP(16'h19831,4);
TASK_PP(16'h19832,4);
TASK_PP(16'h19833,4);
TASK_PP(16'h19834,4);
TASK_PP(16'h19835,4);
TASK_PP(16'h19836,4);
TASK_PP(16'h19837,4);
TASK_PP(16'h19838,4);
TASK_PP(16'h19839,4);
TASK_PP(16'h1983A,4);
TASK_PP(16'h1983B,4);
TASK_PP(16'h1983C,4);
TASK_PP(16'h1983D,4);
TASK_PP(16'h1983E,4);
TASK_PP(16'h1983F,4);
TASK_PP(16'h19840,4);
TASK_PP(16'h19841,4);
TASK_PP(16'h19842,4);
TASK_PP(16'h19843,4);
TASK_PP(16'h19844,4);
TASK_PP(16'h19845,4);
TASK_PP(16'h19846,4);
TASK_PP(16'h19847,4);
TASK_PP(16'h19848,4);
TASK_PP(16'h19849,4);
TASK_PP(16'h1984A,4);
TASK_PP(16'h1984B,4);
TASK_PP(16'h1984C,4);
TASK_PP(16'h1984D,4);
TASK_PP(16'h1984E,4);
TASK_PP(16'h1984F,4);
TASK_PP(16'h19850,4);
TASK_PP(16'h19851,4);
TASK_PP(16'h19852,4);
TASK_PP(16'h19853,4);
TASK_PP(16'h19854,4);
TASK_PP(16'h19855,4);
TASK_PP(16'h19856,4);
TASK_PP(16'h19857,4);
TASK_PP(16'h19858,4);
TASK_PP(16'h19859,4);
TASK_PP(16'h1985A,4);
TASK_PP(16'h1985B,4);
TASK_PP(16'h1985C,4);
TASK_PP(16'h1985D,4);
TASK_PP(16'h1985E,4);
TASK_PP(16'h1985F,4);
TASK_PP(16'h19860,4);
TASK_PP(16'h19861,4);
TASK_PP(16'h19862,4);
TASK_PP(16'h19863,4);
TASK_PP(16'h19864,4);
TASK_PP(16'h19865,4);
TASK_PP(16'h19866,4);
TASK_PP(16'h19867,4);
TASK_PP(16'h19868,4);
TASK_PP(16'h19869,4);
TASK_PP(16'h1986A,4);
TASK_PP(16'h1986B,4);
TASK_PP(16'h1986C,4);
TASK_PP(16'h1986D,4);
TASK_PP(16'h1986E,4);
TASK_PP(16'h1986F,4);
TASK_PP(16'h19870,4);
TASK_PP(16'h19871,4);
TASK_PP(16'h19872,4);
TASK_PP(16'h19873,4);
TASK_PP(16'h19874,4);
TASK_PP(16'h19875,4);
TASK_PP(16'h19876,4);
TASK_PP(16'h19877,4);
TASK_PP(16'h19878,4);
TASK_PP(16'h19879,4);
TASK_PP(16'h1987A,4);
TASK_PP(16'h1987B,4);
TASK_PP(16'h1987C,4);
TASK_PP(16'h1987D,4);
TASK_PP(16'h1987E,4);
TASK_PP(16'h1987F,4);
TASK_PP(16'h19880,4);
TASK_PP(16'h19881,4);
TASK_PP(16'h19882,4);
TASK_PP(16'h19883,4);
TASK_PP(16'h19884,4);
TASK_PP(16'h19885,4);
TASK_PP(16'h19886,4);
TASK_PP(16'h19887,4);
TASK_PP(16'h19888,4);
TASK_PP(16'h19889,4);
TASK_PP(16'h1988A,4);
TASK_PP(16'h1988B,4);
TASK_PP(16'h1988C,4);
TASK_PP(16'h1988D,4);
TASK_PP(16'h1988E,4);
TASK_PP(16'h1988F,4);
TASK_PP(16'h19890,4);
TASK_PP(16'h19891,4);
TASK_PP(16'h19892,4);
TASK_PP(16'h19893,4);
TASK_PP(16'h19894,4);
TASK_PP(16'h19895,4);
TASK_PP(16'h19896,4);
TASK_PP(16'h19897,4);
TASK_PP(16'h19898,4);
TASK_PP(16'h19899,4);
TASK_PP(16'h1989A,4);
TASK_PP(16'h1989B,4);
TASK_PP(16'h1989C,4);
TASK_PP(16'h1989D,4);
TASK_PP(16'h1989E,4);
TASK_PP(16'h1989F,4);
TASK_PP(16'h198A0,4);
TASK_PP(16'h198A1,4);
TASK_PP(16'h198A2,4);
TASK_PP(16'h198A3,4);
TASK_PP(16'h198A4,4);
TASK_PP(16'h198A5,4);
TASK_PP(16'h198A6,4);
TASK_PP(16'h198A7,4);
TASK_PP(16'h198A8,4);
TASK_PP(16'h198A9,4);
TASK_PP(16'h198AA,4);
TASK_PP(16'h198AB,4);
TASK_PP(16'h198AC,4);
TASK_PP(16'h198AD,4);
TASK_PP(16'h198AE,4);
TASK_PP(16'h198AF,4);
TASK_PP(16'h198B0,4);
TASK_PP(16'h198B1,4);
TASK_PP(16'h198B2,4);
TASK_PP(16'h198B3,4);
TASK_PP(16'h198B4,4);
TASK_PP(16'h198B5,4);
TASK_PP(16'h198B6,4);
TASK_PP(16'h198B7,4);
TASK_PP(16'h198B8,4);
TASK_PP(16'h198B9,4);
TASK_PP(16'h198BA,4);
TASK_PP(16'h198BB,4);
TASK_PP(16'h198BC,4);
TASK_PP(16'h198BD,4);
TASK_PP(16'h198BE,4);
TASK_PP(16'h198BF,4);
TASK_PP(16'h198C0,4);
TASK_PP(16'h198C1,4);
TASK_PP(16'h198C2,4);
TASK_PP(16'h198C3,4);
TASK_PP(16'h198C4,4);
TASK_PP(16'h198C5,4);
TASK_PP(16'h198C6,4);
TASK_PP(16'h198C7,4);
TASK_PP(16'h198C8,4);
TASK_PP(16'h198C9,4);
TASK_PP(16'h198CA,4);
TASK_PP(16'h198CB,4);
TASK_PP(16'h198CC,4);
TASK_PP(16'h198CD,4);
TASK_PP(16'h198CE,4);
TASK_PP(16'h198CF,4);
TASK_PP(16'h198D0,4);
TASK_PP(16'h198D1,4);
TASK_PP(16'h198D2,4);
TASK_PP(16'h198D3,4);
TASK_PP(16'h198D4,4);
TASK_PP(16'h198D5,4);
TASK_PP(16'h198D6,4);
TASK_PP(16'h198D7,4);
TASK_PP(16'h198D8,4);
TASK_PP(16'h198D9,4);
TASK_PP(16'h198DA,4);
TASK_PP(16'h198DB,4);
TASK_PP(16'h198DC,4);
TASK_PP(16'h198DD,4);
TASK_PP(16'h198DE,4);
TASK_PP(16'h198DF,4);
TASK_PP(16'h198E0,4);
TASK_PP(16'h198E1,4);
TASK_PP(16'h198E2,4);
TASK_PP(16'h198E3,4);
TASK_PP(16'h198E4,4);
TASK_PP(16'h198E5,4);
TASK_PP(16'h198E6,4);
TASK_PP(16'h198E7,4);
TASK_PP(16'h198E8,4);
TASK_PP(16'h198E9,4);
TASK_PP(16'h198EA,4);
TASK_PP(16'h198EB,4);
TASK_PP(16'h198EC,4);
TASK_PP(16'h198ED,4);
TASK_PP(16'h198EE,4);
TASK_PP(16'h198EF,4);
TASK_PP(16'h198F0,4);
TASK_PP(16'h198F1,4);
TASK_PP(16'h198F2,4);
TASK_PP(16'h198F3,4);
TASK_PP(16'h198F4,4);
TASK_PP(16'h198F5,4);
TASK_PP(16'h198F6,4);
TASK_PP(16'h198F7,4);
TASK_PP(16'h198F8,4);
TASK_PP(16'h198F9,4);
TASK_PP(16'h198FA,4);
TASK_PP(16'h198FB,4);
TASK_PP(16'h198FC,4);
TASK_PP(16'h198FD,4);
TASK_PP(16'h198FE,4);
TASK_PP(16'h198FF,4);
TASK_PP(16'h19900,4);
TASK_PP(16'h19901,4);
TASK_PP(16'h19902,4);
TASK_PP(16'h19903,4);
TASK_PP(16'h19904,4);
TASK_PP(16'h19905,4);
TASK_PP(16'h19906,4);
TASK_PP(16'h19907,4);
TASK_PP(16'h19908,4);
TASK_PP(16'h19909,4);
TASK_PP(16'h1990A,4);
TASK_PP(16'h1990B,4);
TASK_PP(16'h1990C,4);
TASK_PP(16'h1990D,4);
TASK_PP(16'h1990E,4);
TASK_PP(16'h1990F,4);
TASK_PP(16'h19910,4);
TASK_PP(16'h19911,4);
TASK_PP(16'h19912,4);
TASK_PP(16'h19913,4);
TASK_PP(16'h19914,4);
TASK_PP(16'h19915,4);
TASK_PP(16'h19916,4);
TASK_PP(16'h19917,4);
TASK_PP(16'h19918,4);
TASK_PP(16'h19919,4);
TASK_PP(16'h1991A,4);
TASK_PP(16'h1991B,4);
TASK_PP(16'h1991C,4);
TASK_PP(16'h1991D,4);
TASK_PP(16'h1991E,4);
TASK_PP(16'h1991F,4);
TASK_PP(16'h19920,4);
TASK_PP(16'h19921,4);
TASK_PP(16'h19922,4);
TASK_PP(16'h19923,4);
TASK_PP(16'h19924,4);
TASK_PP(16'h19925,4);
TASK_PP(16'h19926,4);
TASK_PP(16'h19927,4);
TASK_PP(16'h19928,4);
TASK_PP(16'h19929,4);
TASK_PP(16'h1992A,4);
TASK_PP(16'h1992B,4);
TASK_PP(16'h1992C,4);
TASK_PP(16'h1992D,4);
TASK_PP(16'h1992E,4);
TASK_PP(16'h1992F,4);
TASK_PP(16'h19930,4);
TASK_PP(16'h19931,4);
TASK_PP(16'h19932,4);
TASK_PP(16'h19933,4);
TASK_PP(16'h19934,4);
TASK_PP(16'h19935,4);
TASK_PP(16'h19936,4);
TASK_PP(16'h19937,4);
TASK_PP(16'h19938,4);
TASK_PP(16'h19939,4);
TASK_PP(16'h1993A,4);
TASK_PP(16'h1993B,4);
TASK_PP(16'h1993C,4);
TASK_PP(16'h1993D,4);
TASK_PP(16'h1993E,4);
TASK_PP(16'h1993F,4);
TASK_PP(16'h19940,4);
TASK_PP(16'h19941,4);
TASK_PP(16'h19942,4);
TASK_PP(16'h19943,4);
TASK_PP(16'h19944,4);
TASK_PP(16'h19945,4);
TASK_PP(16'h19946,4);
TASK_PP(16'h19947,4);
TASK_PP(16'h19948,4);
TASK_PP(16'h19949,4);
TASK_PP(16'h1994A,4);
TASK_PP(16'h1994B,4);
TASK_PP(16'h1994C,4);
TASK_PP(16'h1994D,4);
TASK_PP(16'h1994E,4);
TASK_PP(16'h1994F,4);
TASK_PP(16'h19950,4);
TASK_PP(16'h19951,4);
TASK_PP(16'h19952,4);
TASK_PP(16'h19953,4);
TASK_PP(16'h19954,4);
TASK_PP(16'h19955,4);
TASK_PP(16'h19956,4);
TASK_PP(16'h19957,4);
TASK_PP(16'h19958,4);
TASK_PP(16'h19959,4);
TASK_PP(16'h1995A,4);
TASK_PP(16'h1995B,4);
TASK_PP(16'h1995C,4);
TASK_PP(16'h1995D,4);
TASK_PP(16'h1995E,4);
TASK_PP(16'h1995F,4);
TASK_PP(16'h19960,4);
TASK_PP(16'h19961,4);
TASK_PP(16'h19962,4);
TASK_PP(16'h19963,4);
TASK_PP(16'h19964,4);
TASK_PP(16'h19965,4);
TASK_PP(16'h19966,4);
TASK_PP(16'h19967,4);
TASK_PP(16'h19968,4);
TASK_PP(16'h19969,4);
TASK_PP(16'h1996A,4);
TASK_PP(16'h1996B,4);
TASK_PP(16'h1996C,4);
TASK_PP(16'h1996D,4);
TASK_PP(16'h1996E,4);
TASK_PP(16'h1996F,4);
TASK_PP(16'h19970,4);
TASK_PP(16'h19971,4);
TASK_PP(16'h19972,4);
TASK_PP(16'h19973,4);
TASK_PP(16'h19974,4);
TASK_PP(16'h19975,4);
TASK_PP(16'h19976,4);
TASK_PP(16'h19977,4);
TASK_PP(16'h19978,4);
TASK_PP(16'h19979,4);
TASK_PP(16'h1997A,4);
TASK_PP(16'h1997B,4);
TASK_PP(16'h1997C,4);
TASK_PP(16'h1997D,4);
TASK_PP(16'h1997E,4);
TASK_PP(16'h1997F,4);
TASK_PP(16'h19980,4);
TASK_PP(16'h19981,4);
TASK_PP(16'h19982,4);
TASK_PP(16'h19983,4);
TASK_PP(16'h19984,4);
TASK_PP(16'h19985,4);
TASK_PP(16'h19986,4);
TASK_PP(16'h19987,4);
TASK_PP(16'h19988,4);
TASK_PP(16'h19989,4);
TASK_PP(16'h1998A,4);
TASK_PP(16'h1998B,4);
TASK_PP(16'h1998C,4);
TASK_PP(16'h1998D,4);
TASK_PP(16'h1998E,4);
TASK_PP(16'h1998F,4);
TASK_PP(16'h19990,4);
TASK_PP(16'h19991,4);
TASK_PP(16'h19992,4);
TASK_PP(16'h19993,4);
TASK_PP(16'h19994,4);
TASK_PP(16'h19995,4);
TASK_PP(16'h19996,4);
TASK_PP(16'h19997,4);
TASK_PP(16'h19998,4);
TASK_PP(16'h19999,4);
TASK_PP(16'h1999A,4);
TASK_PP(16'h1999B,4);
TASK_PP(16'h1999C,4);
TASK_PP(16'h1999D,4);
TASK_PP(16'h1999E,4);
TASK_PP(16'h1999F,4);
TASK_PP(16'h199A0,4);
TASK_PP(16'h199A1,4);
TASK_PP(16'h199A2,4);
TASK_PP(16'h199A3,4);
TASK_PP(16'h199A4,4);
TASK_PP(16'h199A5,4);
TASK_PP(16'h199A6,4);
TASK_PP(16'h199A7,4);
TASK_PP(16'h199A8,4);
TASK_PP(16'h199A9,4);
TASK_PP(16'h199AA,4);
TASK_PP(16'h199AB,4);
TASK_PP(16'h199AC,4);
TASK_PP(16'h199AD,4);
TASK_PP(16'h199AE,4);
TASK_PP(16'h199AF,4);
TASK_PP(16'h199B0,4);
TASK_PP(16'h199B1,4);
TASK_PP(16'h199B2,4);
TASK_PP(16'h199B3,4);
TASK_PP(16'h199B4,4);
TASK_PP(16'h199B5,4);
TASK_PP(16'h199B6,4);
TASK_PP(16'h199B7,4);
TASK_PP(16'h199B8,4);
TASK_PP(16'h199B9,4);
TASK_PP(16'h199BA,4);
TASK_PP(16'h199BB,4);
TASK_PP(16'h199BC,4);
TASK_PP(16'h199BD,4);
TASK_PP(16'h199BE,4);
TASK_PP(16'h199BF,4);
TASK_PP(16'h199C0,4);
TASK_PP(16'h199C1,4);
TASK_PP(16'h199C2,4);
TASK_PP(16'h199C3,4);
TASK_PP(16'h199C4,4);
TASK_PP(16'h199C5,4);
TASK_PP(16'h199C6,4);
TASK_PP(16'h199C7,4);
TASK_PP(16'h199C8,4);
TASK_PP(16'h199C9,4);
TASK_PP(16'h199CA,4);
TASK_PP(16'h199CB,4);
TASK_PP(16'h199CC,4);
TASK_PP(16'h199CD,4);
TASK_PP(16'h199CE,4);
TASK_PP(16'h199CF,4);
TASK_PP(16'h199D0,4);
TASK_PP(16'h199D1,4);
TASK_PP(16'h199D2,4);
TASK_PP(16'h199D3,4);
TASK_PP(16'h199D4,4);
TASK_PP(16'h199D5,4);
TASK_PP(16'h199D6,4);
TASK_PP(16'h199D7,4);
TASK_PP(16'h199D8,4);
TASK_PP(16'h199D9,4);
TASK_PP(16'h199DA,4);
TASK_PP(16'h199DB,4);
TASK_PP(16'h199DC,4);
TASK_PP(16'h199DD,4);
TASK_PP(16'h199DE,4);
TASK_PP(16'h199DF,4);
TASK_PP(16'h199E0,4);
TASK_PP(16'h199E1,4);
TASK_PP(16'h199E2,4);
TASK_PP(16'h199E3,4);
TASK_PP(16'h199E4,4);
TASK_PP(16'h199E5,4);
TASK_PP(16'h199E6,4);
TASK_PP(16'h199E7,4);
TASK_PP(16'h199E8,4);
TASK_PP(16'h199E9,4);
TASK_PP(16'h199EA,4);
TASK_PP(16'h199EB,4);
TASK_PP(16'h199EC,4);
TASK_PP(16'h199ED,4);
TASK_PP(16'h199EE,4);
TASK_PP(16'h199EF,4);
TASK_PP(16'h199F0,4);
TASK_PP(16'h199F1,4);
TASK_PP(16'h199F2,4);
TASK_PP(16'h199F3,4);
TASK_PP(16'h199F4,4);
TASK_PP(16'h199F5,4);
TASK_PP(16'h199F6,4);
TASK_PP(16'h199F7,4);
TASK_PP(16'h199F8,4);
TASK_PP(16'h199F9,4);
TASK_PP(16'h199FA,4);
TASK_PP(16'h199FB,4);
TASK_PP(16'h199FC,4);
TASK_PP(16'h199FD,4);
TASK_PP(16'h199FE,4);
TASK_PP(16'h199FF,4);
TASK_PP(16'h19A00,4);
TASK_PP(16'h19A01,4);
TASK_PP(16'h19A02,4);
TASK_PP(16'h19A03,4);
TASK_PP(16'h19A04,4);
TASK_PP(16'h19A05,4);
TASK_PP(16'h19A06,4);
TASK_PP(16'h19A07,4);
TASK_PP(16'h19A08,4);
TASK_PP(16'h19A09,4);
TASK_PP(16'h19A0A,4);
TASK_PP(16'h19A0B,4);
TASK_PP(16'h19A0C,4);
TASK_PP(16'h19A0D,4);
TASK_PP(16'h19A0E,4);
TASK_PP(16'h19A0F,4);
TASK_PP(16'h19A10,4);
TASK_PP(16'h19A11,4);
TASK_PP(16'h19A12,4);
TASK_PP(16'h19A13,4);
TASK_PP(16'h19A14,4);
TASK_PP(16'h19A15,4);
TASK_PP(16'h19A16,4);
TASK_PP(16'h19A17,4);
TASK_PP(16'h19A18,4);
TASK_PP(16'h19A19,4);
TASK_PP(16'h19A1A,4);
TASK_PP(16'h19A1B,4);
TASK_PP(16'h19A1C,4);
TASK_PP(16'h19A1D,4);
TASK_PP(16'h19A1E,4);
TASK_PP(16'h19A1F,4);
TASK_PP(16'h19A20,4);
TASK_PP(16'h19A21,4);
TASK_PP(16'h19A22,4);
TASK_PP(16'h19A23,4);
TASK_PP(16'h19A24,4);
TASK_PP(16'h19A25,4);
TASK_PP(16'h19A26,4);
TASK_PP(16'h19A27,4);
TASK_PP(16'h19A28,4);
TASK_PP(16'h19A29,4);
TASK_PP(16'h19A2A,4);
TASK_PP(16'h19A2B,4);
TASK_PP(16'h19A2C,4);
TASK_PP(16'h19A2D,4);
TASK_PP(16'h19A2E,4);
TASK_PP(16'h19A2F,4);
TASK_PP(16'h19A30,4);
TASK_PP(16'h19A31,4);
TASK_PP(16'h19A32,4);
TASK_PP(16'h19A33,4);
TASK_PP(16'h19A34,4);
TASK_PP(16'h19A35,4);
TASK_PP(16'h19A36,4);
TASK_PP(16'h19A37,4);
TASK_PP(16'h19A38,4);
TASK_PP(16'h19A39,4);
TASK_PP(16'h19A3A,4);
TASK_PP(16'h19A3B,4);
TASK_PP(16'h19A3C,4);
TASK_PP(16'h19A3D,4);
TASK_PP(16'h19A3E,4);
TASK_PP(16'h19A3F,4);
TASK_PP(16'h19A40,4);
TASK_PP(16'h19A41,4);
TASK_PP(16'h19A42,4);
TASK_PP(16'h19A43,4);
TASK_PP(16'h19A44,4);
TASK_PP(16'h19A45,4);
TASK_PP(16'h19A46,4);
TASK_PP(16'h19A47,4);
TASK_PP(16'h19A48,4);
TASK_PP(16'h19A49,4);
TASK_PP(16'h19A4A,4);
TASK_PP(16'h19A4B,4);
TASK_PP(16'h19A4C,4);
TASK_PP(16'h19A4D,4);
TASK_PP(16'h19A4E,4);
TASK_PP(16'h19A4F,4);
TASK_PP(16'h19A50,4);
TASK_PP(16'h19A51,4);
TASK_PP(16'h19A52,4);
TASK_PP(16'h19A53,4);
TASK_PP(16'h19A54,4);
TASK_PP(16'h19A55,4);
TASK_PP(16'h19A56,4);
TASK_PP(16'h19A57,4);
TASK_PP(16'h19A58,4);
TASK_PP(16'h19A59,4);
TASK_PP(16'h19A5A,4);
TASK_PP(16'h19A5B,4);
TASK_PP(16'h19A5C,4);
TASK_PP(16'h19A5D,4);
TASK_PP(16'h19A5E,4);
TASK_PP(16'h19A5F,4);
TASK_PP(16'h19A60,4);
TASK_PP(16'h19A61,4);
TASK_PP(16'h19A62,4);
TASK_PP(16'h19A63,4);
TASK_PP(16'h19A64,4);
TASK_PP(16'h19A65,4);
TASK_PP(16'h19A66,4);
TASK_PP(16'h19A67,4);
TASK_PP(16'h19A68,4);
TASK_PP(16'h19A69,4);
TASK_PP(16'h19A6A,4);
TASK_PP(16'h19A6B,4);
TASK_PP(16'h19A6C,4);
TASK_PP(16'h19A6D,4);
TASK_PP(16'h19A6E,4);
TASK_PP(16'h19A6F,4);
TASK_PP(16'h19A70,4);
TASK_PP(16'h19A71,4);
TASK_PP(16'h19A72,4);
TASK_PP(16'h19A73,4);
TASK_PP(16'h19A74,4);
TASK_PP(16'h19A75,4);
TASK_PP(16'h19A76,4);
TASK_PP(16'h19A77,4);
TASK_PP(16'h19A78,4);
TASK_PP(16'h19A79,4);
TASK_PP(16'h19A7A,4);
TASK_PP(16'h19A7B,4);
TASK_PP(16'h19A7C,4);
TASK_PP(16'h19A7D,4);
TASK_PP(16'h19A7E,4);
TASK_PP(16'h19A7F,4);
TASK_PP(16'h19A80,4);
TASK_PP(16'h19A81,4);
TASK_PP(16'h19A82,4);
TASK_PP(16'h19A83,4);
TASK_PP(16'h19A84,4);
TASK_PP(16'h19A85,4);
TASK_PP(16'h19A86,4);
TASK_PP(16'h19A87,4);
TASK_PP(16'h19A88,4);
TASK_PP(16'h19A89,4);
TASK_PP(16'h19A8A,4);
TASK_PP(16'h19A8B,4);
TASK_PP(16'h19A8C,4);
TASK_PP(16'h19A8D,4);
TASK_PP(16'h19A8E,4);
TASK_PP(16'h19A8F,4);
TASK_PP(16'h19A90,4);
TASK_PP(16'h19A91,4);
TASK_PP(16'h19A92,4);
TASK_PP(16'h19A93,4);
TASK_PP(16'h19A94,4);
TASK_PP(16'h19A95,4);
TASK_PP(16'h19A96,4);
TASK_PP(16'h19A97,4);
TASK_PP(16'h19A98,4);
TASK_PP(16'h19A99,4);
TASK_PP(16'h19A9A,4);
TASK_PP(16'h19A9B,4);
TASK_PP(16'h19A9C,4);
TASK_PP(16'h19A9D,4);
TASK_PP(16'h19A9E,4);
TASK_PP(16'h19A9F,4);
TASK_PP(16'h19AA0,4);
TASK_PP(16'h19AA1,4);
TASK_PP(16'h19AA2,4);
TASK_PP(16'h19AA3,4);
TASK_PP(16'h19AA4,4);
TASK_PP(16'h19AA5,4);
TASK_PP(16'h19AA6,4);
TASK_PP(16'h19AA7,4);
TASK_PP(16'h19AA8,4);
TASK_PP(16'h19AA9,4);
TASK_PP(16'h19AAA,4);
TASK_PP(16'h19AAB,4);
TASK_PP(16'h19AAC,4);
TASK_PP(16'h19AAD,4);
TASK_PP(16'h19AAE,4);
TASK_PP(16'h19AAF,4);
TASK_PP(16'h19AB0,4);
TASK_PP(16'h19AB1,4);
TASK_PP(16'h19AB2,4);
TASK_PP(16'h19AB3,4);
TASK_PP(16'h19AB4,4);
TASK_PP(16'h19AB5,4);
TASK_PP(16'h19AB6,4);
TASK_PP(16'h19AB7,4);
TASK_PP(16'h19AB8,4);
TASK_PP(16'h19AB9,4);
TASK_PP(16'h19ABA,4);
TASK_PP(16'h19ABB,4);
TASK_PP(16'h19ABC,4);
TASK_PP(16'h19ABD,4);
TASK_PP(16'h19ABE,4);
TASK_PP(16'h19ABF,4);
TASK_PP(16'h19AC0,4);
TASK_PP(16'h19AC1,4);
TASK_PP(16'h19AC2,4);
TASK_PP(16'h19AC3,4);
TASK_PP(16'h19AC4,4);
TASK_PP(16'h19AC5,4);
TASK_PP(16'h19AC6,4);
TASK_PP(16'h19AC7,4);
TASK_PP(16'h19AC8,4);
TASK_PP(16'h19AC9,4);
TASK_PP(16'h19ACA,4);
TASK_PP(16'h19ACB,4);
TASK_PP(16'h19ACC,4);
TASK_PP(16'h19ACD,4);
TASK_PP(16'h19ACE,4);
TASK_PP(16'h19ACF,4);
TASK_PP(16'h19AD0,4);
TASK_PP(16'h19AD1,4);
TASK_PP(16'h19AD2,4);
TASK_PP(16'h19AD3,4);
TASK_PP(16'h19AD4,4);
TASK_PP(16'h19AD5,4);
TASK_PP(16'h19AD6,4);
TASK_PP(16'h19AD7,4);
TASK_PP(16'h19AD8,4);
TASK_PP(16'h19AD9,4);
TASK_PP(16'h19ADA,4);
TASK_PP(16'h19ADB,4);
TASK_PP(16'h19ADC,4);
TASK_PP(16'h19ADD,4);
TASK_PP(16'h19ADE,4);
TASK_PP(16'h19ADF,4);
TASK_PP(16'h19AE0,4);
TASK_PP(16'h19AE1,4);
TASK_PP(16'h19AE2,4);
TASK_PP(16'h19AE3,4);
TASK_PP(16'h19AE4,4);
TASK_PP(16'h19AE5,4);
TASK_PP(16'h19AE6,4);
TASK_PP(16'h19AE7,4);
TASK_PP(16'h19AE8,4);
TASK_PP(16'h19AE9,4);
TASK_PP(16'h19AEA,4);
TASK_PP(16'h19AEB,4);
TASK_PP(16'h19AEC,4);
TASK_PP(16'h19AED,4);
TASK_PP(16'h19AEE,4);
TASK_PP(16'h19AEF,4);
TASK_PP(16'h19AF0,4);
TASK_PP(16'h19AF1,4);
TASK_PP(16'h19AF2,4);
TASK_PP(16'h19AF3,4);
TASK_PP(16'h19AF4,4);
TASK_PP(16'h19AF5,4);
TASK_PP(16'h19AF6,4);
TASK_PP(16'h19AF7,4);
TASK_PP(16'h19AF8,4);
TASK_PP(16'h19AF9,4);
TASK_PP(16'h19AFA,4);
TASK_PP(16'h19AFB,4);
TASK_PP(16'h19AFC,4);
TASK_PP(16'h19AFD,4);
TASK_PP(16'h19AFE,4);
TASK_PP(16'h19AFF,4);
TASK_PP(16'h19B00,4);
TASK_PP(16'h19B01,4);
TASK_PP(16'h19B02,4);
TASK_PP(16'h19B03,4);
TASK_PP(16'h19B04,4);
TASK_PP(16'h19B05,4);
TASK_PP(16'h19B06,4);
TASK_PP(16'h19B07,4);
TASK_PP(16'h19B08,4);
TASK_PP(16'h19B09,4);
TASK_PP(16'h19B0A,4);
TASK_PP(16'h19B0B,4);
TASK_PP(16'h19B0C,4);
TASK_PP(16'h19B0D,4);
TASK_PP(16'h19B0E,4);
TASK_PP(16'h19B0F,4);
TASK_PP(16'h19B10,4);
TASK_PP(16'h19B11,4);
TASK_PP(16'h19B12,4);
TASK_PP(16'h19B13,4);
TASK_PP(16'h19B14,4);
TASK_PP(16'h19B15,4);
TASK_PP(16'h19B16,4);
TASK_PP(16'h19B17,4);
TASK_PP(16'h19B18,4);
TASK_PP(16'h19B19,4);
TASK_PP(16'h19B1A,4);
TASK_PP(16'h19B1B,4);
TASK_PP(16'h19B1C,4);
TASK_PP(16'h19B1D,4);
TASK_PP(16'h19B1E,4);
TASK_PP(16'h19B1F,4);
TASK_PP(16'h19B20,4);
TASK_PP(16'h19B21,4);
TASK_PP(16'h19B22,4);
TASK_PP(16'h19B23,4);
TASK_PP(16'h19B24,4);
TASK_PP(16'h19B25,4);
TASK_PP(16'h19B26,4);
TASK_PP(16'h19B27,4);
TASK_PP(16'h19B28,4);
TASK_PP(16'h19B29,4);
TASK_PP(16'h19B2A,4);
TASK_PP(16'h19B2B,4);
TASK_PP(16'h19B2C,4);
TASK_PP(16'h19B2D,4);
TASK_PP(16'h19B2E,4);
TASK_PP(16'h19B2F,4);
TASK_PP(16'h19B30,4);
TASK_PP(16'h19B31,4);
TASK_PP(16'h19B32,4);
TASK_PP(16'h19B33,4);
TASK_PP(16'h19B34,4);
TASK_PP(16'h19B35,4);
TASK_PP(16'h19B36,4);
TASK_PP(16'h19B37,4);
TASK_PP(16'h19B38,4);
TASK_PP(16'h19B39,4);
TASK_PP(16'h19B3A,4);
TASK_PP(16'h19B3B,4);
TASK_PP(16'h19B3C,4);
TASK_PP(16'h19B3D,4);
TASK_PP(16'h19B3E,4);
TASK_PP(16'h19B3F,4);
TASK_PP(16'h19B40,4);
TASK_PP(16'h19B41,4);
TASK_PP(16'h19B42,4);
TASK_PP(16'h19B43,4);
TASK_PP(16'h19B44,4);
TASK_PP(16'h19B45,4);
TASK_PP(16'h19B46,4);
TASK_PP(16'h19B47,4);
TASK_PP(16'h19B48,4);
TASK_PP(16'h19B49,4);
TASK_PP(16'h19B4A,4);
TASK_PP(16'h19B4B,4);
TASK_PP(16'h19B4C,4);
TASK_PP(16'h19B4D,4);
TASK_PP(16'h19B4E,4);
TASK_PP(16'h19B4F,4);
TASK_PP(16'h19B50,4);
TASK_PP(16'h19B51,4);
TASK_PP(16'h19B52,4);
TASK_PP(16'h19B53,4);
TASK_PP(16'h19B54,4);
TASK_PP(16'h19B55,4);
TASK_PP(16'h19B56,4);
TASK_PP(16'h19B57,4);
TASK_PP(16'h19B58,4);
TASK_PP(16'h19B59,4);
TASK_PP(16'h19B5A,4);
TASK_PP(16'h19B5B,4);
TASK_PP(16'h19B5C,4);
TASK_PP(16'h19B5D,4);
TASK_PP(16'h19B5E,4);
TASK_PP(16'h19B5F,4);
TASK_PP(16'h19B60,4);
TASK_PP(16'h19B61,4);
TASK_PP(16'h19B62,4);
TASK_PP(16'h19B63,4);
TASK_PP(16'h19B64,4);
TASK_PP(16'h19B65,4);
TASK_PP(16'h19B66,4);
TASK_PP(16'h19B67,4);
TASK_PP(16'h19B68,4);
TASK_PP(16'h19B69,4);
TASK_PP(16'h19B6A,4);
TASK_PP(16'h19B6B,4);
TASK_PP(16'h19B6C,4);
TASK_PP(16'h19B6D,4);
TASK_PP(16'h19B6E,4);
TASK_PP(16'h19B6F,4);
TASK_PP(16'h19B70,4);
TASK_PP(16'h19B71,4);
TASK_PP(16'h19B72,4);
TASK_PP(16'h19B73,4);
TASK_PP(16'h19B74,4);
TASK_PP(16'h19B75,4);
TASK_PP(16'h19B76,4);
TASK_PP(16'h19B77,4);
TASK_PP(16'h19B78,4);
TASK_PP(16'h19B79,4);
TASK_PP(16'h19B7A,4);
TASK_PP(16'h19B7B,4);
TASK_PP(16'h19B7C,4);
TASK_PP(16'h19B7D,4);
TASK_PP(16'h19B7E,4);
TASK_PP(16'h19B7F,4);
TASK_PP(16'h19B80,4);
TASK_PP(16'h19B81,4);
TASK_PP(16'h19B82,4);
TASK_PP(16'h19B83,4);
TASK_PP(16'h19B84,4);
TASK_PP(16'h19B85,4);
TASK_PP(16'h19B86,4);
TASK_PP(16'h19B87,4);
TASK_PP(16'h19B88,4);
TASK_PP(16'h19B89,4);
TASK_PP(16'h19B8A,4);
TASK_PP(16'h19B8B,4);
TASK_PP(16'h19B8C,4);
TASK_PP(16'h19B8D,4);
TASK_PP(16'h19B8E,4);
TASK_PP(16'h19B8F,4);
TASK_PP(16'h19B90,4);
TASK_PP(16'h19B91,4);
TASK_PP(16'h19B92,4);
TASK_PP(16'h19B93,4);
TASK_PP(16'h19B94,4);
TASK_PP(16'h19B95,4);
TASK_PP(16'h19B96,4);
TASK_PP(16'h19B97,4);
TASK_PP(16'h19B98,4);
TASK_PP(16'h19B99,4);
TASK_PP(16'h19B9A,4);
TASK_PP(16'h19B9B,4);
TASK_PP(16'h19B9C,4);
TASK_PP(16'h19B9D,4);
TASK_PP(16'h19B9E,4);
TASK_PP(16'h19B9F,4);
TASK_PP(16'h19BA0,4);
TASK_PP(16'h19BA1,4);
TASK_PP(16'h19BA2,4);
TASK_PP(16'h19BA3,4);
TASK_PP(16'h19BA4,4);
TASK_PP(16'h19BA5,4);
TASK_PP(16'h19BA6,4);
TASK_PP(16'h19BA7,4);
TASK_PP(16'h19BA8,4);
TASK_PP(16'h19BA9,4);
TASK_PP(16'h19BAA,4);
TASK_PP(16'h19BAB,4);
TASK_PP(16'h19BAC,4);
TASK_PP(16'h19BAD,4);
TASK_PP(16'h19BAE,4);
TASK_PP(16'h19BAF,4);
TASK_PP(16'h19BB0,4);
TASK_PP(16'h19BB1,4);
TASK_PP(16'h19BB2,4);
TASK_PP(16'h19BB3,4);
TASK_PP(16'h19BB4,4);
TASK_PP(16'h19BB5,4);
TASK_PP(16'h19BB6,4);
TASK_PP(16'h19BB7,4);
TASK_PP(16'h19BB8,4);
TASK_PP(16'h19BB9,4);
TASK_PP(16'h19BBA,4);
TASK_PP(16'h19BBB,4);
TASK_PP(16'h19BBC,4);
TASK_PP(16'h19BBD,4);
TASK_PP(16'h19BBE,4);
TASK_PP(16'h19BBF,4);
TASK_PP(16'h19BC0,4);
TASK_PP(16'h19BC1,4);
TASK_PP(16'h19BC2,4);
TASK_PP(16'h19BC3,4);
TASK_PP(16'h19BC4,4);
TASK_PP(16'h19BC5,4);
TASK_PP(16'h19BC6,4);
TASK_PP(16'h19BC7,4);
TASK_PP(16'h19BC8,4);
TASK_PP(16'h19BC9,4);
TASK_PP(16'h19BCA,4);
TASK_PP(16'h19BCB,4);
TASK_PP(16'h19BCC,4);
TASK_PP(16'h19BCD,4);
TASK_PP(16'h19BCE,4);
TASK_PP(16'h19BCF,4);
TASK_PP(16'h19BD0,4);
TASK_PP(16'h19BD1,4);
TASK_PP(16'h19BD2,4);
TASK_PP(16'h19BD3,4);
TASK_PP(16'h19BD4,4);
TASK_PP(16'h19BD5,4);
TASK_PP(16'h19BD6,4);
TASK_PP(16'h19BD7,4);
TASK_PP(16'h19BD8,4);
TASK_PP(16'h19BD9,4);
TASK_PP(16'h19BDA,4);
TASK_PP(16'h19BDB,4);
TASK_PP(16'h19BDC,4);
TASK_PP(16'h19BDD,4);
TASK_PP(16'h19BDE,4);
TASK_PP(16'h19BDF,4);
TASK_PP(16'h19BE0,4);
TASK_PP(16'h19BE1,4);
TASK_PP(16'h19BE2,4);
TASK_PP(16'h19BE3,4);
TASK_PP(16'h19BE4,4);
TASK_PP(16'h19BE5,4);
TASK_PP(16'h19BE6,4);
TASK_PP(16'h19BE7,4);
TASK_PP(16'h19BE8,4);
TASK_PP(16'h19BE9,4);
TASK_PP(16'h19BEA,4);
TASK_PP(16'h19BEB,4);
TASK_PP(16'h19BEC,4);
TASK_PP(16'h19BED,4);
TASK_PP(16'h19BEE,4);
TASK_PP(16'h19BEF,4);
TASK_PP(16'h19BF0,4);
TASK_PP(16'h19BF1,4);
TASK_PP(16'h19BF2,4);
TASK_PP(16'h19BF3,4);
TASK_PP(16'h19BF4,4);
TASK_PP(16'h19BF5,4);
TASK_PP(16'h19BF6,4);
TASK_PP(16'h19BF7,4);
TASK_PP(16'h19BF8,4);
TASK_PP(16'h19BF9,4);
TASK_PP(16'h19BFA,4);
TASK_PP(16'h19BFB,4);
TASK_PP(16'h19BFC,4);
TASK_PP(16'h19BFD,4);
TASK_PP(16'h19BFE,4);
TASK_PP(16'h19BFF,4);
TASK_PP(16'h19C00,4);
TASK_PP(16'h19C01,4);
TASK_PP(16'h19C02,4);
TASK_PP(16'h19C03,4);
TASK_PP(16'h19C04,4);
TASK_PP(16'h19C05,4);
TASK_PP(16'h19C06,4);
TASK_PP(16'h19C07,4);
TASK_PP(16'h19C08,4);
TASK_PP(16'h19C09,4);
TASK_PP(16'h19C0A,4);
TASK_PP(16'h19C0B,4);
TASK_PP(16'h19C0C,4);
TASK_PP(16'h19C0D,4);
TASK_PP(16'h19C0E,4);
TASK_PP(16'h19C0F,4);
TASK_PP(16'h19C10,4);
TASK_PP(16'h19C11,4);
TASK_PP(16'h19C12,4);
TASK_PP(16'h19C13,4);
TASK_PP(16'h19C14,4);
TASK_PP(16'h19C15,4);
TASK_PP(16'h19C16,4);
TASK_PP(16'h19C17,4);
TASK_PP(16'h19C18,4);
TASK_PP(16'h19C19,4);
TASK_PP(16'h19C1A,4);
TASK_PP(16'h19C1B,4);
TASK_PP(16'h19C1C,4);
TASK_PP(16'h19C1D,4);
TASK_PP(16'h19C1E,4);
TASK_PP(16'h19C1F,4);
TASK_PP(16'h19C20,4);
TASK_PP(16'h19C21,4);
TASK_PP(16'h19C22,4);
TASK_PP(16'h19C23,4);
TASK_PP(16'h19C24,4);
TASK_PP(16'h19C25,4);
TASK_PP(16'h19C26,4);
TASK_PP(16'h19C27,4);
TASK_PP(16'h19C28,4);
TASK_PP(16'h19C29,4);
TASK_PP(16'h19C2A,4);
TASK_PP(16'h19C2B,4);
TASK_PP(16'h19C2C,4);
TASK_PP(16'h19C2D,4);
TASK_PP(16'h19C2E,4);
TASK_PP(16'h19C2F,4);
TASK_PP(16'h19C30,4);
TASK_PP(16'h19C31,4);
TASK_PP(16'h19C32,4);
TASK_PP(16'h19C33,4);
TASK_PP(16'h19C34,4);
TASK_PP(16'h19C35,4);
TASK_PP(16'h19C36,4);
TASK_PP(16'h19C37,4);
TASK_PP(16'h19C38,4);
TASK_PP(16'h19C39,4);
TASK_PP(16'h19C3A,4);
TASK_PP(16'h19C3B,4);
TASK_PP(16'h19C3C,4);
TASK_PP(16'h19C3D,4);
TASK_PP(16'h19C3E,4);
TASK_PP(16'h19C3F,4);
TASK_PP(16'h19C40,4);
TASK_PP(16'h19C41,4);
TASK_PP(16'h19C42,4);
TASK_PP(16'h19C43,4);
TASK_PP(16'h19C44,4);
TASK_PP(16'h19C45,4);
TASK_PP(16'h19C46,4);
TASK_PP(16'h19C47,4);
TASK_PP(16'h19C48,4);
TASK_PP(16'h19C49,4);
TASK_PP(16'h19C4A,4);
TASK_PP(16'h19C4B,4);
TASK_PP(16'h19C4C,4);
TASK_PP(16'h19C4D,4);
TASK_PP(16'h19C4E,4);
TASK_PP(16'h19C4F,4);
TASK_PP(16'h19C50,4);
TASK_PP(16'h19C51,4);
TASK_PP(16'h19C52,4);
TASK_PP(16'h19C53,4);
TASK_PP(16'h19C54,4);
TASK_PP(16'h19C55,4);
TASK_PP(16'h19C56,4);
TASK_PP(16'h19C57,4);
TASK_PP(16'h19C58,4);
TASK_PP(16'h19C59,4);
TASK_PP(16'h19C5A,4);
TASK_PP(16'h19C5B,4);
TASK_PP(16'h19C5C,4);
TASK_PP(16'h19C5D,4);
TASK_PP(16'h19C5E,4);
TASK_PP(16'h19C5F,4);
TASK_PP(16'h19C60,4);
TASK_PP(16'h19C61,4);
TASK_PP(16'h19C62,4);
TASK_PP(16'h19C63,4);
TASK_PP(16'h19C64,4);
TASK_PP(16'h19C65,4);
TASK_PP(16'h19C66,4);
TASK_PP(16'h19C67,4);
TASK_PP(16'h19C68,4);
TASK_PP(16'h19C69,4);
TASK_PP(16'h19C6A,4);
TASK_PP(16'h19C6B,4);
TASK_PP(16'h19C6C,4);
TASK_PP(16'h19C6D,4);
TASK_PP(16'h19C6E,4);
TASK_PP(16'h19C6F,4);
TASK_PP(16'h19C70,4);
TASK_PP(16'h19C71,4);
TASK_PP(16'h19C72,4);
TASK_PP(16'h19C73,4);
TASK_PP(16'h19C74,4);
TASK_PP(16'h19C75,4);
TASK_PP(16'h19C76,4);
TASK_PP(16'h19C77,4);
TASK_PP(16'h19C78,4);
TASK_PP(16'h19C79,4);
TASK_PP(16'h19C7A,4);
TASK_PP(16'h19C7B,4);
TASK_PP(16'h19C7C,4);
TASK_PP(16'h19C7D,4);
TASK_PP(16'h19C7E,4);
TASK_PP(16'h19C7F,4);
TASK_PP(16'h19C80,4);
TASK_PP(16'h19C81,4);
TASK_PP(16'h19C82,4);
TASK_PP(16'h19C83,4);
TASK_PP(16'h19C84,4);
TASK_PP(16'h19C85,4);
TASK_PP(16'h19C86,4);
TASK_PP(16'h19C87,4);
TASK_PP(16'h19C88,4);
TASK_PP(16'h19C89,4);
TASK_PP(16'h19C8A,4);
TASK_PP(16'h19C8B,4);
TASK_PP(16'h19C8C,4);
TASK_PP(16'h19C8D,4);
TASK_PP(16'h19C8E,4);
TASK_PP(16'h19C8F,4);
TASK_PP(16'h19C90,4);
TASK_PP(16'h19C91,4);
TASK_PP(16'h19C92,4);
TASK_PP(16'h19C93,4);
TASK_PP(16'h19C94,4);
TASK_PP(16'h19C95,4);
TASK_PP(16'h19C96,4);
TASK_PP(16'h19C97,4);
TASK_PP(16'h19C98,4);
TASK_PP(16'h19C99,4);
TASK_PP(16'h19C9A,4);
TASK_PP(16'h19C9B,4);
TASK_PP(16'h19C9C,4);
TASK_PP(16'h19C9D,4);
TASK_PP(16'h19C9E,4);
TASK_PP(16'h19C9F,4);
TASK_PP(16'h19CA0,4);
TASK_PP(16'h19CA1,4);
TASK_PP(16'h19CA2,4);
TASK_PP(16'h19CA3,4);
TASK_PP(16'h19CA4,4);
TASK_PP(16'h19CA5,4);
TASK_PP(16'h19CA6,4);
TASK_PP(16'h19CA7,4);
TASK_PP(16'h19CA8,4);
TASK_PP(16'h19CA9,4);
TASK_PP(16'h19CAA,4);
TASK_PP(16'h19CAB,4);
TASK_PP(16'h19CAC,4);
TASK_PP(16'h19CAD,4);
TASK_PP(16'h19CAE,4);
TASK_PP(16'h19CAF,4);
TASK_PP(16'h19CB0,4);
TASK_PP(16'h19CB1,4);
TASK_PP(16'h19CB2,4);
TASK_PP(16'h19CB3,4);
TASK_PP(16'h19CB4,4);
TASK_PP(16'h19CB5,4);
TASK_PP(16'h19CB6,4);
TASK_PP(16'h19CB7,4);
TASK_PP(16'h19CB8,4);
TASK_PP(16'h19CB9,4);
TASK_PP(16'h19CBA,4);
TASK_PP(16'h19CBB,4);
TASK_PP(16'h19CBC,4);
TASK_PP(16'h19CBD,4);
TASK_PP(16'h19CBE,4);
TASK_PP(16'h19CBF,4);
TASK_PP(16'h19CC0,4);
TASK_PP(16'h19CC1,4);
TASK_PP(16'h19CC2,4);
TASK_PP(16'h19CC3,4);
TASK_PP(16'h19CC4,4);
TASK_PP(16'h19CC5,4);
TASK_PP(16'h19CC6,4);
TASK_PP(16'h19CC7,4);
TASK_PP(16'h19CC8,4);
TASK_PP(16'h19CC9,4);
TASK_PP(16'h19CCA,4);
TASK_PP(16'h19CCB,4);
TASK_PP(16'h19CCC,4);
TASK_PP(16'h19CCD,4);
TASK_PP(16'h19CCE,4);
TASK_PP(16'h19CCF,4);
TASK_PP(16'h19CD0,4);
TASK_PP(16'h19CD1,4);
TASK_PP(16'h19CD2,4);
TASK_PP(16'h19CD3,4);
TASK_PP(16'h19CD4,4);
TASK_PP(16'h19CD5,4);
TASK_PP(16'h19CD6,4);
TASK_PP(16'h19CD7,4);
TASK_PP(16'h19CD8,4);
TASK_PP(16'h19CD9,4);
TASK_PP(16'h19CDA,4);
TASK_PP(16'h19CDB,4);
TASK_PP(16'h19CDC,4);
TASK_PP(16'h19CDD,4);
TASK_PP(16'h19CDE,4);
TASK_PP(16'h19CDF,4);
TASK_PP(16'h19CE0,4);
TASK_PP(16'h19CE1,4);
TASK_PP(16'h19CE2,4);
TASK_PP(16'h19CE3,4);
TASK_PP(16'h19CE4,4);
TASK_PP(16'h19CE5,4);
TASK_PP(16'h19CE6,4);
TASK_PP(16'h19CE7,4);
TASK_PP(16'h19CE8,4);
TASK_PP(16'h19CE9,4);
TASK_PP(16'h19CEA,4);
TASK_PP(16'h19CEB,4);
TASK_PP(16'h19CEC,4);
TASK_PP(16'h19CED,4);
TASK_PP(16'h19CEE,4);
TASK_PP(16'h19CEF,4);
TASK_PP(16'h19CF0,4);
TASK_PP(16'h19CF1,4);
TASK_PP(16'h19CF2,4);
TASK_PP(16'h19CF3,4);
TASK_PP(16'h19CF4,4);
TASK_PP(16'h19CF5,4);
TASK_PP(16'h19CF6,4);
TASK_PP(16'h19CF7,4);
TASK_PP(16'h19CF8,4);
TASK_PP(16'h19CF9,4);
TASK_PP(16'h19CFA,4);
TASK_PP(16'h19CFB,4);
TASK_PP(16'h19CFC,4);
TASK_PP(16'h19CFD,4);
TASK_PP(16'h19CFE,4);
TASK_PP(16'h19CFF,4);
TASK_PP(16'h19D00,4);
TASK_PP(16'h19D01,4);
TASK_PP(16'h19D02,4);
TASK_PP(16'h19D03,4);
TASK_PP(16'h19D04,4);
TASK_PP(16'h19D05,4);
TASK_PP(16'h19D06,4);
TASK_PP(16'h19D07,4);
TASK_PP(16'h19D08,4);
TASK_PP(16'h19D09,4);
TASK_PP(16'h19D0A,4);
TASK_PP(16'h19D0B,4);
TASK_PP(16'h19D0C,4);
TASK_PP(16'h19D0D,4);
TASK_PP(16'h19D0E,4);
TASK_PP(16'h19D0F,4);
TASK_PP(16'h19D10,4);
TASK_PP(16'h19D11,4);
TASK_PP(16'h19D12,4);
TASK_PP(16'h19D13,4);
TASK_PP(16'h19D14,4);
TASK_PP(16'h19D15,4);
TASK_PP(16'h19D16,4);
TASK_PP(16'h19D17,4);
TASK_PP(16'h19D18,4);
TASK_PP(16'h19D19,4);
TASK_PP(16'h19D1A,4);
TASK_PP(16'h19D1B,4);
TASK_PP(16'h19D1C,4);
TASK_PP(16'h19D1D,4);
TASK_PP(16'h19D1E,4);
TASK_PP(16'h19D1F,4);
TASK_PP(16'h19D20,4);
TASK_PP(16'h19D21,4);
TASK_PP(16'h19D22,4);
TASK_PP(16'h19D23,4);
TASK_PP(16'h19D24,4);
TASK_PP(16'h19D25,4);
TASK_PP(16'h19D26,4);
TASK_PP(16'h19D27,4);
TASK_PP(16'h19D28,4);
TASK_PP(16'h19D29,4);
TASK_PP(16'h19D2A,4);
TASK_PP(16'h19D2B,4);
TASK_PP(16'h19D2C,4);
TASK_PP(16'h19D2D,4);
TASK_PP(16'h19D2E,4);
TASK_PP(16'h19D2F,4);
TASK_PP(16'h19D30,4);
TASK_PP(16'h19D31,4);
TASK_PP(16'h19D32,4);
TASK_PP(16'h19D33,4);
TASK_PP(16'h19D34,4);
TASK_PP(16'h19D35,4);
TASK_PP(16'h19D36,4);
TASK_PP(16'h19D37,4);
TASK_PP(16'h19D38,4);
TASK_PP(16'h19D39,4);
TASK_PP(16'h19D3A,4);
TASK_PP(16'h19D3B,4);
TASK_PP(16'h19D3C,4);
TASK_PP(16'h19D3D,4);
TASK_PP(16'h19D3E,4);
TASK_PP(16'h19D3F,4);
TASK_PP(16'h19D40,4);
TASK_PP(16'h19D41,4);
TASK_PP(16'h19D42,4);
TASK_PP(16'h19D43,4);
TASK_PP(16'h19D44,4);
TASK_PP(16'h19D45,4);
TASK_PP(16'h19D46,4);
TASK_PP(16'h19D47,4);
TASK_PP(16'h19D48,4);
TASK_PP(16'h19D49,4);
TASK_PP(16'h19D4A,4);
TASK_PP(16'h19D4B,4);
TASK_PP(16'h19D4C,4);
TASK_PP(16'h19D4D,4);
TASK_PP(16'h19D4E,4);
TASK_PP(16'h19D4F,4);
TASK_PP(16'h19D50,4);
TASK_PP(16'h19D51,4);
TASK_PP(16'h19D52,4);
TASK_PP(16'h19D53,4);
TASK_PP(16'h19D54,4);
TASK_PP(16'h19D55,4);
TASK_PP(16'h19D56,4);
TASK_PP(16'h19D57,4);
TASK_PP(16'h19D58,4);
TASK_PP(16'h19D59,4);
TASK_PP(16'h19D5A,4);
TASK_PP(16'h19D5B,4);
TASK_PP(16'h19D5C,4);
TASK_PP(16'h19D5D,4);
TASK_PP(16'h19D5E,4);
TASK_PP(16'h19D5F,4);
TASK_PP(16'h19D60,4);
TASK_PP(16'h19D61,4);
TASK_PP(16'h19D62,4);
TASK_PP(16'h19D63,4);
TASK_PP(16'h19D64,4);
TASK_PP(16'h19D65,4);
TASK_PP(16'h19D66,4);
TASK_PP(16'h19D67,4);
TASK_PP(16'h19D68,4);
TASK_PP(16'h19D69,4);
TASK_PP(16'h19D6A,4);
TASK_PP(16'h19D6B,4);
TASK_PP(16'h19D6C,4);
TASK_PP(16'h19D6D,4);
TASK_PP(16'h19D6E,4);
TASK_PP(16'h19D6F,4);
TASK_PP(16'h19D70,4);
TASK_PP(16'h19D71,4);
TASK_PP(16'h19D72,4);
TASK_PP(16'h19D73,4);
TASK_PP(16'h19D74,4);
TASK_PP(16'h19D75,4);
TASK_PP(16'h19D76,4);
TASK_PP(16'h19D77,4);
TASK_PP(16'h19D78,4);
TASK_PP(16'h19D79,4);
TASK_PP(16'h19D7A,4);
TASK_PP(16'h19D7B,4);
TASK_PP(16'h19D7C,4);
TASK_PP(16'h19D7D,4);
TASK_PP(16'h19D7E,4);
TASK_PP(16'h19D7F,4);
TASK_PP(16'h19D80,4);
TASK_PP(16'h19D81,4);
TASK_PP(16'h19D82,4);
TASK_PP(16'h19D83,4);
TASK_PP(16'h19D84,4);
TASK_PP(16'h19D85,4);
TASK_PP(16'h19D86,4);
TASK_PP(16'h19D87,4);
TASK_PP(16'h19D88,4);
TASK_PP(16'h19D89,4);
TASK_PP(16'h19D8A,4);
TASK_PP(16'h19D8B,4);
TASK_PP(16'h19D8C,4);
TASK_PP(16'h19D8D,4);
TASK_PP(16'h19D8E,4);
TASK_PP(16'h19D8F,4);
TASK_PP(16'h19D90,4);
TASK_PP(16'h19D91,4);
TASK_PP(16'h19D92,4);
TASK_PP(16'h19D93,4);
TASK_PP(16'h19D94,4);
TASK_PP(16'h19D95,4);
TASK_PP(16'h19D96,4);
TASK_PP(16'h19D97,4);
TASK_PP(16'h19D98,4);
TASK_PP(16'h19D99,4);
TASK_PP(16'h19D9A,4);
TASK_PP(16'h19D9B,4);
TASK_PP(16'h19D9C,4);
TASK_PP(16'h19D9D,4);
TASK_PP(16'h19D9E,4);
TASK_PP(16'h19D9F,4);
TASK_PP(16'h19DA0,4);
TASK_PP(16'h19DA1,4);
TASK_PP(16'h19DA2,4);
TASK_PP(16'h19DA3,4);
TASK_PP(16'h19DA4,4);
TASK_PP(16'h19DA5,4);
TASK_PP(16'h19DA6,4);
TASK_PP(16'h19DA7,4);
TASK_PP(16'h19DA8,4);
TASK_PP(16'h19DA9,4);
TASK_PP(16'h19DAA,4);
TASK_PP(16'h19DAB,4);
TASK_PP(16'h19DAC,4);
TASK_PP(16'h19DAD,4);
TASK_PP(16'h19DAE,4);
TASK_PP(16'h19DAF,4);
TASK_PP(16'h19DB0,4);
TASK_PP(16'h19DB1,4);
TASK_PP(16'h19DB2,4);
TASK_PP(16'h19DB3,4);
TASK_PP(16'h19DB4,4);
TASK_PP(16'h19DB5,4);
TASK_PP(16'h19DB6,4);
TASK_PP(16'h19DB7,4);
TASK_PP(16'h19DB8,4);
TASK_PP(16'h19DB9,4);
TASK_PP(16'h19DBA,4);
TASK_PP(16'h19DBB,4);
TASK_PP(16'h19DBC,4);
TASK_PP(16'h19DBD,4);
TASK_PP(16'h19DBE,4);
TASK_PP(16'h19DBF,4);
TASK_PP(16'h19DC0,4);
TASK_PP(16'h19DC1,4);
TASK_PP(16'h19DC2,4);
TASK_PP(16'h19DC3,4);
TASK_PP(16'h19DC4,4);
TASK_PP(16'h19DC5,4);
TASK_PP(16'h19DC6,4);
TASK_PP(16'h19DC7,4);
TASK_PP(16'h19DC8,4);
TASK_PP(16'h19DC9,4);
TASK_PP(16'h19DCA,4);
TASK_PP(16'h19DCB,4);
TASK_PP(16'h19DCC,4);
TASK_PP(16'h19DCD,4);
TASK_PP(16'h19DCE,4);
TASK_PP(16'h19DCF,4);
TASK_PP(16'h19DD0,4);
TASK_PP(16'h19DD1,4);
TASK_PP(16'h19DD2,4);
TASK_PP(16'h19DD3,4);
TASK_PP(16'h19DD4,4);
TASK_PP(16'h19DD5,4);
TASK_PP(16'h19DD6,4);
TASK_PP(16'h19DD7,4);
TASK_PP(16'h19DD8,4);
TASK_PP(16'h19DD9,4);
TASK_PP(16'h19DDA,4);
TASK_PP(16'h19DDB,4);
TASK_PP(16'h19DDC,4);
TASK_PP(16'h19DDD,4);
TASK_PP(16'h19DDE,4);
TASK_PP(16'h19DDF,4);
TASK_PP(16'h19DE0,4);
TASK_PP(16'h19DE1,4);
TASK_PP(16'h19DE2,4);
TASK_PP(16'h19DE3,4);
TASK_PP(16'h19DE4,4);
TASK_PP(16'h19DE5,4);
TASK_PP(16'h19DE6,4);
TASK_PP(16'h19DE7,4);
TASK_PP(16'h19DE8,4);
TASK_PP(16'h19DE9,4);
TASK_PP(16'h19DEA,4);
TASK_PP(16'h19DEB,4);
TASK_PP(16'h19DEC,4);
TASK_PP(16'h19DED,4);
TASK_PP(16'h19DEE,4);
TASK_PP(16'h19DEF,4);
TASK_PP(16'h19DF0,4);
TASK_PP(16'h19DF1,4);
TASK_PP(16'h19DF2,4);
TASK_PP(16'h19DF3,4);
TASK_PP(16'h19DF4,4);
TASK_PP(16'h19DF5,4);
TASK_PP(16'h19DF6,4);
TASK_PP(16'h19DF7,4);
TASK_PP(16'h19DF8,4);
TASK_PP(16'h19DF9,4);
TASK_PP(16'h19DFA,4);
TASK_PP(16'h19DFB,4);
TASK_PP(16'h19DFC,4);
TASK_PP(16'h19DFD,4);
TASK_PP(16'h19DFE,4);
TASK_PP(16'h19DFF,4);
TASK_PP(16'h19E00,4);
TASK_PP(16'h19E01,4);
TASK_PP(16'h19E02,4);
TASK_PP(16'h19E03,4);
TASK_PP(16'h19E04,4);
TASK_PP(16'h19E05,4);
TASK_PP(16'h19E06,4);
TASK_PP(16'h19E07,4);
TASK_PP(16'h19E08,4);
TASK_PP(16'h19E09,4);
TASK_PP(16'h19E0A,4);
TASK_PP(16'h19E0B,4);
TASK_PP(16'h19E0C,4);
TASK_PP(16'h19E0D,4);
TASK_PP(16'h19E0E,4);
TASK_PP(16'h19E0F,4);
TASK_PP(16'h19E10,4);
TASK_PP(16'h19E11,4);
TASK_PP(16'h19E12,4);
TASK_PP(16'h19E13,4);
TASK_PP(16'h19E14,4);
TASK_PP(16'h19E15,4);
TASK_PP(16'h19E16,4);
TASK_PP(16'h19E17,4);
TASK_PP(16'h19E18,4);
TASK_PP(16'h19E19,4);
TASK_PP(16'h19E1A,4);
TASK_PP(16'h19E1B,4);
TASK_PP(16'h19E1C,4);
TASK_PP(16'h19E1D,4);
TASK_PP(16'h19E1E,4);
TASK_PP(16'h19E1F,4);
TASK_PP(16'h19E20,4);
TASK_PP(16'h19E21,4);
TASK_PP(16'h19E22,4);
TASK_PP(16'h19E23,4);
TASK_PP(16'h19E24,4);
TASK_PP(16'h19E25,4);
TASK_PP(16'h19E26,4);
TASK_PP(16'h19E27,4);
TASK_PP(16'h19E28,4);
TASK_PP(16'h19E29,4);
TASK_PP(16'h19E2A,4);
TASK_PP(16'h19E2B,4);
TASK_PP(16'h19E2C,4);
TASK_PP(16'h19E2D,4);
TASK_PP(16'h19E2E,4);
TASK_PP(16'h19E2F,4);
TASK_PP(16'h19E30,4);
TASK_PP(16'h19E31,4);
TASK_PP(16'h19E32,4);
TASK_PP(16'h19E33,4);
TASK_PP(16'h19E34,4);
TASK_PP(16'h19E35,4);
TASK_PP(16'h19E36,4);
TASK_PP(16'h19E37,4);
TASK_PP(16'h19E38,4);
TASK_PP(16'h19E39,4);
TASK_PP(16'h19E3A,4);
TASK_PP(16'h19E3B,4);
TASK_PP(16'h19E3C,4);
TASK_PP(16'h19E3D,4);
TASK_PP(16'h19E3E,4);
TASK_PP(16'h19E3F,4);
TASK_PP(16'h19E40,4);
TASK_PP(16'h19E41,4);
TASK_PP(16'h19E42,4);
TASK_PP(16'h19E43,4);
TASK_PP(16'h19E44,4);
TASK_PP(16'h19E45,4);
TASK_PP(16'h19E46,4);
TASK_PP(16'h19E47,4);
TASK_PP(16'h19E48,4);
TASK_PP(16'h19E49,4);
TASK_PP(16'h19E4A,4);
TASK_PP(16'h19E4B,4);
TASK_PP(16'h19E4C,4);
TASK_PP(16'h19E4D,4);
TASK_PP(16'h19E4E,4);
TASK_PP(16'h19E4F,4);
TASK_PP(16'h19E50,4);
TASK_PP(16'h19E51,4);
TASK_PP(16'h19E52,4);
TASK_PP(16'h19E53,4);
TASK_PP(16'h19E54,4);
TASK_PP(16'h19E55,4);
TASK_PP(16'h19E56,4);
TASK_PP(16'h19E57,4);
TASK_PP(16'h19E58,4);
TASK_PP(16'h19E59,4);
TASK_PP(16'h19E5A,4);
TASK_PP(16'h19E5B,4);
TASK_PP(16'h19E5C,4);
TASK_PP(16'h19E5D,4);
TASK_PP(16'h19E5E,4);
TASK_PP(16'h19E5F,4);
TASK_PP(16'h19E60,4);
TASK_PP(16'h19E61,4);
TASK_PP(16'h19E62,4);
TASK_PP(16'h19E63,4);
TASK_PP(16'h19E64,4);
TASK_PP(16'h19E65,4);
TASK_PP(16'h19E66,4);
TASK_PP(16'h19E67,4);
TASK_PP(16'h19E68,4);
TASK_PP(16'h19E69,4);
TASK_PP(16'h19E6A,4);
TASK_PP(16'h19E6B,4);
TASK_PP(16'h19E6C,4);
TASK_PP(16'h19E6D,4);
TASK_PP(16'h19E6E,4);
TASK_PP(16'h19E6F,4);
TASK_PP(16'h19E70,4);
TASK_PP(16'h19E71,4);
TASK_PP(16'h19E72,4);
TASK_PP(16'h19E73,4);
TASK_PP(16'h19E74,4);
TASK_PP(16'h19E75,4);
TASK_PP(16'h19E76,4);
TASK_PP(16'h19E77,4);
TASK_PP(16'h19E78,4);
TASK_PP(16'h19E79,4);
TASK_PP(16'h19E7A,4);
TASK_PP(16'h19E7B,4);
TASK_PP(16'h19E7C,4);
TASK_PP(16'h19E7D,4);
TASK_PP(16'h19E7E,4);
TASK_PP(16'h19E7F,4);
TASK_PP(16'h19E80,4);
TASK_PP(16'h19E81,4);
TASK_PP(16'h19E82,4);
TASK_PP(16'h19E83,4);
TASK_PP(16'h19E84,4);
TASK_PP(16'h19E85,4);
TASK_PP(16'h19E86,4);
TASK_PP(16'h19E87,4);
TASK_PP(16'h19E88,4);
TASK_PP(16'h19E89,4);
TASK_PP(16'h19E8A,4);
TASK_PP(16'h19E8B,4);
TASK_PP(16'h19E8C,4);
TASK_PP(16'h19E8D,4);
TASK_PP(16'h19E8E,4);
TASK_PP(16'h19E8F,4);
TASK_PP(16'h19E90,4);
TASK_PP(16'h19E91,4);
TASK_PP(16'h19E92,4);
TASK_PP(16'h19E93,4);
TASK_PP(16'h19E94,4);
TASK_PP(16'h19E95,4);
TASK_PP(16'h19E96,4);
TASK_PP(16'h19E97,4);
TASK_PP(16'h19E98,4);
TASK_PP(16'h19E99,4);
TASK_PP(16'h19E9A,4);
TASK_PP(16'h19E9B,4);
TASK_PP(16'h19E9C,4);
TASK_PP(16'h19E9D,4);
TASK_PP(16'h19E9E,4);
TASK_PP(16'h19E9F,4);
TASK_PP(16'h19EA0,4);
TASK_PP(16'h19EA1,4);
TASK_PP(16'h19EA2,4);
TASK_PP(16'h19EA3,4);
TASK_PP(16'h19EA4,4);
TASK_PP(16'h19EA5,4);
TASK_PP(16'h19EA6,4);
TASK_PP(16'h19EA7,4);
TASK_PP(16'h19EA8,4);
TASK_PP(16'h19EA9,4);
TASK_PP(16'h19EAA,4);
TASK_PP(16'h19EAB,4);
TASK_PP(16'h19EAC,4);
TASK_PP(16'h19EAD,4);
TASK_PP(16'h19EAE,4);
TASK_PP(16'h19EAF,4);
TASK_PP(16'h19EB0,4);
TASK_PP(16'h19EB1,4);
TASK_PP(16'h19EB2,4);
TASK_PP(16'h19EB3,4);
TASK_PP(16'h19EB4,4);
TASK_PP(16'h19EB5,4);
TASK_PP(16'h19EB6,4);
TASK_PP(16'h19EB7,4);
TASK_PP(16'h19EB8,4);
TASK_PP(16'h19EB9,4);
TASK_PP(16'h19EBA,4);
TASK_PP(16'h19EBB,4);
TASK_PP(16'h19EBC,4);
TASK_PP(16'h19EBD,4);
TASK_PP(16'h19EBE,4);
TASK_PP(16'h19EBF,4);
TASK_PP(16'h19EC0,4);
TASK_PP(16'h19EC1,4);
TASK_PP(16'h19EC2,4);
TASK_PP(16'h19EC3,4);
TASK_PP(16'h19EC4,4);
TASK_PP(16'h19EC5,4);
TASK_PP(16'h19EC6,4);
TASK_PP(16'h19EC7,4);
TASK_PP(16'h19EC8,4);
TASK_PP(16'h19EC9,4);
TASK_PP(16'h19ECA,4);
TASK_PP(16'h19ECB,4);
TASK_PP(16'h19ECC,4);
TASK_PP(16'h19ECD,4);
TASK_PP(16'h19ECE,4);
TASK_PP(16'h19ECF,4);
TASK_PP(16'h19ED0,4);
TASK_PP(16'h19ED1,4);
TASK_PP(16'h19ED2,4);
TASK_PP(16'h19ED3,4);
TASK_PP(16'h19ED4,4);
TASK_PP(16'h19ED5,4);
TASK_PP(16'h19ED6,4);
TASK_PP(16'h19ED7,4);
TASK_PP(16'h19ED8,4);
TASK_PP(16'h19ED9,4);
TASK_PP(16'h19EDA,4);
TASK_PP(16'h19EDB,4);
TASK_PP(16'h19EDC,4);
TASK_PP(16'h19EDD,4);
TASK_PP(16'h19EDE,4);
TASK_PP(16'h19EDF,4);
TASK_PP(16'h19EE0,4);
TASK_PP(16'h19EE1,4);
TASK_PP(16'h19EE2,4);
TASK_PP(16'h19EE3,4);
TASK_PP(16'h19EE4,4);
TASK_PP(16'h19EE5,4);
TASK_PP(16'h19EE6,4);
TASK_PP(16'h19EE7,4);
TASK_PP(16'h19EE8,4);
TASK_PP(16'h19EE9,4);
TASK_PP(16'h19EEA,4);
TASK_PP(16'h19EEB,4);
TASK_PP(16'h19EEC,4);
TASK_PP(16'h19EED,4);
TASK_PP(16'h19EEE,4);
TASK_PP(16'h19EEF,4);
TASK_PP(16'h19EF0,4);
TASK_PP(16'h19EF1,4);
TASK_PP(16'h19EF2,4);
TASK_PP(16'h19EF3,4);
TASK_PP(16'h19EF4,4);
TASK_PP(16'h19EF5,4);
TASK_PP(16'h19EF6,4);
TASK_PP(16'h19EF7,4);
TASK_PP(16'h19EF8,4);
TASK_PP(16'h19EF9,4);
TASK_PP(16'h19EFA,4);
TASK_PP(16'h19EFB,4);
TASK_PP(16'h19EFC,4);
TASK_PP(16'h19EFD,4);
TASK_PP(16'h19EFE,4);
TASK_PP(16'h19EFF,4);
TASK_PP(16'h19F00,4);
TASK_PP(16'h19F01,4);
TASK_PP(16'h19F02,4);
TASK_PP(16'h19F03,4);
TASK_PP(16'h19F04,4);
TASK_PP(16'h19F05,4);
TASK_PP(16'h19F06,4);
TASK_PP(16'h19F07,4);
TASK_PP(16'h19F08,4);
TASK_PP(16'h19F09,4);
TASK_PP(16'h19F0A,4);
TASK_PP(16'h19F0B,4);
TASK_PP(16'h19F0C,4);
TASK_PP(16'h19F0D,4);
TASK_PP(16'h19F0E,4);
TASK_PP(16'h19F0F,4);
TASK_PP(16'h19F10,4);
TASK_PP(16'h19F11,4);
TASK_PP(16'h19F12,4);
TASK_PP(16'h19F13,4);
TASK_PP(16'h19F14,4);
TASK_PP(16'h19F15,4);
TASK_PP(16'h19F16,4);
TASK_PP(16'h19F17,4);
TASK_PP(16'h19F18,4);
TASK_PP(16'h19F19,4);
TASK_PP(16'h19F1A,4);
TASK_PP(16'h19F1B,4);
TASK_PP(16'h19F1C,4);
TASK_PP(16'h19F1D,4);
TASK_PP(16'h19F1E,4);
TASK_PP(16'h19F1F,4);
TASK_PP(16'h19F20,4);
TASK_PP(16'h19F21,4);
TASK_PP(16'h19F22,4);
TASK_PP(16'h19F23,4);
TASK_PP(16'h19F24,4);
TASK_PP(16'h19F25,4);
TASK_PP(16'h19F26,4);
TASK_PP(16'h19F27,4);
TASK_PP(16'h19F28,4);
TASK_PP(16'h19F29,4);
TASK_PP(16'h19F2A,4);
TASK_PP(16'h19F2B,4);
TASK_PP(16'h19F2C,4);
TASK_PP(16'h19F2D,4);
TASK_PP(16'h19F2E,4);
TASK_PP(16'h19F2F,4);
TASK_PP(16'h19F30,4);
TASK_PP(16'h19F31,4);
TASK_PP(16'h19F32,4);
TASK_PP(16'h19F33,4);
TASK_PP(16'h19F34,4);
TASK_PP(16'h19F35,4);
TASK_PP(16'h19F36,4);
TASK_PP(16'h19F37,4);
TASK_PP(16'h19F38,4);
TASK_PP(16'h19F39,4);
TASK_PP(16'h19F3A,4);
TASK_PP(16'h19F3B,4);
TASK_PP(16'h19F3C,4);
TASK_PP(16'h19F3D,4);
TASK_PP(16'h19F3E,4);
TASK_PP(16'h19F3F,4);
TASK_PP(16'h19F40,4);
TASK_PP(16'h19F41,4);
TASK_PP(16'h19F42,4);
TASK_PP(16'h19F43,4);
TASK_PP(16'h19F44,4);
TASK_PP(16'h19F45,4);
TASK_PP(16'h19F46,4);
TASK_PP(16'h19F47,4);
TASK_PP(16'h19F48,4);
TASK_PP(16'h19F49,4);
TASK_PP(16'h19F4A,4);
TASK_PP(16'h19F4B,4);
TASK_PP(16'h19F4C,4);
TASK_PP(16'h19F4D,4);
TASK_PP(16'h19F4E,4);
TASK_PP(16'h19F4F,4);
TASK_PP(16'h19F50,4);
TASK_PP(16'h19F51,4);
TASK_PP(16'h19F52,4);
TASK_PP(16'h19F53,4);
TASK_PP(16'h19F54,4);
TASK_PP(16'h19F55,4);
TASK_PP(16'h19F56,4);
TASK_PP(16'h19F57,4);
TASK_PP(16'h19F58,4);
TASK_PP(16'h19F59,4);
TASK_PP(16'h19F5A,4);
TASK_PP(16'h19F5B,4);
TASK_PP(16'h19F5C,4);
TASK_PP(16'h19F5D,4);
TASK_PP(16'h19F5E,4);
TASK_PP(16'h19F5F,4);
TASK_PP(16'h19F60,4);
TASK_PP(16'h19F61,4);
TASK_PP(16'h19F62,4);
TASK_PP(16'h19F63,4);
TASK_PP(16'h19F64,4);
TASK_PP(16'h19F65,4);
TASK_PP(16'h19F66,4);
TASK_PP(16'h19F67,4);
TASK_PP(16'h19F68,4);
TASK_PP(16'h19F69,4);
TASK_PP(16'h19F6A,4);
TASK_PP(16'h19F6B,4);
TASK_PP(16'h19F6C,4);
TASK_PP(16'h19F6D,4);
TASK_PP(16'h19F6E,4);
TASK_PP(16'h19F6F,4);
TASK_PP(16'h19F70,4);
TASK_PP(16'h19F71,4);
TASK_PP(16'h19F72,4);
TASK_PP(16'h19F73,4);
TASK_PP(16'h19F74,4);
TASK_PP(16'h19F75,4);
TASK_PP(16'h19F76,4);
TASK_PP(16'h19F77,4);
TASK_PP(16'h19F78,4);
TASK_PP(16'h19F79,4);
TASK_PP(16'h19F7A,4);
TASK_PP(16'h19F7B,4);
TASK_PP(16'h19F7C,4);
TASK_PP(16'h19F7D,4);
TASK_PP(16'h19F7E,4);
TASK_PP(16'h19F7F,4);
TASK_PP(16'h19F80,4);
TASK_PP(16'h19F81,4);
TASK_PP(16'h19F82,4);
TASK_PP(16'h19F83,4);
TASK_PP(16'h19F84,4);
TASK_PP(16'h19F85,4);
TASK_PP(16'h19F86,4);
TASK_PP(16'h19F87,4);
TASK_PP(16'h19F88,4);
TASK_PP(16'h19F89,4);
TASK_PP(16'h19F8A,4);
TASK_PP(16'h19F8B,4);
TASK_PP(16'h19F8C,4);
TASK_PP(16'h19F8D,4);
TASK_PP(16'h19F8E,4);
TASK_PP(16'h19F8F,4);
TASK_PP(16'h19F90,4);
TASK_PP(16'h19F91,4);
TASK_PP(16'h19F92,4);
TASK_PP(16'h19F93,4);
TASK_PP(16'h19F94,4);
TASK_PP(16'h19F95,4);
TASK_PP(16'h19F96,4);
TASK_PP(16'h19F97,4);
TASK_PP(16'h19F98,4);
TASK_PP(16'h19F99,4);
TASK_PP(16'h19F9A,4);
TASK_PP(16'h19F9B,4);
TASK_PP(16'h19F9C,4);
TASK_PP(16'h19F9D,4);
TASK_PP(16'h19F9E,4);
TASK_PP(16'h19F9F,4);
TASK_PP(16'h19FA0,4);
TASK_PP(16'h19FA1,4);
TASK_PP(16'h19FA2,4);
TASK_PP(16'h19FA3,4);
TASK_PP(16'h19FA4,4);
TASK_PP(16'h19FA5,4);
TASK_PP(16'h19FA6,4);
TASK_PP(16'h19FA7,4);
TASK_PP(16'h19FA8,4);
TASK_PP(16'h19FA9,4);
TASK_PP(16'h19FAA,4);
TASK_PP(16'h19FAB,4);
TASK_PP(16'h19FAC,4);
TASK_PP(16'h19FAD,4);
TASK_PP(16'h19FAE,4);
TASK_PP(16'h19FAF,4);
TASK_PP(16'h19FB0,4);
TASK_PP(16'h19FB1,4);
TASK_PP(16'h19FB2,4);
TASK_PP(16'h19FB3,4);
TASK_PP(16'h19FB4,4);
TASK_PP(16'h19FB5,4);
TASK_PP(16'h19FB6,4);
TASK_PP(16'h19FB7,4);
TASK_PP(16'h19FB8,4);
TASK_PP(16'h19FB9,4);
TASK_PP(16'h19FBA,4);
TASK_PP(16'h19FBB,4);
TASK_PP(16'h19FBC,4);
TASK_PP(16'h19FBD,4);
TASK_PP(16'h19FBE,4);
TASK_PP(16'h19FBF,4);
TASK_PP(16'h19FC0,4);
TASK_PP(16'h19FC1,4);
TASK_PP(16'h19FC2,4);
TASK_PP(16'h19FC3,4);
TASK_PP(16'h19FC4,4);
TASK_PP(16'h19FC5,4);
TASK_PP(16'h19FC6,4);
TASK_PP(16'h19FC7,4);
TASK_PP(16'h19FC8,4);
TASK_PP(16'h19FC9,4);
TASK_PP(16'h19FCA,4);
TASK_PP(16'h19FCB,4);
TASK_PP(16'h19FCC,4);
TASK_PP(16'h19FCD,4);
TASK_PP(16'h19FCE,4);
TASK_PP(16'h19FCF,4);
TASK_PP(16'h19FD0,4);
TASK_PP(16'h19FD1,4);
TASK_PP(16'h19FD2,4);
TASK_PP(16'h19FD3,4);
TASK_PP(16'h19FD4,4);
TASK_PP(16'h19FD5,4);
TASK_PP(16'h19FD6,4);
TASK_PP(16'h19FD7,4);
TASK_PP(16'h19FD8,4);
TASK_PP(16'h19FD9,4);
TASK_PP(16'h19FDA,4);
TASK_PP(16'h19FDB,4);
TASK_PP(16'h19FDC,4);
TASK_PP(16'h19FDD,4);
TASK_PP(16'h19FDE,4);
TASK_PP(16'h19FDF,4);
TASK_PP(16'h19FE0,4);
TASK_PP(16'h19FE1,4);
TASK_PP(16'h19FE2,4);
TASK_PP(16'h19FE3,4);
TASK_PP(16'h19FE4,4);
TASK_PP(16'h19FE5,4);
TASK_PP(16'h19FE6,4);
TASK_PP(16'h19FE7,4);
TASK_PP(16'h19FE8,4);
TASK_PP(16'h19FE9,4);
TASK_PP(16'h19FEA,4);
TASK_PP(16'h19FEB,4);
TASK_PP(16'h19FEC,4);
TASK_PP(16'h19FED,4);
TASK_PP(16'h19FEE,4);
TASK_PP(16'h19FEF,4);
TASK_PP(16'h19FF0,4);
TASK_PP(16'h19FF1,4);
TASK_PP(16'h19FF2,4);
TASK_PP(16'h19FF3,4);
TASK_PP(16'h19FF4,4);
TASK_PP(16'h19FF5,4);
TASK_PP(16'h19FF6,4);
TASK_PP(16'h19FF7,4);
TASK_PP(16'h19FF8,4);
TASK_PP(16'h19FF9,4);
TASK_PP(16'h19FFA,4);
TASK_PP(16'h19FFB,4);
TASK_PP(16'h19FFC,4);
TASK_PP(16'h19FFD,4);
TASK_PP(16'h19FFE,4);
TASK_PP(16'h19FFF,4);
TASK_PP(16'h1A000,4);
TASK_PP(16'h1A001,4);
TASK_PP(16'h1A002,4);
TASK_PP(16'h1A003,4);
TASK_PP(16'h1A004,4);
TASK_PP(16'h1A005,4);
TASK_PP(16'h1A006,4);
TASK_PP(16'h1A007,4);
TASK_PP(16'h1A008,4);
TASK_PP(16'h1A009,4);
TASK_PP(16'h1A00A,4);
TASK_PP(16'h1A00B,4);
TASK_PP(16'h1A00C,4);
TASK_PP(16'h1A00D,4);
TASK_PP(16'h1A00E,4);
TASK_PP(16'h1A00F,4);
TASK_PP(16'h1A010,4);
TASK_PP(16'h1A011,4);
TASK_PP(16'h1A012,4);
TASK_PP(16'h1A013,4);
TASK_PP(16'h1A014,4);
TASK_PP(16'h1A015,4);
TASK_PP(16'h1A016,4);
TASK_PP(16'h1A017,4);
TASK_PP(16'h1A018,4);
TASK_PP(16'h1A019,4);
TASK_PP(16'h1A01A,4);
TASK_PP(16'h1A01B,4);
TASK_PP(16'h1A01C,4);
TASK_PP(16'h1A01D,4);
TASK_PP(16'h1A01E,4);
TASK_PP(16'h1A01F,4);
TASK_PP(16'h1A020,4);
TASK_PP(16'h1A021,4);
TASK_PP(16'h1A022,4);
TASK_PP(16'h1A023,4);
TASK_PP(16'h1A024,4);
TASK_PP(16'h1A025,4);
TASK_PP(16'h1A026,4);
TASK_PP(16'h1A027,4);
TASK_PP(16'h1A028,4);
TASK_PP(16'h1A029,4);
TASK_PP(16'h1A02A,4);
TASK_PP(16'h1A02B,4);
TASK_PP(16'h1A02C,4);
TASK_PP(16'h1A02D,4);
TASK_PP(16'h1A02E,4);
TASK_PP(16'h1A02F,4);
TASK_PP(16'h1A030,4);
TASK_PP(16'h1A031,4);
TASK_PP(16'h1A032,4);
TASK_PP(16'h1A033,4);
TASK_PP(16'h1A034,4);
TASK_PP(16'h1A035,4);
TASK_PP(16'h1A036,4);
TASK_PP(16'h1A037,4);
TASK_PP(16'h1A038,4);
TASK_PP(16'h1A039,4);
TASK_PP(16'h1A03A,4);
TASK_PP(16'h1A03B,4);
TASK_PP(16'h1A03C,4);
TASK_PP(16'h1A03D,4);
TASK_PP(16'h1A03E,4);
TASK_PP(16'h1A03F,4);
TASK_PP(16'h1A040,4);
TASK_PP(16'h1A041,4);
TASK_PP(16'h1A042,4);
TASK_PP(16'h1A043,4);
TASK_PP(16'h1A044,4);
TASK_PP(16'h1A045,4);
TASK_PP(16'h1A046,4);
TASK_PP(16'h1A047,4);
TASK_PP(16'h1A048,4);
TASK_PP(16'h1A049,4);
TASK_PP(16'h1A04A,4);
TASK_PP(16'h1A04B,4);
TASK_PP(16'h1A04C,4);
TASK_PP(16'h1A04D,4);
TASK_PP(16'h1A04E,4);
TASK_PP(16'h1A04F,4);
TASK_PP(16'h1A050,4);
TASK_PP(16'h1A051,4);
TASK_PP(16'h1A052,4);
TASK_PP(16'h1A053,4);
TASK_PP(16'h1A054,4);
TASK_PP(16'h1A055,4);
TASK_PP(16'h1A056,4);
TASK_PP(16'h1A057,4);
TASK_PP(16'h1A058,4);
TASK_PP(16'h1A059,4);
TASK_PP(16'h1A05A,4);
TASK_PP(16'h1A05B,4);
TASK_PP(16'h1A05C,4);
TASK_PP(16'h1A05D,4);
TASK_PP(16'h1A05E,4);
TASK_PP(16'h1A05F,4);
TASK_PP(16'h1A060,4);
TASK_PP(16'h1A061,4);
TASK_PP(16'h1A062,4);
TASK_PP(16'h1A063,4);
TASK_PP(16'h1A064,4);
TASK_PP(16'h1A065,4);
TASK_PP(16'h1A066,4);
TASK_PP(16'h1A067,4);
TASK_PP(16'h1A068,4);
TASK_PP(16'h1A069,4);
TASK_PP(16'h1A06A,4);
TASK_PP(16'h1A06B,4);
TASK_PP(16'h1A06C,4);
TASK_PP(16'h1A06D,4);
TASK_PP(16'h1A06E,4);
TASK_PP(16'h1A06F,4);
TASK_PP(16'h1A070,4);
TASK_PP(16'h1A071,4);
TASK_PP(16'h1A072,4);
TASK_PP(16'h1A073,4);
TASK_PP(16'h1A074,4);
TASK_PP(16'h1A075,4);
TASK_PP(16'h1A076,4);
TASK_PP(16'h1A077,4);
TASK_PP(16'h1A078,4);
TASK_PP(16'h1A079,4);
TASK_PP(16'h1A07A,4);
TASK_PP(16'h1A07B,4);
TASK_PP(16'h1A07C,4);
TASK_PP(16'h1A07D,4);
TASK_PP(16'h1A07E,4);
TASK_PP(16'h1A07F,4);
TASK_PP(16'h1A080,4);
TASK_PP(16'h1A081,4);
TASK_PP(16'h1A082,4);
TASK_PP(16'h1A083,4);
TASK_PP(16'h1A084,4);
TASK_PP(16'h1A085,4);
TASK_PP(16'h1A086,4);
TASK_PP(16'h1A087,4);
TASK_PP(16'h1A088,4);
TASK_PP(16'h1A089,4);
TASK_PP(16'h1A08A,4);
TASK_PP(16'h1A08B,4);
TASK_PP(16'h1A08C,4);
TASK_PP(16'h1A08D,4);
TASK_PP(16'h1A08E,4);
TASK_PP(16'h1A08F,4);
TASK_PP(16'h1A090,4);
TASK_PP(16'h1A091,4);
TASK_PP(16'h1A092,4);
TASK_PP(16'h1A093,4);
TASK_PP(16'h1A094,4);
TASK_PP(16'h1A095,4);
TASK_PP(16'h1A096,4);
TASK_PP(16'h1A097,4);
TASK_PP(16'h1A098,4);
TASK_PP(16'h1A099,4);
TASK_PP(16'h1A09A,4);
TASK_PP(16'h1A09B,4);
TASK_PP(16'h1A09C,4);
TASK_PP(16'h1A09D,4);
TASK_PP(16'h1A09E,4);
TASK_PP(16'h1A09F,4);
TASK_PP(16'h1A0A0,4);
TASK_PP(16'h1A0A1,4);
TASK_PP(16'h1A0A2,4);
TASK_PP(16'h1A0A3,4);
TASK_PP(16'h1A0A4,4);
TASK_PP(16'h1A0A5,4);
TASK_PP(16'h1A0A6,4);
TASK_PP(16'h1A0A7,4);
TASK_PP(16'h1A0A8,4);
TASK_PP(16'h1A0A9,4);
TASK_PP(16'h1A0AA,4);
TASK_PP(16'h1A0AB,4);
TASK_PP(16'h1A0AC,4);
TASK_PP(16'h1A0AD,4);
TASK_PP(16'h1A0AE,4);
TASK_PP(16'h1A0AF,4);
TASK_PP(16'h1A0B0,4);
TASK_PP(16'h1A0B1,4);
TASK_PP(16'h1A0B2,4);
TASK_PP(16'h1A0B3,4);
TASK_PP(16'h1A0B4,4);
TASK_PP(16'h1A0B5,4);
TASK_PP(16'h1A0B6,4);
TASK_PP(16'h1A0B7,4);
TASK_PP(16'h1A0B8,4);
TASK_PP(16'h1A0B9,4);
TASK_PP(16'h1A0BA,4);
TASK_PP(16'h1A0BB,4);
TASK_PP(16'h1A0BC,4);
TASK_PP(16'h1A0BD,4);
TASK_PP(16'h1A0BE,4);
TASK_PP(16'h1A0BF,4);
TASK_PP(16'h1A0C0,4);
TASK_PP(16'h1A0C1,4);
TASK_PP(16'h1A0C2,4);
TASK_PP(16'h1A0C3,4);
TASK_PP(16'h1A0C4,4);
TASK_PP(16'h1A0C5,4);
TASK_PP(16'h1A0C6,4);
TASK_PP(16'h1A0C7,4);
TASK_PP(16'h1A0C8,4);
TASK_PP(16'h1A0C9,4);
TASK_PP(16'h1A0CA,4);
TASK_PP(16'h1A0CB,4);
TASK_PP(16'h1A0CC,4);
TASK_PP(16'h1A0CD,4);
TASK_PP(16'h1A0CE,4);
TASK_PP(16'h1A0CF,4);
TASK_PP(16'h1A0D0,4);
TASK_PP(16'h1A0D1,4);
TASK_PP(16'h1A0D2,4);
TASK_PP(16'h1A0D3,4);
TASK_PP(16'h1A0D4,4);
TASK_PP(16'h1A0D5,4);
TASK_PP(16'h1A0D6,4);
TASK_PP(16'h1A0D7,4);
TASK_PP(16'h1A0D8,4);
TASK_PP(16'h1A0D9,4);
TASK_PP(16'h1A0DA,4);
TASK_PP(16'h1A0DB,4);
TASK_PP(16'h1A0DC,4);
TASK_PP(16'h1A0DD,4);
TASK_PP(16'h1A0DE,4);
TASK_PP(16'h1A0DF,4);
TASK_PP(16'h1A0E0,4);
TASK_PP(16'h1A0E1,4);
TASK_PP(16'h1A0E2,4);
TASK_PP(16'h1A0E3,4);
TASK_PP(16'h1A0E4,4);
TASK_PP(16'h1A0E5,4);
TASK_PP(16'h1A0E6,4);
TASK_PP(16'h1A0E7,4);
TASK_PP(16'h1A0E8,4);
TASK_PP(16'h1A0E9,4);
TASK_PP(16'h1A0EA,4);
TASK_PP(16'h1A0EB,4);
TASK_PP(16'h1A0EC,4);
TASK_PP(16'h1A0ED,4);
TASK_PP(16'h1A0EE,4);
TASK_PP(16'h1A0EF,4);
TASK_PP(16'h1A0F0,4);
TASK_PP(16'h1A0F1,4);
TASK_PP(16'h1A0F2,4);
TASK_PP(16'h1A0F3,4);
TASK_PP(16'h1A0F4,4);
TASK_PP(16'h1A0F5,4);
TASK_PP(16'h1A0F6,4);
TASK_PP(16'h1A0F7,4);
TASK_PP(16'h1A0F8,4);
TASK_PP(16'h1A0F9,4);
TASK_PP(16'h1A0FA,4);
TASK_PP(16'h1A0FB,4);
TASK_PP(16'h1A0FC,4);
TASK_PP(16'h1A0FD,4);
TASK_PP(16'h1A0FE,4);
TASK_PP(16'h1A0FF,4);
TASK_PP(16'h1A100,4);
TASK_PP(16'h1A101,4);
TASK_PP(16'h1A102,4);
TASK_PP(16'h1A103,4);
TASK_PP(16'h1A104,4);
TASK_PP(16'h1A105,4);
TASK_PP(16'h1A106,4);
TASK_PP(16'h1A107,4);
TASK_PP(16'h1A108,4);
TASK_PP(16'h1A109,4);
TASK_PP(16'h1A10A,4);
TASK_PP(16'h1A10B,4);
TASK_PP(16'h1A10C,4);
TASK_PP(16'h1A10D,4);
TASK_PP(16'h1A10E,4);
TASK_PP(16'h1A10F,4);
TASK_PP(16'h1A110,4);
TASK_PP(16'h1A111,4);
TASK_PP(16'h1A112,4);
TASK_PP(16'h1A113,4);
TASK_PP(16'h1A114,4);
TASK_PP(16'h1A115,4);
TASK_PP(16'h1A116,4);
TASK_PP(16'h1A117,4);
TASK_PP(16'h1A118,4);
TASK_PP(16'h1A119,4);
TASK_PP(16'h1A11A,4);
TASK_PP(16'h1A11B,4);
TASK_PP(16'h1A11C,4);
TASK_PP(16'h1A11D,4);
TASK_PP(16'h1A11E,4);
TASK_PP(16'h1A11F,4);
TASK_PP(16'h1A120,4);
TASK_PP(16'h1A121,4);
TASK_PP(16'h1A122,4);
TASK_PP(16'h1A123,4);
TASK_PP(16'h1A124,4);
TASK_PP(16'h1A125,4);
TASK_PP(16'h1A126,4);
TASK_PP(16'h1A127,4);
TASK_PP(16'h1A128,4);
TASK_PP(16'h1A129,4);
TASK_PP(16'h1A12A,4);
TASK_PP(16'h1A12B,4);
TASK_PP(16'h1A12C,4);
TASK_PP(16'h1A12D,4);
TASK_PP(16'h1A12E,4);
TASK_PP(16'h1A12F,4);
TASK_PP(16'h1A130,4);
TASK_PP(16'h1A131,4);
TASK_PP(16'h1A132,4);
TASK_PP(16'h1A133,4);
TASK_PP(16'h1A134,4);
TASK_PP(16'h1A135,4);
TASK_PP(16'h1A136,4);
TASK_PP(16'h1A137,4);
TASK_PP(16'h1A138,4);
TASK_PP(16'h1A139,4);
TASK_PP(16'h1A13A,4);
TASK_PP(16'h1A13B,4);
TASK_PP(16'h1A13C,4);
TASK_PP(16'h1A13D,4);
TASK_PP(16'h1A13E,4);
TASK_PP(16'h1A13F,4);
TASK_PP(16'h1A140,4);
TASK_PP(16'h1A141,4);
TASK_PP(16'h1A142,4);
TASK_PP(16'h1A143,4);
TASK_PP(16'h1A144,4);
TASK_PP(16'h1A145,4);
TASK_PP(16'h1A146,4);
TASK_PP(16'h1A147,4);
TASK_PP(16'h1A148,4);
TASK_PP(16'h1A149,4);
TASK_PP(16'h1A14A,4);
TASK_PP(16'h1A14B,4);
TASK_PP(16'h1A14C,4);
TASK_PP(16'h1A14D,4);
TASK_PP(16'h1A14E,4);
TASK_PP(16'h1A14F,4);
TASK_PP(16'h1A150,4);
TASK_PP(16'h1A151,4);
TASK_PP(16'h1A152,4);
TASK_PP(16'h1A153,4);
TASK_PP(16'h1A154,4);
TASK_PP(16'h1A155,4);
TASK_PP(16'h1A156,4);
TASK_PP(16'h1A157,4);
TASK_PP(16'h1A158,4);
TASK_PP(16'h1A159,4);
TASK_PP(16'h1A15A,4);
TASK_PP(16'h1A15B,4);
TASK_PP(16'h1A15C,4);
TASK_PP(16'h1A15D,4);
TASK_PP(16'h1A15E,4);
TASK_PP(16'h1A15F,4);
TASK_PP(16'h1A160,4);
TASK_PP(16'h1A161,4);
TASK_PP(16'h1A162,4);
TASK_PP(16'h1A163,4);
TASK_PP(16'h1A164,4);
TASK_PP(16'h1A165,4);
TASK_PP(16'h1A166,4);
TASK_PP(16'h1A167,4);
TASK_PP(16'h1A168,4);
TASK_PP(16'h1A169,4);
TASK_PP(16'h1A16A,4);
TASK_PP(16'h1A16B,4);
TASK_PP(16'h1A16C,4);
TASK_PP(16'h1A16D,4);
TASK_PP(16'h1A16E,4);
TASK_PP(16'h1A16F,4);
TASK_PP(16'h1A170,4);
TASK_PP(16'h1A171,4);
TASK_PP(16'h1A172,4);
TASK_PP(16'h1A173,4);
TASK_PP(16'h1A174,4);
TASK_PP(16'h1A175,4);
TASK_PP(16'h1A176,4);
TASK_PP(16'h1A177,4);
TASK_PP(16'h1A178,4);
TASK_PP(16'h1A179,4);
TASK_PP(16'h1A17A,4);
TASK_PP(16'h1A17B,4);
TASK_PP(16'h1A17C,4);
TASK_PP(16'h1A17D,4);
TASK_PP(16'h1A17E,4);
TASK_PP(16'h1A17F,4);
TASK_PP(16'h1A180,4);
TASK_PP(16'h1A181,4);
TASK_PP(16'h1A182,4);
TASK_PP(16'h1A183,4);
TASK_PP(16'h1A184,4);
TASK_PP(16'h1A185,4);
TASK_PP(16'h1A186,4);
TASK_PP(16'h1A187,4);
TASK_PP(16'h1A188,4);
TASK_PP(16'h1A189,4);
TASK_PP(16'h1A18A,4);
TASK_PP(16'h1A18B,4);
TASK_PP(16'h1A18C,4);
TASK_PP(16'h1A18D,4);
TASK_PP(16'h1A18E,4);
TASK_PP(16'h1A18F,4);
TASK_PP(16'h1A190,4);
TASK_PP(16'h1A191,4);
TASK_PP(16'h1A192,4);
TASK_PP(16'h1A193,4);
TASK_PP(16'h1A194,4);
TASK_PP(16'h1A195,4);
TASK_PP(16'h1A196,4);
TASK_PP(16'h1A197,4);
TASK_PP(16'h1A198,4);
TASK_PP(16'h1A199,4);
TASK_PP(16'h1A19A,4);
TASK_PP(16'h1A19B,4);
TASK_PP(16'h1A19C,4);
TASK_PP(16'h1A19D,4);
TASK_PP(16'h1A19E,4);
TASK_PP(16'h1A19F,4);
TASK_PP(16'h1A1A0,4);
TASK_PP(16'h1A1A1,4);
TASK_PP(16'h1A1A2,4);
TASK_PP(16'h1A1A3,4);
TASK_PP(16'h1A1A4,4);
TASK_PP(16'h1A1A5,4);
TASK_PP(16'h1A1A6,4);
TASK_PP(16'h1A1A7,4);
TASK_PP(16'h1A1A8,4);
TASK_PP(16'h1A1A9,4);
TASK_PP(16'h1A1AA,4);
TASK_PP(16'h1A1AB,4);
TASK_PP(16'h1A1AC,4);
TASK_PP(16'h1A1AD,4);
TASK_PP(16'h1A1AE,4);
TASK_PP(16'h1A1AF,4);
TASK_PP(16'h1A1B0,4);
TASK_PP(16'h1A1B1,4);
TASK_PP(16'h1A1B2,4);
TASK_PP(16'h1A1B3,4);
TASK_PP(16'h1A1B4,4);
TASK_PP(16'h1A1B5,4);
TASK_PP(16'h1A1B6,4);
TASK_PP(16'h1A1B7,4);
TASK_PP(16'h1A1B8,4);
TASK_PP(16'h1A1B9,4);
TASK_PP(16'h1A1BA,4);
TASK_PP(16'h1A1BB,4);
TASK_PP(16'h1A1BC,4);
TASK_PP(16'h1A1BD,4);
TASK_PP(16'h1A1BE,4);
TASK_PP(16'h1A1BF,4);
TASK_PP(16'h1A1C0,4);
TASK_PP(16'h1A1C1,4);
TASK_PP(16'h1A1C2,4);
TASK_PP(16'h1A1C3,4);
TASK_PP(16'h1A1C4,4);
TASK_PP(16'h1A1C5,4);
TASK_PP(16'h1A1C6,4);
TASK_PP(16'h1A1C7,4);
TASK_PP(16'h1A1C8,4);
TASK_PP(16'h1A1C9,4);
TASK_PP(16'h1A1CA,4);
TASK_PP(16'h1A1CB,4);
TASK_PP(16'h1A1CC,4);
TASK_PP(16'h1A1CD,4);
TASK_PP(16'h1A1CE,4);
TASK_PP(16'h1A1CF,4);
TASK_PP(16'h1A1D0,4);
TASK_PP(16'h1A1D1,4);
TASK_PP(16'h1A1D2,4);
TASK_PP(16'h1A1D3,4);
TASK_PP(16'h1A1D4,4);
TASK_PP(16'h1A1D5,4);
TASK_PP(16'h1A1D6,4);
TASK_PP(16'h1A1D7,4);
TASK_PP(16'h1A1D8,4);
TASK_PP(16'h1A1D9,4);
TASK_PP(16'h1A1DA,4);
TASK_PP(16'h1A1DB,4);
TASK_PP(16'h1A1DC,4);
TASK_PP(16'h1A1DD,4);
TASK_PP(16'h1A1DE,4);
TASK_PP(16'h1A1DF,4);
TASK_PP(16'h1A1E0,4);
TASK_PP(16'h1A1E1,4);
TASK_PP(16'h1A1E2,4);
TASK_PP(16'h1A1E3,4);
TASK_PP(16'h1A1E4,4);
TASK_PP(16'h1A1E5,4);
TASK_PP(16'h1A1E6,4);
TASK_PP(16'h1A1E7,4);
TASK_PP(16'h1A1E8,4);
TASK_PP(16'h1A1E9,4);
TASK_PP(16'h1A1EA,4);
TASK_PP(16'h1A1EB,4);
TASK_PP(16'h1A1EC,4);
TASK_PP(16'h1A1ED,4);
TASK_PP(16'h1A1EE,4);
TASK_PP(16'h1A1EF,4);
TASK_PP(16'h1A1F0,4);
TASK_PP(16'h1A1F1,4);
TASK_PP(16'h1A1F2,4);
TASK_PP(16'h1A1F3,4);
TASK_PP(16'h1A1F4,4);
TASK_PP(16'h1A1F5,4);
TASK_PP(16'h1A1F6,4);
TASK_PP(16'h1A1F7,4);
TASK_PP(16'h1A1F8,4);
TASK_PP(16'h1A1F9,4);
TASK_PP(16'h1A1FA,4);
TASK_PP(16'h1A1FB,4);
TASK_PP(16'h1A1FC,4);
TASK_PP(16'h1A1FD,4);
TASK_PP(16'h1A1FE,4);
TASK_PP(16'h1A1FF,4);
TASK_PP(16'h1A200,4);
TASK_PP(16'h1A201,4);
TASK_PP(16'h1A202,4);
TASK_PP(16'h1A203,4);
TASK_PP(16'h1A204,4);
TASK_PP(16'h1A205,4);
TASK_PP(16'h1A206,4);
TASK_PP(16'h1A207,4);
TASK_PP(16'h1A208,4);
TASK_PP(16'h1A209,4);
TASK_PP(16'h1A20A,4);
TASK_PP(16'h1A20B,4);
TASK_PP(16'h1A20C,4);
TASK_PP(16'h1A20D,4);
TASK_PP(16'h1A20E,4);
TASK_PP(16'h1A20F,4);
TASK_PP(16'h1A210,4);
TASK_PP(16'h1A211,4);
TASK_PP(16'h1A212,4);
TASK_PP(16'h1A213,4);
TASK_PP(16'h1A214,4);
TASK_PP(16'h1A215,4);
TASK_PP(16'h1A216,4);
TASK_PP(16'h1A217,4);
TASK_PP(16'h1A218,4);
TASK_PP(16'h1A219,4);
TASK_PP(16'h1A21A,4);
TASK_PP(16'h1A21B,4);
TASK_PP(16'h1A21C,4);
TASK_PP(16'h1A21D,4);
TASK_PP(16'h1A21E,4);
TASK_PP(16'h1A21F,4);
TASK_PP(16'h1A220,4);
TASK_PP(16'h1A221,4);
TASK_PP(16'h1A222,4);
TASK_PP(16'h1A223,4);
TASK_PP(16'h1A224,4);
TASK_PP(16'h1A225,4);
TASK_PP(16'h1A226,4);
TASK_PP(16'h1A227,4);
TASK_PP(16'h1A228,4);
TASK_PP(16'h1A229,4);
TASK_PP(16'h1A22A,4);
TASK_PP(16'h1A22B,4);
TASK_PP(16'h1A22C,4);
TASK_PP(16'h1A22D,4);
TASK_PP(16'h1A22E,4);
TASK_PP(16'h1A22F,4);
TASK_PP(16'h1A230,4);
TASK_PP(16'h1A231,4);
TASK_PP(16'h1A232,4);
TASK_PP(16'h1A233,4);
TASK_PP(16'h1A234,4);
TASK_PP(16'h1A235,4);
TASK_PP(16'h1A236,4);
TASK_PP(16'h1A237,4);
TASK_PP(16'h1A238,4);
TASK_PP(16'h1A239,4);
TASK_PP(16'h1A23A,4);
TASK_PP(16'h1A23B,4);
TASK_PP(16'h1A23C,4);
TASK_PP(16'h1A23D,4);
TASK_PP(16'h1A23E,4);
TASK_PP(16'h1A23F,4);
TASK_PP(16'h1A240,4);
TASK_PP(16'h1A241,4);
TASK_PP(16'h1A242,4);
TASK_PP(16'h1A243,4);
TASK_PP(16'h1A244,4);
TASK_PP(16'h1A245,4);
TASK_PP(16'h1A246,4);
TASK_PP(16'h1A247,4);
TASK_PP(16'h1A248,4);
TASK_PP(16'h1A249,4);
TASK_PP(16'h1A24A,4);
TASK_PP(16'h1A24B,4);
TASK_PP(16'h1A24C,4);
TASK_PP(16'h1A24D,4);
TASK_PP(16'h1A24E,4);
TASK_PP(16'h1A24F,4);
TASK_PP(16'h1A250,4);
TASK_PP(16'h1A251,4);
TASK_PP(16'h1A252,4);
TASK_PP(16'h1A253,4);
TASK_PP(16'h1A254,4);
TASK_PP(16'h1A255,4);
TASK_PP(16'h1A256,4);
TASK_PP(16'h1A257,4);
TASK_PP(16'h1A258,4);
TASK_PP(16'h1A259,4);
TASK_PP(16'h1A25A,4);
TASK_PP(16'h1A25B,4);
TASK_PP(16'h1A25C,4);
TASK_PP(16'h1A25D,4);
TASK_PP(16'h1A25E,4);
TASK_PP(16'h1A25F,4);
TASK_PP(16'h1A260,4);
TASK_PP(16'h1A261,4);
TASK_PP(16'h1A262,4);
TASK_PP(16'h1A263,4);
TASK_PP(16'h1A264,4);
TASK_PP(16'h1A265,4);
TASK_PP(16'h1A266,4);
TASK_PP(16'h1A267,4);
TASK_PP(16'h1A268,4);
TASK_PP(16'h1A269,4);
TASK_PP(16'h1A26A,4);
TASK_PP(16'h1A26B,4);
TASK_PP(16'h1A26C,4);
TASK_PP(16'h1A26D,4);
TASK_PP(16'h1A26E,4);
TASK_PP(16'h1A26F,4);
TASK_PP(16'h1A270,4);
TASK_PP(16'h1A271,4);
TASK_PP(16'h1A272,4);
TASK_PP(16'h1A273,4);
TASK_PP(16'h1A274,4);
TASK_PP(16'h1A275,4);
TASK_PP(16'h1A276,4);
TASK_PP(16'h1A277,4);
TASK_PP(16'h1A278,4);
TASK_PP(16'h1A279,4);
TASK_PP(16'h1A27A,4);
TASK_PP(16'h1A27B,4);
TASK_PP(16'h1A27C,4);
TASK_PP(16'h1A27D,4);
TASK_PP(16'h1A27E,4);
TASK_PP(16'h1A27F,4);
TASK_PP(16'h1A280,4);
TASK_PP(16'h1A281,4);
TASK_PP(16'h1A282,4);
TASK_PP(16'h1A283,4);
TASK_PP(16'h1A284,4);
TASK_PP(16'h1A285,4);
TASK_PP(16'h1A286,4);
TASK_PP(16'h1A287,4);
TASK_PP(16'h1A288,4);
TASK_PP(16'h1A289,4);
TASK_PP(16'h1A28A,4);
TASK_PP(16'h1A28B,4);
TASK_PP(16'h1A28C,4);
TASK_PP(16'h1A28D,4);
TASK_PP(16'h1A28E,4);
TASK_PP(16'h1A28F,4);
TASK_PP(16'h1A290,4);
TASK_PP(16'h1A291,4);
TASK_PP(16'h1A292,4);
TASK_PP(16'h1A293,4);
TASK_PP(16'h1A294,4);
TASK_PP(16'h1A295,4);
TASK_PP(16'h1A296,4);
TASK_PP(16'h1A297,4);
TASK_PP(16'h1A298,4);
TASK_PP(16'h1A299,4);
TASK_PP(16'h1A29A,4);
TASK_PP(16'h1A29B,4);
TASK_PP(16'h1A29C,4);
TASK_PP(16'h1A29D,4);
TASK_PP(16'h1A29E,4);
TASK_PP(16'h1A29F,4);
TASK_PP(16'h1A2A0,4);
TASK_PP(16'h1A2A1,4);
TASK_PP(16'h1A2A2,4);
TASK_PP(16'h1A2A3,4);
TASK_PP(16'h1A2A4,4);
TASK_PP(16'h1A2A5,4);
TASK_PP(16'h1A2A6,4);
TASK_PP(16'h1A2A7,4);
TASK_PP(16'h1A2A8,4);
TASK_PP(16'h1A2A9,4);
TASK_PP(16'h1A2AA,4);
TASK_PP(16'h1A2AB,4);
TASK_PP(16'h1A2AC,4);
TASK_PP(16'h1A2AD,4);
TASK_PP(16'h1A2AE,4);
TASK_PP(16'h1A2AF,4);
TASK_PP(16'h1A2B0,4);
TASK_PP(16'h1A2B1,4);
TASK_PP(16'h1A2B2,4);
TASK_PP(16'h1A2B3,4);
TASK_PP(16'h1A2B4,4);
TASK_PP(16'h1A2B5,4);
TASK_PP(16'h1A2B6,4);
TASK_PP(16'h1A2B7,4);
TASK_PP(16'h1A2B8,4);
TASK_PP(16'h1A2B9,4);
TASK_PP(16'h1A2BA,4);
TASK_PP(16'h1A2BB,4);
TASK_PP(16'h1A2BC,4);
TASK_PP(16'h1A2BD,4);
TASK_PP(16'h1A2BE,4);
TASK_PP(16'h1A2BF,4);
TASK_PP(16'h1A2C0,4);
TASK_PP(16'h1A2C1,4);
TASK_PP(16'h1A2C2,4);
TASK_PP(16'h1A2C3,4);
TASK_PP(16'h1A2C4,4);
TASK_PP(16'h1A2C5,4);
TASK_PP(16'h1A2C6,4);
TASK_PP(16'h1A2C7,4);
TASK_PP(16'h1A2C8,4);
TASK_PP(16'h1A2C9,4);
TASK_PP(16'h1A2CA,4);
TASK_PP(16'h1A2CB,4);
TASK_PP(16'h1A2CC,4);
TASK_PP(16'h1A2CD,4);
TASK_PP(16'h1A2CE,4);
TASK_PP(16'h1A2CF,4);
TASK_PP(16'h1A2D0,4);
TASK_PP(16'h1A2D1,4);
TASK_PP(16'h1A2D2,4);
TASK_PP(16'h1A2D3,4);
TASK_PP(16'h1A2D4,4);
TASK_PP(16'h1A2D5,4);
TASK_PP(16'h1A2D6,4);
TASK_PP(16'h1A2D7,4);
TASK_PP(16'h1A2D8,4);
TASK_PP(16'h1A2D9,4);
TASK_PP(16'h1A2DA,4);
TASK_PP(16'h1A2DB,4);
TASK_PP(16'h1A2DC,4);
TASK_PP(16'h1A2DD,4);
TASK_PP(16'h1A2DE,4);
TASK_PP(16'h1A2DF,4);
TASK_PP(16'h1A2E0,4);
TASK_PP(16'h1A2E1,4);
TASK_PP(16'h1A2E2,4);
TASK_PP(16'h1A2E3,4);
TASK_PP(16'h1A2E4,4);
TASK_PP(16'h1A2E5,4);
TASK_PP(16'h1A2E6,4);
TASK_PP(16'h1A2E7,4);
TASK_PP(16'h1A2E8,4);
TASK_PP(16'h1A2E9,4);
TASK_PP(16'h1A2EA,4);
TASK_PP(16'h1A2EB,4);
TASK_PP(16'h1A2EC,4);
TASK_PP(16'h1A2ED,4);
TASK_PP(16'h1A2EE,4);
TASK_PP(16'h1A2EF,4);
TASK_PP(16'h1A2F0,4);
TASK_PP(16'h1A2F1,4);
TASK_PP(16'h1A2F2,4);
TASK_PP(16'h1A2F3,4);
TASK_PP(16'h1A2F4,4);
TASK_PP(16'h1A2F5,4);
TASK_PP(16'h1A2F6,4);
TASK_PP(16'h1A2F7,4);
TASK_PP(16'h1A2F8,4);
TASK_PP(16'h1A2F9,4);
TASK_PP(16'h1A2FA,4);
TASK_PP(16'h1A2FB,4);
TASK_PP(16'h1A2FC,4);
TASK_PP(16'h1A2FD,4);
TASK_PP(16'h1A2FE,4);
TASK_PP(16'h1A2FF,4);
TASK_PP(16'h1A300,4);
TASK_PP(16'h1A301,4);
TASK_PP(16'h1A302,4);
TASK_PP(16'h1A303,4);
TASK_PP(16'h1A304,4);
TASK_PP(16'h1A305,4);
TASK_PP(16'h1A306,4);
TASK_PP(16'h1A307,4);
TASK_PP(16'h1A308,4);
TASK_PP(16'h1A309,4);
TASK_PP(16'h1A30A,4);
TASK_PP(16'h1A30B,4);
TASK_PP(16'h1A30C,4);
TASK_PP(16'h1A30D,4);
TASK_PP(16'h1A30E,4);
TASK_PP(16'h1A30F,4);
TASK_PP(16'h1A310,4);
TASK_PP(16'h1A311,4);
TASK_PP(16'h1A312,4);
TASK_PP(16'h1A313,4);
TASK_PP(16'h1A314,4);
TASK_PP(16'h1A315,4);
TASK_PP(16'h1A316,4);
TASK_PP(16'h1A317,4);
TASK_PP(16'h1A318,4);
TASK_PP(16'h1A319,4);
TASK_PP(16'h1A31A,4);
TASK_PP(16'h1A31B,4);
TASK_PP(16'h1A31C,4);
TASK_PP(16'h1A31D,4);
TASK_PP(16'h1A31E,4);
TASK_PP(16'h1A31F,4);
TASK_PP(16'h1A320,4);
TASK_PP(16'h1A321,4);
TASK_PP(16'h1A322,4);
TASK_PP(16'h1A323,4);
TASK_PP(16'h1A324,4);
TASK_PP(16'h1A325,4);
TASK_PP(16'h1A326,4);
TASK_PP(16'h1A327,4);
TASK_PP(16'h1A328,4);
TASK_PP(16'h1A329,4);
TASK_PP(16'h1A32A,4);
TASK_PP(16'h1A32B,4);
TASK_PP(16'h1A32C,4);
TASK_PP(16'h1A32D,4);
TASK_PP(16'h1A32E,4);
TASK_PP(16'h1A32F,4);
TASK_PP(16'h1A330,4);
TASK_PP(16'h1A331,4);
TASK_PP(16'h1A332,4);
TASK_PP(16'h1A333,4);
TASK_PP(16'h1A334,4);
TASK_PP(16'h1A335,4);
TASK_PP(16'h1A336,4);
TASK_PP(16'h1A337,4);
TASK_PP(16'h1A338,4);
TASK_PP(16'h1A339,4);
TASK_PP(16'h1A33A,4);
TASK_PP(16'h1A33B,4);
TASK_PP(16'h1A33C,4);
TASK_PP(16'h1A33D,4);
TASK_PP(16'h1A33E,4);
TASK_PP(16'h1A33F,4);
TASK_PP(16'h1A340,4);
TASK_PP(16'h1A341,4);
TASK_PP(16'h1A342,4);
TASK_PP(16'h1A343,4);
TASK_PP(16'h1A344,4);
TASK_PP(16'h1A345,4);
TASK_PP(16'h1A346,4);
TASK_PP(16'h1A347,4);
TASK_PP(16'h1A348,4);
TASK_PP(16'h1A349,4);
TASK_PP(16'h1A34A,4);
TASK_PP(16'h1A34B,4);
TASK_PP(16'h1A34C,4);
TASK_PP(16'h1A34D,4);
TASK_PP(16'h1A34E,4);
TASK_PP(16'h1A34F,4);
TASK_PP(16'h1A350,4);
TASK_PP(16'h1A351,4);
TASK_PP(16'h1A352,4);
TASK_PP(16'h1A353,4);
TASK_PP(16'h1A354,4);
TASK_PP(16'h1A355,4);
TASK_PP(16'h1A356,4);
TASK_PP(16'h1A357,4);
TASK_PP(16'h1A358,4);
TASK_PP(16'h1A359,4);
TASK_PP(16'h1A35A,4);
TASK_PP(16'h1A35B,4);
TASK_PP(16'h1A35C,4);
TASK_PP(16'h1A35D,4);
TASK_PP(16'h1A35E,4);
TASK_PP(16'h1A35F,4);
TASK_PP(16'h1A360,4);
TASK_PP(16'h1A361,4);
TASK_PP(16'h1A362,4);
TASK_PP(16'h1A363,4);
TASK_PP(16'h1A364,4);
TASK_PP(16'h1A365,4);
TASK_PP(16'h1A366,4);
TASK_PP(16'h1A367,4);
TASK_PP(16'h1A368,4);
TASK_PP(16'h1A369,4);
TASK_PP(16'h1A36A,4);
TASK_PP(16'h1A36B,4);
TASK_PP(16'h1A36C,4);
TASK_PP(16'h1A36D,4);
TASK_PP(16'h1A36E,4);
TASK_PP(16'h1A36F,4);
TASK_PP(16'h1A370,4);
TASK_PP(16'h1A371,4);
TASK_PP(16'h1A372,4);
TASK_PP(16'h1A373,4);
TASK_PP(16'h1A374,4);
TASK_PP(16'h1A375,4);
TASK_PP(16'h1A376,4);
TASK_PP(16'h1A377,4);
TASK_PP(16'h1A378,4);
TASK_PP(16'h1A379,4);
TASK_PP(16'h1A37A,4);
TASK_PP(16'h1A37B,4);
TASK_PP(16'h1A37C,4);
TASK_PP(16'h1A37D,4);
TASK_PP(16'h1A37E,4);
TASK_PP(16'h1A37F,4);
TASK_PP(16'h1A380,4);
TASK_PP(16'h1A381,4);
TASK_PP(16'h1A382,4);
TASK_PP(16'h1A383,4);
TASK_PP(16'h1A384,4);
TASK_PP(16'h1A385,4);
TASK_PP(16'h1A386,4);
TASK_PP(16'h1A387,4);
TASK_PP(16'h1A388,4);
TASK_PP(16'h1A389,4);
TASK_PP(16'h1A38A,4);
TASK_PP(16'h1A38B,4);
TASK_PP(16'h1A38C,4);
TASK_PP(16'h1A38D,4);
TASK_PP(16'h1A38E,4);
TASK_PP(16'h1A38F,4);
TASK_PP(16'h1A390,4);
TASK_PP(16'h1A391,4);
TASK_PP(16'h1A392,4);
TASK_PP(16'h1A393,4);
TASK_PP(16'h1A394,4);
TASK_PP(16'h1A395,4);
TASK_PP(16'h1A396,4);
TASK_PP(16'h1A397,4);
TASK_PP(16'h1A398,4);
TASK_PP(16'h1A399,4);
TASK_PP(16'h1A39A,4);
TASK_PP(16'h1A39B,4);
TASK_PP(16'h1A39C,4);
TASK_PP(16'h1A39D,4);
TASK_PP(16'h1A39E,4);
TASK_PP(16'h1A39F,4);
TASK_PP(16'h1A3A0,4);
TASK_PP(16'h1A3A1,4);
TASK_PP(16'h1A3A2,4);
TASK_PP(16'h1A3A3,4);
TASK_PP(16'h1A3A4,4);
TASK_PP(16'h1A3A5,4);
TASK_PP(16'h1A3A6,4);
TASK_PP(16'h1A3A7,4);
TASK_PP(16'h1A3A8,4);
TASK_PP(16'h1A3A9,4);
TASK_PP(16'h1A3AA,4);
TASK_PP(16'h1A3AB,4);
TASK_PP(16'h1A3AC,4);
TASK_PP(16'h1A3AD,4);
TASK_PP(16'h1A3AE,4);
TASK_PP(16'h1A3AF,4);
TASK_PP(16'h1A3B0,4);
TASK_PP(16'h1A3B1,4);
TASK_PP(16'h1A3B2,4);
TASK_PP(16'h1A3B3,4);
TASK_PP(16'h1A3B4,4);
TASK_PP(16'h1A3B5,4);
TASK_PP(16'h1A3B6,4);
TASK_PP(16'h1A3B7,4);
TASK_PP(16'h1A3B8,4);
TASK_PP(16'h1A3B9,4);
TASK_PP(16'h1A3BA,4);
TASK_PP(16'h1A3BB,4);
TASK_PP(16'h1A3BC,4);
TASK_PP(16'h1A3BD,4);
TASK_PP(16'h1A3BE,4);
TASK_PP(16'h1A3BF,4);
TASK_PP(16'h1A3C0,4);
TASK_PP(16'h1A3C1,4);
TASK_PP(16'h1A3C2,4);
TASK_PP(16'h1A3C3,4);
TASK_PP(16'h1A3C4,4);
TASK_PP(16'h1A3C5,4);
TASK_PP(16'h1A3C6,4);
TASK_PP(16'h1A3C7,4);
TASK_PP(16'h1A3C8,4);
TASK_PP(16'h1A3C9,4);
TASK_PP(16'h1A3CA,4);
TASK_PP(16'h1A3CB,4);
TASK_PP(16'h1A3CC,4);
TASK_PP(16'h1A3CD,4);
TASK_PP(16'h1A3CE,4);
TASK_PP(16'h1A3CF,4);
TASK_PP(16'h1A3D0,4);
TASK_PP(16'h1A3D1,4);
TASK_PP(16'h1A3D2,4);
TASK_PP(16'h1A3D3,4);
TASK_PP(16'h1A3D4,4);
TASK_PP(16'h1A3D5,4);
TASK_PP(16'h1A3D6,4);
TASK_PP(16'h1A3D7,4);
TASK_PP(16'h1A3D8,4);
TASK_PP(16'h1A3D9,4);
TASK_PP(16'h1A3DA,4);
TASK_PP(16'h1A3DB,4);
TASK_PP(16'h1A3DC,4);
TASK_PP(16'h1A3DD,4);
TASK_PP(16'h1A3DE,4);
TASK_PP(16'h1A3DF,4);
TASK_PP(16'h1A3E0,4);
TASK_PP(16'h1A3E1,4);
TASK_PP(16'h1A3E2,4);
TASK_PP(16'h1A3E3,4);
TASK_PP(16'h1A3E4,4);
TASK_PP(16'h1A3E5,4);
TASK_PP(16'h1A3E6,4);
TASK_PP(16'h1A3E7,4);
TASK_PP(16'h1A3E8,4);
TASK_PP(16'h1A3E9,4);
TASK_PP(16'h1A3EA,4);
TASK_PP(16'h1A3EB,4);
TASK_PP(16'h1A3EC,4);
TASK_PP(16'h1A3ED,4);
TASK_PP(16'h1A3EE,4);
TASK_PP(16'h1A3EF,4);
TASK_PP(16'h1A3F0,4);
TASK_PP(16'h1A3F1,4);
TASK_PP(16'h1A3F2,4);
TASK_PP(16'h1A3F3,4);
TASK_PP(16'h1A3F4,4);
TASK_PP(16'h1A3F5,4);
TASK_PP(16'h1A3F6,4);
TASK_PP(16'h1A3F7,4);
TASK_PP(16'h1A3F8,4);
TASK_PP(16'h1A3F9,4);
TASK_PP(16'h1A3FA,4);
TASK_PP(16'h1A3FB,4);
TASK_PP(16'h1A3FC,4);
TASK_PP(16'h1A3FD,4);
TASK_PP(16'h1A3FE,4);
TASK_PP(16'h1A3FF,4);
TASK_PP(16'h1A400,4);
TASK_PP(16'h1A401,4);
TASK_PP(16'h1A402,4);
TASK_PP(16'h1A403,4);
TASK_PP(16'h1A404,4);
TASK_PP(16'h1A405,4);
TASK_PP(16'h1A406,4);
TASK_PP(16'h1A407,4);
TASK_PP(16'h1A408,4);
TASK_PP(16'h1A409,4);
TASK_PP(16'h1A40A,4);
TASK_PP(16'h1A40B,4);
TASK_PP(16'h1A40C,4);
TASK_PP(16'h1A40D,4);
TASK_PP(16'h1A40E,4);
TASK_PP(16'h1A40F,4);
TASK_PP(16'h1A410,4);
TASK_PP(16'h1A411,4);
TASK_PP(16'h1A412,4);
TASK_PP(16'h1A413,4);
TASK_PP(16'h1A414,4);
TASK_PP(16'h1A415,4);
TASK_PP(16'h1A416,4);
TASK_PP(16'h1A417,4);
TASK_PP(16'h1A418,4);
TASK_PP(16'h1A419,4);
TASK_PP(16'h1A41A,4);
TASK_PP(16'h1A41B,4);
TASK_PP(16'h1A41C,4);
TASK_PP(16'h1A41D,4);
TASK_PP(16'h1A41E,4);
TASK_PP(16'h1A41F,4);
TASK_PP(16'h1A420,4);
TASK_PP(16'h1A421,4);
TASK_PP(16'h1A422,4);
TASK_PP(16'h1A423,4);
TASK_PP(16'h1A424,4);
TASK_PP(16'h1A425,4);
TASK_PP(16'h1A426,4);
TASK_PP(16'h1A427,4);
TASK_PP(16'h1A428,4);
TASK_PP(16'h1A429,4);
TASK_PP(16'h1A42A,4);
TASK_PP(16'h1A42B,4);
TASK_PP(16'h1A42C,4);
TASK_PP(16'h1A42D,4);
TASK_PP(16'h1A42E,4);
TASK_PP(16'h1A42F,4);
TASK_PP(16'h1A430,4);
TASK_PP(16'h1A431,4);
TASK_PP(16'h1A432,4);
TASK_PP(16'h1A433,4);
TASK_PP(16'h1A434,4);
TASK_PP(16'h1A435,4);
TASK_PP(16'h1A436,4);
TASK_PP(16'h1A437,4);
TASK_PP(16'h1A438,4);
TASK_PP(16'h1A439,4);
TASK_PP(16'h1A43A,4);
TASK_PP(16'h1A43B,4);
TASK_PP(16'h1A43C,4);
TASK_PP(16'h1A43D,4);
TASK_PP(16'h1A43E,4);
TASK_PP(16'h1A43F,4);
TASK_PP(16'h1A440,4);
TASK_PP(16'h1A441,4);
TASK_PP(16'h1A442,4);
TASK_PP(16'h1A443,4);
TASK_PP(16'h1A444,4);
TASK_PP(16'h1A445,4);
TASK_PP(16'h1A446,4);
TASK_PP(16'h1A447,4);
TASK_PP(16'h1A448,4);
TASK_PP(16'h1A449,4);
TASK_PP(16'h1A44A,4);
TASK_PP(16'h1A44B,4);
TASK_PP(16'h1A44C,4);
TASK_PP(16'h1A44D,4);
TASK_PP(16'h1A44E,4);
TASK_PP(16'h1A44F,4);
TASK_PP(16'h1A450,4);
TASK_PP(16'h1A451,4);
TASK_PP(16'h1A452,4);
TASK_PP(16'h1A453,4);
TASK_PP(16'h1A454,4);
TASK_PP(16'h1A455,4);
TASK_PP(16'h1A456,4);
TASK_PP(16'h1A457,4);
TASK_PP(16'h1A458,4);
TASK_PP(16'h1A459,4);
TASK_PP(16'h1A45A,4);
TASK_PP(16'h1A45B,4);
TASK_PP(16'h1A45C,4);
TASK_PP(16'h1A45D,4);
TASK_PP(16'h1A45E,4);
TASK_PP(16'h1A45F,4);
TASK_PP(16'h1A460,4);
TASK_PP(16'h1A461,4);
TASK_PP(16'h1A462,4);
TASK_PP(16'h1A463,4);
TASK_PP(16'h1A464,4);
TASK_PP(16'h1A465,4);
TASK_PP(16'h1A466,4);
TASK_PP(16'h1A467,4);
TASK_PP(16'h1A468,4);
TASK_PP(16'h1A469,4);
TASK_PP(16'h1A46A,4);
TASK_PP(16'h1A46B,4);
TASK_PP(16'h1A46C,4);
TASK_PP(16'h1A46D,4);
TASK_PP(16'h1A46E,4);
TASK_PP(16'h1A46F,4);
TASK_PP(16'h1A470,4);
TASK_PP(16'h1A471,4);
TASK_PP(16'h1A472,4);
TASK_PP(16'h1A473,4);
TASK_PP(16'h1A474,4);
TASK_PP(16'h1A475,4);
TASK_PP(16'h1A476,4);
TASK_PP(16'h1A477,4);
TASK_PP(16'h1A478,4);
TASK_PP(16'h1A479,4);
TASK_PP(16'h1A47A,4);
TASK_PP(16'h1A47B,4);
TASK_PP(16'h1A47C,4);
TASK_PP(16'h1A47D,4);
TASK_PP(16'h1A47E,4);
TASK_PP(16'h1A47F,4);
TASK_PP(16'h1A480,4);
TASK_PP(16'h1A481,4);
TASK_PP(16'h1A482,4);
TASK_PP(16'h1A483,4);
TASK_PP(16'h1A484,4);
TASK_PP(16'h1A485,4);
TASK_PP(16'h1A486,4);
TASK_PP(16'h1A487,4);
TASK_PP(16'h1A488,4);
TASK_PP(16'h1A489,4);
TASK_PP(16'h1A48A,4);
TASK_PP(16'h1A48B,4);
TASK_PP(16'h1A48C,4);
TASK_PP(16'h1A48D,4);
TASK_PP(16'h1A48E,4);
TASK_PP(16'h1A48F,4);
TASK_PP(16'h1A490,4);
TASK_PP(16'h1A491,4);
TASK_PP(16'h1A492,4);
TASK_PP(16'h1A493,4);
TASK_PP(16'h1A494,4);
TASK_PP(16'h1A495,4);
TASK_PP(16'h1A496,4);
TASK_PP(16'h1A497,4);
TASK_PP(16'h1A498,4);
TASK_PP(16'h1A499,4);
TASK_PP(16'h1A49A,4);
TASK_PP(16'h1A49B,4);
TASK_PP(16'h1A49C,4);
TASK_PP(16'h1A49D,4);
TASK_PP(16'h1A49E,4);
TASK_PP(16'h1A49F,4);
TASK_PP(16'h1A4A0,4);
TASK_PP(16'h1A4A1,4);
TASK_PP(16'h1A4A2,4);
TASK_PP(16'h1A4A3,4);
TASK_PP(16'h1A4A4,4);
TASK_PP(16'h1A4A5,4);
TASK_PP(16'h1A4A6,4);
TASK_PP(16'h1A4A7,4);
TASK_PP(16'h1A4A8,4);
TASK_PP(16'h1A4A9,4);
TASK_PP(16'h1A4AA,4);
TASK_PP(16'h1A4AB,4);
TASK_PP(16'h1A4AC,4);
TASK_PP(16'h1A4AD,4);
TASK_PP(16'h1A4AE,4);
TASK_PP(16'h1A4AF,4);
TASK_PP(16'h1A4B0,4);
TASK_PP(16'h1A4B1,4);
TASK_PP(16'h1A4B2,4);
TASK_PP(16'h1A4B3,4);
TASK_PP(16'h1A4B4,4);
TASK_PP(16'h1A4B5,4);
TASK_PP(16'h1A4B6,4);
TASK_PP(16'h1A4B7,4);
TASK_PP(16'h1A4B8,4);
TASK_PP(16'h1A4B9,4);
TASK_PP(16'h1A4BA,4);
TASK_PP(16'h1A4BB,4);
TASK_PP(16'h1A4BC,4);
TASK_PP(16'h1A4BD,4);
TASK_PP(16'h1A4BE,4);
TASK_PP(16'h1A4BF,4);
TASK_PP(16'h1A4C0,4);
TASK_PP(16'h1A4C1,4);
TASK_PP(16'h1A4C2,4);
TASK_PP(16'h1A4C3,4);
TASK_PP(16'h1A4C4,4);
TASK_PP(16'h1A4C5,4);
TASK_PP(16'h1A4C6,4);
TASK_PP(16'h1A4C7,4);
TASK_PP(16'h1A4C8,4);
TASK_PP(16'h1A4C9,4);
TASK_PP(16'h1A4CA,4);
TASK_PP(16'h1A4CB,4);
TASK_PP(16'h1A4CC,4);
TASK_PP(16'h1A4CD,4);
TASK_PP(16'h1A4CE,4);
TASK_PP(16'h1A4CF,4);
TASK_PP(16'h1A4D0,4);
TASK_PP(16'h1A4D1,4);
TASK_PP(16'h1A4D2,4);
TASK_PP(16'h1A4D3,4);
TASK_PP(16'h1A4D4,4);
TASK_PP(16'h1A4D5,4);
TASK_PP(16'h1A4D6,4);
TASK_PP(16'h1A4D7,4);
TASK_PP(16'h1A4D8,4);
TASK_PP(16'h1A4D9,4);
TASK_PP(16'h1A4DA,4);
TASK_PP(16'h1A4DB,4);
TASK_PP(16'h1A4DC,4);
TASK_PP(16'h1A4DD,4);
TASK_PP(16'h1A4DE,4);
TASK_PP(16'h1A4DF,4);
TASK_PP(16'h1A4E0,4);
TASK_PP(16'h1A4E1,4);
TASK_PP(16'h1A4E2,4);
TASK_PP(16'h1A4E3,4);
TASK_PP(16'h1A4E4,4);
TASK_PP(16'h1A4E5,4);
TASK_PP(16'h1A4E6,4);
TASK_PP(16'h1A4E7,4);
TASK_PP(16'h1A4E8,4);
TASK_PP(16'h1A4E9,4);
TASK_PP(16'h1A4EA,4);
TASK_PP(16'h1A4EB,4);
TASK_PP(16'h1A4EC,4);
TASK_PP(16'h1A4ED,4);
TASK_PP(16'h1A4EE,4);
TASK_PP(16'h1A4EF,4);
TASK_PP(16'h1A4F0,4);
TASK_PP(16'h1A4F1,4);
TASK_PP(16'h1A4F2,4);
TASK_PP(16'h1A4F3,4);
TASK_PP(16'h1A4F4,4);
TASK_PP(16'h1A4F5,4);
TASK_PP(16'h1A4F6,4);
TASK_PP(16'h1A4F7,4);
TASK_PP(16'h1A4F8,4);
TASK_PP(16'h1A4F9,4);
TASK_PP(16'h1A4FA,4);
TASK_PP(16'h1A4FB,4);
TASK_PP(16'h1A4FC,4);
TASK_PP(16'h1A4FD,4);
TASK_PP(16'h1A4FE,4);
TASK_PP(16'h1A4FF,4);
TASK_PP(16'h1A500,4);
TASK_PP(16'h1A501,4);
TASK_PP(16'h1A502,4);
TASK_PP(16'h1A503,4);
TASK_PP(16'h1A504,4);
TASK_PP(16'h1A505,4);
TASK_PP(16'h1A506,4);
TASK_PP(16'h1A507,4);
TASK_PP(16'h1A508,4);
TASK_PP(16'h1A509,4);
TASK_PP(16'h1A50A,4);
TASK_PP(16'h1A50B,4);
TASK_PP(16'h1A50C,4);
TASK_PP(16'h1A50D,4);
TASK_PP(16'h1A50E,4);
TASK_PP(16'h1A50F,4);
TASK_PP(16'h1A510,4);
TASK_PP(16'h1A511,4);
TASK_PP(16'h1A512,4);
TASK_PP(16'h1A513,4);
TASK_PP(16'h1A514,4);
TASK_PP(16'h1A515,4);
TASK_PP(16'h1A516,4);
TASK_PP(16'h1A517,4);
TASK_PP(16'h1A518,4);
TASK_PP(16'h1A519,4);
TASK_PP(16'h1A51A,4);
TASK_PP(16'h1A51B,4);
TASK_PP(16'h1A51C,4);
TASK_PP(16'h1A51D,4);
TASK_PP(16'h1A51E,4);
TASK_PP(16'h1A51F,4);
TASK_PP(16'h1A520,4);
TASK_PP(16'h1A521,4);
TASK_PP(16'h1A522,4);
TASK_PP(16'h1A523,4);
TASK_PP(16'h1A524,4);
TASK_PP(16'h1A525,4);
TASK_PP(16'h1A526,4);
TASK_PP(16'h1A527,4);
TASK_PP(16'h1A528,4);
TASK_PP(16'h1A529,4);
TASK_PP(16'h1A52A,4);
TASK_PP(16'h1A52B,4);
TASK_PP(16'h1A52C,4);
TASK_PP(16'h1A52D,4);
TASK_PP(16'h1A52E,4);
TASK_PP(16'h1A52F,4);
TASK_PP(16'h1A530,4);
TASK_PP(16'h1A531,4);
TASK_PP(16'h1A532,4);
TASK_PP(16'h1A533,4);
TASK_PP(16'h1A534,4);
TASK_PP(16'h1A535,4);
TASK_PP(16'h1A536,4);
TASK_PP(16'h1A537,4);
TASK_PP(16'h1A538,4);
TASK_PP(16'h1A539,4);
TASK_PP(16'h1A53A,4);
TASK_PP(16'h1A53B,4);
TASK_PP(16'h1A53C,4);
TASK_PP(16'h1A53D,4);
TASK_PP(16'h1A53E,4);
TASK_PP(16'h1A53F,4);
TASK_PP(16'h1A540,4);
TASK_PP(16'h1A541,4);
TASK_PP(16'h1A542,4);
TASK_PP(16'h1A543,4);
TASK_PP(16'h1A544,4);
TASK_PP(16'h1A545,4);
TASK_PP(16'h1A546,4);
TASK_PP(16'h1A547,4);
TASK_PP(16'h1A548,4);
TASK_PP(16'h1A549,4);
TASK_PP(16'h1A54A,4);
TASK_PP(16'h1A54B,4);
TASK_PP(16'h1A54C,4);
TASK_PP(16'h1A54D,4);
TASK_PP(16'h1A54E,4);
TASK_PP(16'h1A54F,4);
TASK_PP(16'h1A550,4);
TASK_PP(16'h1A551,4);
TASK_PP(16'h1A552,4);
TASK_PP(16'h1A553,4);
TASK_PP(16'h1A554,4);
TASK_PP(16'h1A555,4);
TASK_PP(16'h1A556,4);
TASK_PP(16'h1A557,4);
TASK_PP(16'h1A558,4);
TASK_PP(16'h1A559,4);
TASK_PP(16'h1A55A,4);
TASK_PP(16'h1A55B,4);
TASK_PP(16'h1A55C,4);
TASK_PP(16'h1A55D,4);
TASK_PP(16'h1A55E,4);
TASK_PP(16'h1A55F,4);
TASK_PP(16'h1A560,4);
TASK_PP(16'h1A561,4);
TASK_PP(16'h1A562,4);
TASK_PP(16'h1A563,4);
TASK_PP(16'h1A564,4);
TASK_PP(16'h1A565,4);
TASK_PP(16'h1A566,4);
TASK_PP(16'h1A567,4);
TASK_PP(16'h1A568,4);
TASK_PP(16'h1A569,4);
TASK_PP(16'h1A56A,4);
TASK_PP(16'h1A56B,4);
TASK_PP(16'h1A56C,4);
TASK_PP(16'h1A56D,4);
TASK_PP(16'h1A56E,4);
TASK_PP(16'h1A56F,4);
TASK_PP(16'h1A570,4);
TASK_PP(16'h1A571,4);
TASK_PP(16'h1A572,4);
TASK_PP(16'h1A573,4);
TASK_PP(16'h1A574,4);
TASK_PP(16'h1A575,4);
TASK_PP(16'h1A576,4);
TASK_PP(16'h1A577,4);
TASK_PP(16'h1A578,4);
TASK_PP(16'h1A579,4);
TASK_PP(16'h1A57A,4);
TASK_PP(16'h1A57B,4);
TASK_PP(16'h1A57C,4);
TASK_PP(16'h1A57D,4);
TASK_PP(16'h1A57E,4);
TASK_PP(16'h1A57F,4);
TASK_PP(16'h1A580,4);
TASK_PP(16'h1A581,4);
TASK_PP(16'h1A582,4);
TASK_PP(16'h1A583,4);
TASK_PP(16'h1A584,4);
TASK_PP(16'h1A585,4);
TASK_PP(16'h1A586,4);
TASK_PP(16'h1A587,4);
TASK_PP(16'h1A588,4);
TASK_PP(16'h1A589,4);
TASK_PP(16'h1A58A,4);
TASK_PP(16'h1A58B,4);
TASK_PP(16'h1A58C,4);
TASK_PP(16'h1A58D,4);
TASK_PP(16'h1A58E,4);
TASK_PP(16'h1A58F,4);
TASK_PP(16'h1A590,4);
TASK_PP(16'h1A591,4);
TASK_PP(16'h1A592,4);
TASK_PP(16'h1A593,4);
TASK_PP(16'h1A594,4);
TASK_PP(16'h1A595,4);
TASK_PP(16'h1A596,4);
TASK_PP(16'h1A597,4);
TASK_PP(16'h1A598,4);
TASK_PP(16'h1A599,4);
TASK_PP(16'h1A59A,4);
TASK_PP(16'h1A59B,4);
TASK_PP(16'h1A59C,4);
TASK_PP(16'h1A59D,4);
TASK_PP(16'h1A59E,4);
TASK_PP(16'h1A59F,4);
TASK_PP(16'h1A5A0,4);
TASK_PP(16'h1A5A1,4);
TASK_PP(16'h1A5A2,4);
TASK_PP(16'h1A5A3,4);
TASK_PP(16'h1A5A4,4);
TASK_PP(16'h1A5A5,4);
TASK_PP(16'h1A5A6,4);
TASK_PP(16'h1A5A7,4);
TASK_PP(16'h1A5A8,4);
TASK_PP(16'h1A5A9,4);
TASK_PP(16'h1A5AA,4);
TASK_PP(16'h1A5AB,4);
TASK_PP(16'h1A5AC,4);
TASK_PP(16'h1A5AD,4);
TASK_PP(16'h1A5AE,4);
TASK_PP(16'h1A5AF,4);
TASK_PP(16'h1A5B0,4);
TASK_PP(16'h1A5B1,4);
TASK_PP(16'h1A5B2,4);
TASK_PP(16'h1A5B3,4);
TASK_PP(16'h1A5B4,4);
TASK_PP(16'h1A5B5,4);
TASK_PP(16'h1A5B6,4);
TASK_PP(16'h1A5B7,4);
TASK_PP(16'h1A5B8,4);
TASK_PP(16'h1A5B9,4);
TASK_PP(16'h1A5BA,4);
TASK_PP(16'h1A5BB,4);
TASK_PP(16'h1A5BC,4);
TASK_PP(16'h1A5BD,4);
TASK_PP(16'h1A5BE,4);
TASK_PP(16'h1A5BF,4);
TASK_PP(16'h1A5C0,4);
TASK_PP(16'h1A5C1,4);
TASK_PP(16'h1A5C2,4);
TASK_PP(16'h1A5C3,4);
TASK_PP(16'h1A5C4,4);
TASK_PP(16'h1A5C5,4);
TASK_PP(16'h1A5C6,4);
TASK_PP(16'h1A5C7,4);
TASK_PP(16'h1A5C8,4);
TASK_PP(16'h1A5C9,4);
TASK_PP(16'h1A5CA,4);
TASK_PP(16'h1A5CB,4);
TASK_PP(16'h1A5CC,4);
TASK_PP(16'h1A5CD,4);
TASK_PP(16'h1A5CE,4);
TASK_PP(16'h1A5CF,4);
TASK_PP(16'h1A5D0,4);
TASK_PP(16'h1A5D1,4);
TASK_PP(16'h1A5D2,4);
TASK_PP(16'h1A5D3,4);
TASK_PP(16'h1A5D4,4);
TASK_PP(16'h1A5D5,4);
TASK_PP(16'h1A5D6,4);
TASK_PP(16'h1A5D7,4);
TASK_PP(16'h1A5D8,4);
TASK_PP(16'h1A5D9,4);
TASK_PP(16'h1A5DA,4);
TASK_PP(16'h1A5DB,4);
TASK_PP(16'h1A5DC,4);
TASK_PP(16'h1A5DD,4);
TASK_PP(16'h1A5DE,4);
TASK_PP(16'h1A5DF,4);
TASK_PP(16'h1A5E0,4);
TASK_PP(16'h1A5E1,4);
TASK_PP(16'h1A5E2,4);
TASK_PP(16'h1A5E3,4);
TASK_PP(16'h1A5E4,4);
TASK_PP(16'h1A5E5,4);
TASK_PP(16'h1A5E6,4);
TASK_PP(16'h1A5E7,4);
TASK_PP(16'h1A5E8,4);
TASK_PP(16'h1A5E9,4);
TASK_PP(16'h1A5EA,4);
TASK_PP(16'h1A5EB,4);
TASK_PP(16'h1A5EC,4);
TASK_PP(16'h1A5ED,4);
TASK_PP(16'h1A5EE,4);
TASK_PP(16'h1A5EF,4);
TASK_PP(16'h1A5F0,4);
TASK_PP(16'h1A5F1,4);
TASK_PP(16'h1A5F2,4);
TASK_PP(16'h1A5F3,4);
TASK_PP(16'h1A5F4,4);
TASK_PP(16'h1A5F5,4);
TASK_PP(16'h1A5F6,4);
TASK_PP(16'h1A5F7,4);
TASK_PP(16'h1A5F8,4);
TASK_PP(16'h1A5F9,4);
TASK_PP(16'h1A5FA,4);
TASK_PP(16'h1A5FB,4);
TASK_PP(16'h1A5FC,4);
TASK_PP(16'h1A5FD,4);
TASK_PP(16'h1A5FE,4);
TASK_PP(16'h1A5FF,4);
TASK_PP(16'h1A600,4);
TASK_PP(16'h1A601,4);
TASK_PP(16'h1A602,4);
TASK_PP(16'h1A603,4);
TASK_PP(16'h1A604,4);
TASK_PP(16'h1A605,4);
TASK_PP(16'h1A606,4);
TASK_PP(16'h1A607,4);
TASK_PP(16'h1A608,4);
TASK_PP(16'h1A609,4);
TASK_PP(16'h1A60A,4);
TASK_PP(16'h1A60B,4);
TASK_PP(16'h1A60C,4);
TASK_PP(16'h1A60D,4);
TASK_PP(16'h1A60E,4);
TASK_PP(16'h1A60F,4);
TASK_PP(16'h1A610,4);
TASK_PP(16'h1A611,4);
TASK_PP(16'h1A612,4);
TASK_PP(16'h1A613,4);
TASK_PP(16'h1A614,4);
TASK_PP(16'h1A615,4);
TASK_PP(16'h1A616,4);
TASK_PP(16'h1A617,4);
TASK_PP(16'h1A618,4);
TASK_PP(16'h1A619,4);
TASK_PP(16'h1A61A,4);
TASK_PP(16'h1A61B,4);
TASK_PP(16'h1A61C,4);
TASK_PP(16'h1A61D,4);
TASK_PP(16'h1A61E,4);
TASK_PP(16'h1A61F,4);
TASK_PP(16'h1A620,4);
TASK_PP(16'h1A621,4);
TASK_PP(16'h1A622,4);
TASK_PP(16'h1A623,4);
TASK_PP(16'h1A624,4);
TASK_PP(16'h1A625,4);
TASK_PP(16'h1A626,4);
TASK_PP(16'h1A627,4);
TASK_PP(16'h1A628,4);
TASK_PP(16'h1A629,4);
TASK_PP(16'h1A62A,4);
TASK_PP(16'h1A62B,4);
TASK_PP(16'h1A62C,4);
TASK_PP(16'h1A62D,4);
TASK_PP(16'h1A62E,4);
TASK_PP(16'h1A62F,4);
TASK_PP(16'h1A630,4);
TASK_PP(16'h1A631,4);
TASK_PP(16'h1A632,4);
TASK_PP(16'h1A633,4);
TASK_PP(16'h1A634,4);
TASK_PP(16'h1A635,4);
TASK_PP(16'h1A636,4);
TASK_PP(16'h1A637,4);
TASK_PP(16'h1A638,4);
TASK_PP(16'h1A639,4);
TASK_PP(16'h1A63A,4);
TASK_PP(16'h1A63B,4);
TASK_PP(16'h1A63C,4);
TASK_PP(16'h1A63D,4);
TASK_PP(16'h1A63E,4);
TASK_PP(16'h1A63F,4);
TASK_PP(16'h1A640,4);
TASK_PP(16'h1A641,4);
TASK_PP(16'h1A642,4);
TASK_PP(16'h1A643,4);
TASK_PP(16'h1A644,4);
TASK_PP(16'h1A645,4);
TASK_PP(16'h1A646,4);
TASK_PP(16'h1A647,4);
TASK_PP(16'h1A648,4);
TASK_PP(16'h1A649,4);
TASK_PP(16'h1A64A,4);
TASK_PP(16'h1A64B,4);
TASK_PP(16'h1A64C,4);
TASK_PP(16'h1A64D,4);
TASK_PP(16'h1A64E,4);
TASK_PP(16'h1A64F,4);
TASK_PP(16'h1A650,4);
TASK_PP(16'h1A651,4);
TASK_PP(16'h1A652,4);
TASK_PP(16'h1A653,4);
TASK_PP(16'h1A654,4);
TASK_PP(16'h1A655,4);
TASK_PP(16'h1A656,4);
TASK_PP(16'h1A657,4);
TASK_PP(16'h1A658,4);
TASK_PP(16'h1A659,4);
TASK_PP(16'h1A65A,4);
TASK_PP(16'h1A65B,4);
TASK_PP(16'h1A65C,4);
TASK_PP(16'h1A65D,4);
TASK_PP(16'h1A65E,4);
TASK_PP(16'h1A65F,4);
TASK_PP(16'h1A660,4);
TASK_PP(16'h1A661,4);
TASK_PP(16'h1A662,4);
TASK_PP(16'h1A663,4);
TASK_PP(16'h1A664,4);
TASK_PP(16'h1A665,4);
TASK_PP(16'h1A666,4);
TASK_PP(16'h1A667,4);
TASK_PP(16'h1A668,4);
TASK_PP(16'h1A669,4);
TASK_PP(16'h1A66A,4);
TASK_PP(16'h1A66B,4);
TASK_PP(16'h1A66C,4);
TASK_PP(16'h1A66D,4);
TASK_PP(16'h1A66E,4);
TASK_PP(16'h1A66F,4);
TASK_PP(16'h1A670,4);
TASK_PP(16'h1A671,4);
TASK_PP(16'h1A672,4);
TASK_PP(16'h1A673,4);
TASK_PP(16'h1A674,4);
TASK_PP(16'h1A675,4);
TASK_PP(16'h1A676,4);
TASK_PP(16'h1A677,4);
TASK_PP(16'h1A678,4);
TASK_PP(16'h1A679,4);
TASK_PP(16'h1A67A,4);
TASK_PP(16'h1A67B,4);
TASK_PP(16'h1A67C,4);
TASK_PP(16'h1A67D,4);
TASK_PP(16'h1A67E,4);
TASK_PP(16'h1A67F,4);
TASK_PP(16'h1A680,4);
TASK_PP(16'h1A681,4);
TASK_PP(16'h1A682,4);
TASK_PP(16'h1A683,4);
TASK_PP(16'h1A684,4);
TASK_PP(16'h1A685,4);
TASK_PP(16'h1A686,4);
TASK_PP(16'h1A687,4);
TASK_PP(16'h1A688,4);
TASK_PP(16'h1A689,4);
TASK_PP(16'h1A68A,4);
TASK_PP(16'h1A68B,4);
TASK_PP(16'h1A68C,4);
TASK_PP(16'h1A68D,4);
TASK_PP(16'h1A68E,4);
TASK_PP(16'h1A68F,4);
TASK_PP(16'h1A690,4);
TASK_PP(16'h1A691,4);
TASK_PP(16'h1A692,4);
TASK_PP(16'h1A693,4);
TASK_PP(16'h1A694,4);
TASK_PP(16'h1A695,4);
TASK_PP(16'h1A696,4);
TASK_PP(16'h1A697,4);
TASK_PP(16'h1A698,4);
TASK_PP(16'h1A699,4);
TASK_PP(16'h1A69A,4);
TASK_PP(16'h1A69B,4);
TASK_PP(16'h1A69C,4);
TASK_PP(16'h1A69D,4);
TASK_PP(16'h1A69E,4);
TASK_PP(16'h1A69F,4);
TASK_PP(16'h1A6A0,4);
TASK_PP(16'h1A6A1,4);
TASK_PP(16'h1A6A2,4);
TASK_PP(16'h1A6A3,4);
TASK_PP(16'h1A6A4,4);
TASK_PP(16'h1A6A5,4);
TASK_PP(16'h1A6A6,4);
TASK_PP(16'h1A6A7,4);
TASK_PP(16'h1A6A8,4);
TASK_PP(16'h1A6A9,4);
TASK_PP(16'h1A6AA,4);
TASK_PP(16'h1A6AB,4);
TASK_PP(16'h1A6AC,4);
TASK_PP(16'h1A6AD,4);
TASK_PP(16'h1A6AE,4);
TASK_PP(16'h1A6AF,4);
TASK_PP(16'h1A6B0,4);
TASK_PP(16'h1A6B1,4);
TASK_PP(16'h1A6B2,4);
TASK_PP(16'h1A6B3,4);
TASK_PP(16'h1A6B4,4);
TASK_PP(16'h1A6B5,4);
TASK_PP(16'h1A6B6,4);
TASK_PP(16'h1A6B7,4);
TASK_PP(16'h1A6B8,4);
TASK_PP(16'h1A6B9,4);
TASK_PP(16'h1A6BA,4);
TASK_PP(16'h1A6BB,4);
TASK_PP(16'h1A6BC,4);
TASK_PP(16'h1A6BD,4);
TASK_PP(16'h1A6BE,4);
TASK_PP(16'h1A6BF,4);
TASK_PP(16'h1A6C0,4);
TASK_PP(16'h1A6C1,4);
TASK_PP(16'h1A6C2,4);
TASK_PP(16'h1A6C3,4);
TASK_PP(16'h1A6C4,4);
TASK_PP(16'h1A6C5,4);
TASK_PP(16'h1A6C6,4);
TASK_PP(16'h1A6C7,4);
TASK_PP(16'h1A6C8,4);
TASK_PP(16'h1A6C9,4);
TASK_PP(16'h1A6CA,4);
TASK_PP(16'h1A6CB,4);
TASK_PP(16'h1A6CC,4);
TASK_PP(16'h1A6CD,4);
TASK_PP(16'h1A6CE,4);
TASK_PP(16'h1A6CF,4);
TASK_PP(16'h1A6D0,4);
TASK_PP(16'h1A6D1,4);
TASK_PP(16'h1A6D2,4);
TASK_PP(16'h1A6D3,4);
TASK_PP(16'h1A6D4,4);
TASK_PP(16'h1A6D5,4);
TASK_PP(16'h1A6D6,4);
TASK_PP(16'h1A6D7,4);
TASK_PP(16'h1A6D8,4);
TASK_PP(16'h1A6D9,4);
TASK_PP(16'h1A6DA,4);
TASK_PP(16'h1A6DB,4);
TASK_PP(16'h1A6DC,4);
TASK_PP(16'h1A6DD,4);
TASK_PP(16'h1A6DE,4);
TASK_PP(16'h1A6DF,4);
TASK_PP(16'h1A6E0,4);
TASK_PP(16'h1A6E1,4);
TASK_PP(16'h1A6E2,4);
TASK_PP(16'h1A6E3,4);
TASK_PP(16'h1A6E4,4);
TASK_PP(16'h1A6E5,4);
TASK_PP(16'h1A6E6,4);
TASK_PP(16'h1A6E7,4);
TASK_PP(16'h1A6E8,4);
TASK_PP(16'h1A6E9,4);
TASK_PP(16'h1A6EA,4);
TASK_PP(16'h1A6EB,4);
TASK_PP(16'h1A6EC,4);
TASK_PP(16'h1A6ED,4);
TASK_PP(16'h1A6EE,4);
TASK_PP(16'h1A6EF,4);
TASK_PP(16'h1A6F0,4);
TASK_PP(16'h1A6F1,4);
TASK_PP(16'h1A6F2,4);
TASK_PP(16'h1A6F3,4);
TASK_PP(16'h1A6F4,4);
TASK_PP(16'h1A6F5,4);
TASK_PP(16'h1A6F6,4);
TASK_PP(16'h1A6F7,4);
TASK_PP(16'h1A6F8,4);
TASK_PP(16'h1A6F9,4);
TASK_PP(16'h1A6FA,4);
TASK_PP(16'h1A6FB,4);
TASK_PP(16'h1A6FC,4);
TASK_PP(16'h1A6FD,4);
TASK_PP(16'h1A6FE,4);
TASK_PP(16'h1A6FF,4);
TASK_PP(16'h1A700,4);
TASK_PP(16'h1A701,4);
TASK_PP(16'h1A702,4);
TASK_PP(16'h1A703,4);
TASK_PP(16'h1A704,4);
TASK_PP(16'h1A705,4);
TASK_PP(16'h1A706,4);
TASK_PP(16'h1A707,4);
TASK_PP(16'h1A708,4);
TASK_PP(16'h1A709,4);
TASK_PP(16'h1A70A,4);
TASK_PP(16'h1A70B,4);
TASK_PP(16'h1A70C,4);
TASK_PP(16'h1A70D,4);
TASK_PP(16'h1A70E,4);
TASK_PP(16'h1A70F,4);
TASK_PP(16'h1A710,4);
TASK_PP(16'h1A711,4);
TASK_PP(16'h1A712,4);
TASK_PP(16'h1A713,4);
TASK_PP(16'h1A714,4);
TASK_PP(16'h1A715,4);
TASK_PP(16'h1A716,4);
TASK_PP(16'h1A717,4);
TASK_PP(16'h1A718,4);
TASK_PP(16'h1A719,4);
TASK_PP(16'h1A71A,4);
TASK_PP(16'h1A71B,4);
TASK_PP(16'h1A71C,4);
TASK_PP(16'h1A71D,4);
TASK_PP(16'h1A71E,4);
TASK_PP(16'h1A71F,4);
TASK_PP(16'h1A720,4);
TASK_PP(16'h1A721,4);
TASK_PP(16'h1A722,4);
TASK_PP(16'h1A723,4);
TASK_PP(16'h1A724,4);
TASK_PP(16'h1A725,4);
TASK_PP(16'h1A726,4);
TASK_PP(16'h1A727,4);
TASK_PP(16'h1A728,4);
TASK_PP(16'h1A729,4);
TASK_PP(16'h1A72A,4);
TASK_PP(16'h1A72B,4);
TASK_PP(16'h1A72C,4);
TASK_PP(16'h1A72D,4);
TASK_PP(16'h1A72E,4);
TASK_PP(16'h1A72F,4);
TASK_PP(16'h1A730,4);
TASK_PP(16'h1A731,4);
TASK_PP(16'h1A732,4);
TASK_PP(16'h1A733,4);
TASK_PP(16'h1A734,4);
TASK_PP(16'h1A735,4);
TASK_PP(16'h1A736,4);
TASK_PP(16'h1A737,4);
TASK_PP(16'h1A738,4);
TASK_PP(16'h1A739,4);
TASK_PP(16'h1A73A,4);
TASK_PP(16'h1A73B,4);
TASK_PP(16'h1A73C,4);
TASK_PP(16'h1A73D,4);
TASK_PP(16'h1A73E,4);
TASK_PP(16'h1A73F,4);
TASK_PP(16'h1A740,4);
TASK_PP(16'h1A741,4);
TASK_PP(16'h1A742,4);
TASK_PP(16'h1A743,4);
TASK_PP(16'h1A744,4);
TASK_PP(16'h1A745,4);
TASK_PP(16'h1A746,4);
TASK_PP(16'h1A747,4);
TASK_PP(16'h1A748,4);
TASK_PP(16'h1A749,4);
TASK_PP(16'h1A74A,4);
TASK_PP(16'h1A74B,4);
TASK_PP(16'h1A74C,4);
TASK_PP(16'h1A74D,4);
TASK_PP(16'h1A74E,4);
TASK_PP(16'h1A74F,4);
TASK_PP(16'h1A750,4);
TASK_PP(16'h1A751,4);
TASK_PP(16'h1A752,4);
TASK_PP(16'h1A753,4);
TASK_PP(16'h1A754,4);
TASK_PP(16'h1A755,4);
TASK_PP(16'h1A756,4);
TASK_PP(16'h1A757,4);
TASK_PP(16'h1A758,4);
TASK_PP(16'h1A759,4);
TASK_PP(16'h1A75A,4);
TASK_PP(16'h1A75B,4);
TASK_PP(16'h1A75C,4);
TASK_PP(16'h1A75D,4);
TASK_PP(16'h1A75E,4);
TASK_PP(16'h1A75F,4);
TASK_PP(16'h1A760,4);
TASK_PP(16'h1A761,4);
TASK_PP(16'h1A762,4);
TASK_PP(16'h1A763,4);
TASK_PP(16'h1A764,4);
TASK_PP(16'h1A765,4);
TASK_PP(16'h1A766,4);
TASK_PP(16'h1A767,4);
TASK_PP(16'h1A768,4);
TASK_PP(16'h1A769,4);
TASK_PP(16'h1A76A,4);
TASK_PP(16'h1A76B,4);
TASK_PP(16'h1A76C,4);
TASK_PP(16'h1A76D,4);
TASK_PP(16'h1A76E,4);
TASK_PP(16'h1A76F,4);
TASK_PP(16'h1A770,4);
TASK_PP(16'h1A771,4);
TASK_PP(16'h1A772,4);
TASK_PP(16'h1A773,4);
TASK_PP(16'h1A774,4);
TASK_PP(16'h1A775,4);
TASK_PP(16'h1A776,4);
TASK_PP(16'h1A777,4);
TASK_PP(16'h1A778,4);
TASK_PP(16'h1A779,4);
TASK_PP(16'h1A77A,4);
TASK_PP(16'h1A77B,4);
TASK_PP(16'h1A77C,4);
TASK_PP(16'h1A77D,4);
TASK_PP(16'h1A77E,4);
TASK_PP(16'h1A77F,4);
TASK_PP(16'h1A780,4);
TASK_PP(16'h1A781,4);
TASK_PP(16'h1A782,4);
TASK_PP(16'h1A783,4);
TASK_PP(16'h1A784,4);
TASK_PP(16'h1A785,4);
TASK_PP(16'h1A786,4);
TASK_PP(16'h1A787,4);
TASK_PP(16'h1A788,4);
TASK_PP(16'h1A789,4);
TASK_PP(16'h1A78A,4);
TASK_PP(16'h1A78B,4);
TASK_PP(16'h1A78C,4);
TASK_PP(16'h1A78D,4);
TASK_PP(16'h1A78E,4);
TASK_PP(16'h1A78F,4);
TASK_PP(16'h1A790,4);
TASK_PP(16'h1A791,4);
TASK_PP(16'h1A792,4);
TASK_PP(16'h1A793,4);
TASK_PP(16'h1A794,4);
TASK_PP(16'h1A795,4);
TASK_PP(16'h1A796,4);
TASK_PP(16'h1A797,4);
TASK_PP(16'h1A798,4);
TASK_PP(16'h1A799,4);
TASK_PP(16'h1A79A,4);
TASK_PP(16'h1A79B,4);
TASK_PP(16'h1A79C,4);
TASK_PP(16'h1A79D,4);
TASK_PP(16'h1A79E,4);
TASK_PP(16'h1A79F,4);
TASK_PP(16'h1A7A0,4);
TASK_PP(16'h1A7A1,4);
TASK_PP(16'h1A7A2,4);
TASK_PP(16'h1A7A3,4);
TASK_PP(16'h1A7A4,4);
TASK_PP(16'h1A7A5,4);
TASK_PP(16'h1A7A6,4);
TASK_PP(16'h1A7A7,4);
TASK_PP(16'h1A7A8,4);
TASK_PP(16'h1A7A9,4);
TASK_PP(16'h1A7AA,4);
TASK_PP(16'h1A7AB,4);
TASK_PP(16'h1A7AC,4);
TASK_PP(16'h1A7AD,4);
TASK_PP(16'h1A7AE,4);
TASK_PP(16'h1A7AF,4);
TASK_PP(16'h1A7B0,4);
TASK_PP(16'h1A7B1,4);
TASK_PP(16'h1A7B2,4);
TASK_PP(16'h1A7B3,4);
TASK_PP(16'h1A7B4,4);
TASK_PP(16'h1A7B5,4);
TASK_PP(16'h1A7B6,4);
TASK_PP(16'h1A7B7,4);
TASK_PP(16'h1A7B8,4);
TASK_PP(16'h1A7B9,4);
TASK_PP(16'h1A7BA,4);
TASK_PP(16'h1A7BB,4);
TASK_PP(16'h1A7BC,4);
TASK_PP(16'h1A7BD,4);
TASK_PP(16'h1A7BE,4);
TASK_PP(16'h1A7BF,4);
TASK_PP(16'h1A7C0,4);
TASK_PP(16'h1A7C1,4);
TASK_PP(16'h1A7C2,4);
TASK_PP(16'h1A7C3,4);
TASK_PP(16'h1A7C4,4);
TASK_PP(16'h1A7C5,4);
TASK_PP(16'h1A7C6,4);
TASK_PP(16'h1A7C7,4);
TASK_PP(16'h1A7C8,4);
TASK_PP(16'h1A7C9,4);
TASK_PP(16'h1A7CA,4);
TASK_PP(16'h1A7CB,4);
TASK_PP(16'h1A7CC,4);
TASK_PP(16'h1A7CD,4);
TASK_PP(16'h1A7CE,4);
TASK_PP(16'h1A7CF,4);
TASK_PP(16'h1A7D0,4);
TASK_PP(16'h1A7D1,4);
TASK_PP(16'h1A7D2,4);
TASK_PP(16'h1A7D3,4);
TASK_PP(16'h1A7D4,4);
TASK_PP(16'h1A7D5,4);
TASK_PP(16'h1A7D6,4);
TASK_PP(16'h1A7D7,4);
TASK_PP(16'h1A7D8,4);
TASK_PP(16'h1A7D9,4);
TASK_PP(16'h1A7DA,4);
TASK_PP(16'h1A7DB,4);
TASK_PP(16'h1A7DC,4);
TASK_PP(16'h1A7DD,4);
TASK_PP(16'h1A7DE,4);
TASK_PP(16'h1A7DF,4);
TASK_PP(16'h1A7E0,4);
TASK_PP(16'h1A7E1,4);
TASK_PP(16'h1A7E2,4);
TASK_PP(16'h1A7E3,4);
TASK_PP(16'h1A7E4,4);
TASK_PP(16'h1A7E5,4);
TASK_PP(16'h1A7E6,4);
TASK_PP(16'h1A7E7,4);
TASK_PP(16'h1A7E8,4);
TASK_PP(16'h1A7E9,4);
TASK_PP(16'h1A7EA,4);
TASK_PP(16'h1A7EB,4);
TASK_PP(16'h1A7EC,4);
TASK_PP(16'h1A7ED,4);
TASK_PP(16'h1A7EE,4);
TASK_PP(16'h1A7EF,4);
TASK_PP(16'h1A7F0,4);
TASK_PP(16'h1A7F1,4);
TASK_PP(16'h1A7F2,4);
TASK_PP(16'h1A7F3,4);
TASK_PP(16'h1A7F4,4);
TASK_PP(16'h1A7F5,4);
TASK_PP(16'h1A7F6,4);
TASK_PP(16'h1A7F7,4);
TASK_PP(16'h1A7F8,4);
TASK_PP(16'h1A7F9,4);
TASK_PP(16'h1A7FA,4);
TASK_PP(16'h1A7FB,4);
TASK_PP(16'h1A7FC,4);
TASK_PP(16'h1A7FD,4);
TASK_PP(16'h1A7FE,4);
TASK_PP(16'h1A7FF,4);
TASK_PP(16'h1A800,4);
TASK_PP(16'h1A801,4);
TASK_PP(16'h1A802,4);
TASK_PP(16'h1A803,4);
TASK_PP(16'h1A804,4);
TASK_PP(16'h1A805,4);
TASK_PP(16'h1A806,4);
TASK_PP(16'h1A807,4);
TASK_PP(16'h1A808,4);
TASK_PP(16'h1A809,4);
TASK_PP(16'h1A80A,4);
TASK_PP(16'h1A80B,4);
TASK_PP(16'h1A80C,4);
TASK_PP(16'h1A80D,4);
TASK_PP(16'h1A80E,4);
TASK_PP(16'h1A80F,4);
TASK_PP(16'h1A810,4);
TASK_PP(16'h1A811,4);
TASK_PP(16'h1A812,4);
TASK_PP(16'h1A813,4);
TASK_PP(16'h1A814,4);
TASK_PP(16'h1A815,4);
TASK_PP(16'h1A816,4);
TASK_PP(16'h1A817,4);
TASK_PP(16'h1A818,4);
TASK_PP(16'h1A819,4);
TASK_PP(16'h1A81A,4);
TASK_PP(16'h1A81B,4);
TASK_PP(16'h1A81C,4);
TASK_PP(16'h1A81D,4);
TASK_PP(16'h1A81E,4);
TASK_PP(16'h1A81F,4);
TASK_PP(16'h1A820,4);
TASK_PP(16'h1A821,4);
TASK_PP(16'h1A822,4);
TASK_PP(16'h1A823,4);
TASK_PP(16'h1A824,4);
TASK_PP(16'h1A825,4);
TASK_PP(16'h1A826,4);
TASK_PP(16'h1A827,4);
TASK_PP(16'h1A828,4);
TASK_PP(16'h1A829,4);
TASK_PP(16'h1A82A,4);
TASK_PP(16'h1A82B,4);
TASK_PP(16'h1A82C,4);
TASK_PP(16'h1A82D,4);
TASK_PP(16'h1A82E,4);
TASK_PP(16'h1A82F,4);
TASK_PP(16'h1A830,4);
TASK_PP(16'h1A831,4);
TASK_PP(16'h1A832,4);
TASK_PP(16'h1A833,4);
TASK_PP(16'h1A834,4);
TASK_PP(16'h1A835,4);
TASK_PP(16'h1A836,4);
TASK_PP(16'h1A837,4);
TASK_PP(16'h1A838,4);
TASK_PP(16'h1A839,4);
TASK_PP(16'h1A83A,4);
TASK_PP(16'h1A83B,4);
TASK_PP(16'h1A83C,4);
TASK_PP(16'h1A83D,4);
TASK_PP(16'h1A83E,4);
TASK_PP(16'h1A83F,4);
TASK_PP(16'h1A840,4);
TASK_PP(16'h1A841,4);
TASK_PP(16'h1A842,4);
TASK_PP(16'h1A843,4);
TASK_PP(16'h1A844,4);
TASK_PP(16'h1A845,4);
TASK_PP(16'h1A846,4);
TASK_PP(16'h1A847,4);
TASK_PP(16'h1A848,4);
TASK_PP(16'h1A849,4);
TASK_PP(16'h1A84A,4);
TASK_PP(16'h1A84B,4);
TASK_PP(16'h1A84C,4);
TASK_PP(16'h1A84D,4);
TASK_PP(16'h1A84E,4);
TASK_PP(16'h1A84F,4);
TASK_PP(16'h1A850,4);
TASK_PP(16'h1A851,4);
TASK_PP(16'h1A852,4);
TASK_PP(16'h1A853,4);
TASK_PP(16'h1A854,4);
TASK_PP(16'h1A855,4);
TASK_PP(16'h1A856,4);
TASK_PP(16'h1A857,4);
TASK_PP(16'h1A858,4);
TASK_PP(16'h1A859,4);
TASK_PP(16'h1A85A,4);
TASK_PP(16'h1A85B,4);
TASK_PP(16'h1A85C,4);
TASK_PP(16'h1A85D,4);
TASK_PP(16'h1A85E,4);
TASK_PP(16'h1A85F,4);
TASK_PP(16'h1A860,4);
TASK_PP(16'h1A861,4);
TASK_PP(16'h1A862,4);
TASK_PP(16'h1A863,4);
TASK_PP(16'h1A864,4);
TASK_PP(16'h1A865,4);
TASK_PP(16'h1A866,4);
TASK_PP(16'h1A867,4);
TASK_PP(16'h1A868,4);
TASK_PP(16'h1A869,4);
TASK_PP(16'h1A86A,4);
TASK_PP(16'h1A86B,4);
TASK_PP(16'h1A86C,4);
TASK_PP(16'h1A86D,4);
TASK_PP(16'h1A86E,4);
TASK_PP(16'h1A86F,4);
TASK_PP(16'h1A870,4);
TASK_PP(16'h1A871,4);
TASK_PP(16'h1A872,4);
TASK_PP(16'h1A873,4);
TASK_PP(16'h1A874,4);
TASK_PP(16'h1A875,4);
TASK_PP(16'h1A876,4);
TASK_PP(16'h1A877,4);
TASK_PP(16'h1A878,4);
TASK_PP(16'h1A879,4);
TASK_PP(16'h1A87A,4);
TASK_PP(16'h1A87B,4);
TASK_PP(16'h1A87C,4);
TASK_PP(16'h1A87D,4);
TASK_PP(16'h1A87E,4);
TASK_PP(16'h1A87F,4);
TASK_PP(16'h1A880,4);
TASK_PP(16'h1A881,4);
TASK_PP(16'h1A882,4);
TASK_PP(16'h1A883,4);
TASK_PP(16'h1A884,4);
TASK_PP(16'h1A885,4);
TASK_PP(16'h1A886,4);
TASK_PP(16'h1A887,4);
TASK_PP(16'h1A888,4);
TASK_PP(16'h1A889,4);
TASK_PP(16'h1A88A,4);
TASK_PP(16'h1A88B,4);
TASK_PP(16'h1A88C,4);
TASK_PP(16'h1A88D,4);
TASK_PP(16'h1A88E,4);
TASK_PP(16'h1A88F,4);
TASK_PP(16'h1A890,4);
TASK_PP(16'h1A891,4);
TASK_PP(16'h1A892,4);
TASK_PP(16'h1A893,4);
TASK_PP(16'h1A894,4);
TASK_PP(16'h1A895,4);
TASK_PP(16'h1A896,4);
TASK_PP(16'h1A897,4);
TASK_PP(16'h1A898,4);
TASK_PP(16'h1A899,4);
TASK_PP(16'h1A89A,4);
TASK_PP(16'h1A89B,4);
TASK_PP(16'h1A89C,4);
TASK_PP(16'h1A89D,4);
TASK_PP(16'h1A89E,4);
TASK_PP(16'h1A89F,4);
TASK_PP(16'h1A8A0,4);
TASK_PP(16'h1A8A1,4);
TASK_PP(16'h1A8A2,4);
TASK_PP(16'h1A8A3,4);
TASK_PP(16'h1A8A4,4);
TASK_PP(16'h1A8A5,4);
TASK_PP(16'h1A8A6,4);
TASK_PP(16'h1A8A7,4);
TASK_PP(16'h1A8A8,4);
TASK_PP(16'h1A8A9,4);
TASK_PP(16'h1A8AA,4);
TASK_PP(16'h1A8AB,4);
TASK_PP(16'h1A8AC,4);
TASK_PP(16'h1A8AD,4);
TASK_PP(16'h1A8AE,4);
TASK_PP(16'h1A8AF,4);
TASK_PP(16'h1A8B0,4);
TASK_PP(16'h1A8B1,4);
TASK_PP(16'h1A8B2,4);
TASK_PP(16'h1A8B3,4);
TASK_PP(16'h1A8B4,4);
TASK_PP(16'h1A8B5,4);
TASK_PP(16'h1A8B6,4);
TASK_PP(16'h1A8B7,4);
TASK_PP(16'h1A8B8,4);
TASK_PP(16'h1A8B9,4);
TASK_PP(16'h1A8BA,4);
TASK_PP(16'h1A8BB,4);
TASK_PP(16'h1A8BC,4);
TASK_PP(16'h1A8BD,4);
TASK_PP(16'h1A8BE,4);
TASK_PP(16'h1A8BF,4);
TASK_PP(16'h1A8C0,4);
TASK_PP(16'h1A8C1,4);
TASK_PP(16'h1A8C2,4);
TASK_PP(16'h1A8C3,4);
TASK_PP(16'h1A8C4,4);
TASK_PP(16'h1A8C5,4);
TASK_PP(16'h1A8C6,4);
TASK_PP(16'h1A8C7,4);
TASK_PP(16'h1A8C8,4);
TASK_PP(16'h1A8C9,4);
TASK_PP(16'h1A8CA,4);
TASK_PP(16'h1A8CB,4);
TASK_PP(16'h1A8CC,4);
TASK_PP(16'h1A8CD,4);
TASK_PP(16'h1A8CE,4);
TASK_PP(16'h1A8CF,4);
TASK_PP(16'h1A8D0,4);
TASK_PP(16'h1A8D1,4);
TASK_PP(16'h1A8D2,4);
TASK_PP(16'h1A8D3,4);
TASK_PP(16'h1A8D4,4);
TASK_PP(16'h1A8D5,4);
TASK_PP(16'h1A8D6,4);
TASK_PP(16'h1A8D7,4);
TASK_PP(16'h1A8D8,4);
TASK_PP(16'h1A8D9,4);
TASK_PP(16'h1A8DA,4);
TASK_PP(16'h1A8DB,4);
TASK_PP(16'h1A8DC,4);
TASK_PP(16'h1A8DD,4);
TASK_PP(16'h1A8DE,4);
TASK_PP(16'h1A8DF,4);
TASK_PP(16'h1A8E0,4);
TASK_PP(16'h1A8E1,4);
TASK_PP(16'h1A8E2,4);
TASK_PP(16'h1A8E3,4);
TASK_PP(16'h1A8E4,4);
TASK_PP(16'h1A8E5,4);
TASK_PP(16'h1A8E6,4);
TASK_PP(16'h1A8E7,4);
TASK_PP(16'h1A8E8,4);
TASK_PP(16'h1A8E9,4);
TASK_PP(16'h1A8EA,4);
TASK_PP(16'h1A8EB,4);
TASK_PP(16'h1A8EC,4);
TASK_PP(16'h1A8ED,4);
TASK_PP(16'h1A8EE,4);
TASK_PP(16'h1A8EF,4);
TASK_PP(16'h1A8F0,4);
TASK_PP(16'h1A8F1,4);
TASK_PP(16'h1A8F2,4);
TASK_PP(16'h1A8F3,4);
TASK_PP(16'h1A8F4,4);
TASK_PP(16'h1A8F5,4);
TASK_PP(16'h1A8F6,4);
TASK_PP(16'h1A8F7,4);
TASK_PP(16'h1A8F8,4);
TASK_PP(16'h1A8F9,4);
TASK_PP(16'h1A8FA,4);
TASK_PP(16'h1A8FB,4);
TASK_PP(16'h1A8FC,4);
TASK_PP(16'h1A8FD,4);
TASK_PP(16'h1A8FE,4);
TASK_PP(16'h1A8FF,4);
TASK_PP(16'h1A900,4);
TASK_PP(16'h1A901,4);
TASK_PP(16'h1A902,4);
TASK_PP(16'h1A903,4);
TASK_PP(16'h1A904,4);
TASK_PP(16'h1A905,4);
TASK_PP(16'h1A906,4);
TASK_PP(16'h1A907,4);
TASK_PP(16'h1A908,4);
TASK_PP(16'h1A909,4);
TASK_PP(16'h1A90A,4);
TASK_PP(16'h1A90B,4);
TASK_PP(16'h1A90C,4);
TASK_PP(16'h1A90D,4);
TASK_PP(16'h1A90E,4);
TASK_PP(16'h1A90F,4);
TASK_PP(16'h1A910,4);
TASK_PP(16'h1A911,4);
TASK_PP(16'h1A912,4);
TASK_PP(16'h1A913,4);
TASK_PP(16'h1A914,4);
TASK_PP(16'h1A915,4);
TASK_PP(16'h1A916,4);
TASK_PP(16'h1A917,4);
TASK_PP(16'h1A918,4);
TASK_PP(16'h1A919,4);
TASK_PP(16'h1A91A,4);
TASK_PP(16'h1A91B,4);
TASK_PP(16'h1A91C,4);
TASK_PP(16'h1A91D,4);
TASK_PP(16'h1A91E,4);
TASK_PP(16'h1A91F,4);
TASK_PP(16'h1A920,4);
TASK_PP(16'h1A921,4);
TASK_PP(16'h1A922,4);
TASK_PP(16'h1A923,4);
TASK_PP(16'h1A924,4);
TASK_PP(16'h1A925,4);
TASK_PP(16'h1A926,4);
TASK_PP(16'h1A927,4);
TASK_PP(16'h1A928,4);
TASK_PP(16'h1A929,4);
TASK_PP(16'h1A92A,4);
TASK_PP(16'h1A92B,4);
TASK_PP(16'h1A92C,4);
TASK_PP(16'h1A92D,4);
TASK_PP(16'h1A92E,4);
TASK_PP(16'h1A92F,4);
TASK_PP(16'h1A930,4);
TASK_PP(16'h1A931,4);
TASK_PP(16'h1A932,4);
TASK_PP(16'h1A933,4);
TASK_PP(16'h1A934,4);
TASK_PP(16'h1A935,4);
TASK_PP(16'h1A936,4);
TASK_PP(16'h1A937,4);
TASK_PP(16'h1A938,4);
TASK_PP(16'h1A939,4);
TASK_PP(16'h1A93A,4);
TASK_PP(16'h1A93B,4);
TASK_PP(16'h1A93C,4);
TASK_PP(16'h1A93D,4);
TASK_PP(16'h1A93E,4);
TASK_PP(16'h1A93F,4);
TASK_PP(16'h1A940,4);
TASK_PP(16'h1A941,4);
TASK_PP(16'h1A942,4);
TASK_PP(16'h1A943,4);
TASK_PP(16'h1A944,4);
TASK_PP(16'h1A945,4);
TASK_PP(16'h1A946,4);
TASK_PP(16'h1A947,4);
TASK_PP(16'h1A948,4);
TASK_PP(16'h1A949,4);
TASK_PP(16'h1A94A,4);
TASK_PP(16'h1A94B,4);
TASK_PP(16'h1A94C,4);
TASK_PP(16'h1A94D,4);
TASK_PP(16'h1A94E,4);
TASK_PP(16'h1A94F,4);
TASK_PP(16'h1A950,4);
TASK_PP(16'h1A951,4);
TASK_PP(16'h1A952,4);
TASK_PP(16'h1A953,4);
TASK_PP(16'h1A954,4);
TASK_PP(16'h1A955,4);
TASK_PP(16'h1A956,4);
TASK_PP(16'h1A957,4);
TASK_PP(16'h1A958,4);
TASK_PP(16'h1A959,4);
TASK_PP(16'h1A95A,4);
TASK_PP(16'h1A95B,4);
TASK_PP(16'h1A95C,4);
TASK_PP(16'h1A95D,4);
TASK_PP(16'h1A95E,4);
TASK_PP(16'h1A95F,4);
TASK_PP(16'h1A960,4);
TASK_PP(16'h1A961,4);
TASK_PP(16'h1A962,4);
TASK_PP(16'h1A963,4);
TASK_PP(16'h1A964,4);
TASK_PP(16'h1A965,4);
TASK_PP(16'h1A966,4);
TASK_PP(16'h1A967,4);
TASK_PP(16'h1A968,4);
TASK_PP(16'h1A969,4);
TASK_PP(16'h1A96A,4);
TASK_PP(16'h1A96B,4);
TASK_PP(16'h1A96C,4);
TASK_PP(16'h1A96D,4);
TASK_PP(16'h1A96E,4);
TASK_PP(16'h1A96F,4);
TASK_PP(16'h1A970,4);
TASK_PP(16'h1A971,4);
TASK_PP(16'h1A972,4);
TASK_PP(16'h1A973,4);
TASK_PP(16'h1A974,4);
TASK_PP(16'h1A975,4);
TASK_PP(16'h1A976,4);
TASK_PP(16'h1A977,4);
TASK_PP(16'h1A978,4);
TASK_PP(16'h1A979,4);
TASK_PP(16'h1A97A,4);
TASK_PP(16'h1A97B,4);
TASK_PP(16'h1A97C,4);
TASK_PP(16'h1A97D,4);
TASK_PP(16'h1A97E,4);
TASK_PP(16'h1A97F,4);
TASK_PP(16'h1A980,4);
TASK_PP(16'h1A981,4);
TASK_PP(16'h1A982,4);
TASK_PP(16'h1A983,4);
TASK_PP(16'h1A984,4);
TASK_PP(16'h1A985,4);
TASK_PP(16'h1A986,4);
TASK_PP(16'h1A987,4);
TASK_PP(16'h1A988,4);
TASK_PP(16'h1A989,4);
TASK_PP(16'h1A98A,4);
TASK_PP(16'h1A98B,4);
TASK_PP(16'h1A98C,4);
TASK_PP(16'h1A98D,4);
TASK_PP(16'h1A98E,4);
TASK_PP(16'h1A98F,4);
TASK_PP(16'h1A990,4);
TASK_PP(16'h1A991,4);
TASK_PP(16'h1A992,4);
TASK_PP(16'h1A993,4);
TASK_PP(16'h1A994,4);
TASK_PP(16'h1A995,4);
TASK_PP(16'h1A996,4);
TASK_PP(16'h1A997,4);
TASK_PP(16'h1A998,4);
TASK_PP(16'h1A999,4);
TASK_PP(16'h1A99A,4);
TASK_PP(16'h1A99B,4);
TASK_PP(16'h1A99C,4);
TASK_PP(16'h1A99D,4);
TASK_PP(16'h1A99E,4);
TASK_PP(16'h1A99F,4);
TASK_PP(16'h1A9A0,4);
TASK_PP(16'h1A9A1,4);
TASK_PP(16'h1A9A2,4);
TASK_PP(16'h1A9A3,4);
TASK_PP(16'h1A9A4,4);
TASK_PP(16'h1A9A5,4);
TASK_PP(16'h1A9A6,4);
TASK_PP(16'h1A9A7,4);
TASK_PP(16'h1A9A8,4);
TASK_PP(16'h1A9A9,4);
TASK_PP(16'h1A9AA,4);
TASK_PP(16'h1A9AB,4);
TASK_PP(16'h1A9AC,4);
TASK_PP(16'h1A9AD,4);
TASK_PP(16'h1A9AE,4);
TASK_PP(16'h1A9AF,4);
TASK_PP(16'h1A9B0,4);
TASK_PP(16'h1A9B1,4);
TASK_PP(16'h1A9B2,4);
TASK_PP(16'h1A9B3,4);
TASK_PP(16'h1A9B4,4);
TASK_PP(16'h1A9B5,4);
TASK_PP(16'h1A9B6,4);
TASK_PP(16'h1A9B7,4);
TASK_PP(16'h1A9B8,4);
TASK_PP(16'h1A9B9,4);
TASK_PP(16'h1A9BA,4);
TASK_PP(16'h1A9BB,4);
TASK_PP(16'h1A9BC,4);
TASK_PP(16'h1A9BD,4);
TASK_PP(16'h1A9BE,4);
TASK_PP(16'h1A9BF,4);
TASK_PP(16'h1A9C0,4);
TASK_PP(16'h1A9C1,4);
TASK_PP(16'h1A9C2,4);
TASK_PP(16'h1A9C3,4);
TASK_PP(16'h1A9C4,4);
TASK_PP(16'h1A9C5,4);
TASK_PP(16'h1A9C6,4);
TASK_PP(16'h1A9C7,4);
TASK_PP(16'h1A9C8,4);
TASK_PP(16'h1A9C9,4);
TASK_PP(16'h1A9CA,4);
TASK_PP(16'h1A9CB,4);
TASK_PP(16'h1A9CC,4);
TASK_PP(16'h1A9CD,4);
TASK_PP(16'h1A9CE,4);
TASK_PP(16'h1A9CF,4);
TASK_PP(16'h1A9D0,4);
TASK_PP(16'h1A9D1,4);
TASK_PP(16'h1A9D2,4);
TASK_PP(16'h1A9D3,4);
TASK_PP(16'h1A9D4,4);
TASK_PP(16'h1A9D5,4);
TASK_PP(16'h1A9D6,4);
TASK_PP(16'h1A9D7,4);
TASK_PP(16'h1A9D8,4);
TASK_PP(16'h1A9D9,4);
TASK_PP(16'h1A9DA,4);
TASK_PP(16'h1A9DB,4);
TASK_PP(16'h1A9DC,4);
TASK_PP(16'h1A9DD,4);
TASK_PP(16'h1A9DE,4);
TASK_PP(16'h1A9DF,4);
TASK_PP(16'h1A9E0,4);
TASK_PP(16'h1A9E1,4);
TASK_PP(16'h1A9E2,4);
TASK_PP(16'h1A9E3,4);
TASK_PP(16'h1A9E4,4);
TASK_PP(16'h1A9E5,4);
TASK_PP(16'h1A9E6,4);
TASK_PP(16'h1A9E7,4);
TASK_PP(16'h1A9E8,4);
TASK_PP(16'h1A9E9,4);
TASK_PP(16'h1A9EA,4);
TASK_PP(16'h1A9EB,4);
TASK_PP(16'h1A9EC,4);
TASK_PP(16'h1A9ED,4);
TASK_PP(16'h1A9EE,4);
TASK_PP(16'h1A9EF,4);
TASK_PP(16'h1A9F0,4);
TASK_PP(16'h1A9F1,4);
TASK_PP(16'h1A9F2,4);
TASK_PP(16'h1A9F3,4);
TASK_PP(16'h1A9F4,4);
TASK_PP(16'h1A9F5,4);
TASK_PP(16'h1A9F6,4);
TASK_PP(16'h1A9F7,4);
TASK_PP(16'h1A9F8,4);
TASK_PP(16'h1A9F9,4);
TASK_PP(16'h1A9FA,4);
TASK_PP(16'h1A9FB,4);
TASK_PP(16'h1A9FC,4);
TASK_PP(16'h1A9FD,4);
TASK_PP(16'h1A9FE,4);
TASK_PP(16'h1A9FF,4);
TASK_PP(16'h1AA00,4);
TASK_PP(16'h1AA01,4);
TASK_PP(16'h1AA02,4);
TASK_PP(16'h1AA03,4);
TASK_PP(16'h1AA04,4);
TASK_PP(16'h1AA05,4);
TASK_PP(16'h1AA06,4);
TASK_PP(16'h1AA07,4);
TASK_PP(16'h1AA08,4);
TASK_PP(16'h1AA09,4);
TASK_PP(16'h1AA0A,4);
TASK_PP(16'h1AA0B,4);
TASK_PP(16'h1AA0C,4);
TASK_PP(16'h1AA0D,4);
TASK_PP(16'h1AA0E,4);
TASK_PP(16'h1AA0F,4);
TASK_PP(16'h1AA10,4);
TASK_PP(16'h1AA11,4);
TASK_PP(16'h1AA12,4);
TASK_PP(16'h1AA13,4);
TASK_PP(16'h1AA14,4);
TASK_PP(16'h1AA15,4);
TASK_PP(16'h1AA16,4);
TASK_PP(16'h1AA17,4);
TASK_PP(16'h1AA18,4);
TASK_PP(16'h1AA19,4);
TASK_PP(16'h1AA1A,4);
TASK_PP(16'h1AA1B,4);
TASK_PP(16'h1AA1C,4);
TASK_PP(16'h1AA1D,4);
TASK_PP(16'h1AA1E,4);
TASK_PP(16'h1AA1F,4);
TASK_PP(16'h1AA20,4);
TASK_PP(16'h1AA21,4);
TASK_PP(16'h1AA22,4);
TASK_PP(16'h1AA23,4);
TASK_PP(16'h1AA24,4);
TASK_PP(16'h1AA25,4);
TASK_PP(16'h1AA26,4);
TASK_PP(16'h1AA27,4);
TASK_PP(16'h1AA28,4);
TASK_PP(16'h1AA29,4);
TASK_PP(16'h1AA2A,4);
TASK_PP(16'h1AA2B,4);
TASK_PP(16'h1AA2C,4);
TASK_PP(16'h1AA2D,4);
TASK_PP(16'h1AA2E,4);
TASK_PP(16'h1AA2F,4);
TASK_PP(16'h1AA30,4);
TASK_PP(16'h1AA31,4);
TASK_PP(16'h1AA32,4);
TASK_PP(16'h1AA33,4);
TASK_PP(16'h1AA34,4);
TASK_PP(16'h1AA35,4);
TASK_PP(16'h1AA36,4);
TASK_PP(16'h1AA37,4);
TASK_PP(16'h1AA38,4);
TASK_PP(16'h1AA39,4);
TASK_PP(16'h1AA3A,4);
TASK_PP(16'h1AA3B,4);
TASK_PP(16'h1AA3C,4);
TASK_PP(16'h1AA3D,4);
TASK_PP(16'h1AA3E,4);
TASK_PP(16'h1AA3F,4);
TASK_PP(16'h1AA40,4);
TASK_PP(16'h1AA41,4);
TASK_PP(16'h1AA42,4);
TASK_PP(16'h1AA43,4);
TASK_PP(16'h1AA44,4);
TASK_PP(16'h1AA45,4);
TASK_PP(16'h1AA46,4);
TASK_PP(16'h1AA47,4);
TASK_PP(16'h1AA48,4);
TASK_PP(16'h1AA49,4);
TASK_PP(16'h1AA4A,4);
TASK_PP(16'h1AA4B,4);
TASK_PP(16'h1AA4C,4);
TASK_PP(16'h1AA4D,4);
TASK_PP(16'h1AA4E,4);
TASK_PP(16'h1AA4F,4);
TASK_PP(16'h1AA50,4);
TASK_PP(16'h1AA51,4);
TASK_PP(16'h1AA52,4);
TASK_PP(16'h1AA53,4);
TASK_PP(16'h1AA54,4);
TASK_PP(16'h1AA55,4);
TASK_PP(16'h1AA56,4);
TASK_PP(16'h1AA57,4);
TASK_PP(16'h1AA58,4);
TASK_PP(16'h1AA59,4);
TASK_PP(16'h1AA5A,4);
TASK_PP(16'h1AA5B,4);
TASK_PP(16'h1AA5C,4);
TASK_PP(16'h1AA5D,4);
TASK_PP(16'h1AA5E,4);
TASK_PP(16'h1AA5F,4);
TASK_PP(16'h1AA60,4);
TASK_PP(16'h1AA61,4);
TASK_PP(16'h1AA62,4);
TASK_PP(16'h1AA63,4);
TASK_PP(16'h1AA64,4);
TASK_PP(16'h1AA65,4);
TASK_PP(16'h1AA66,4);
TASK_PP(16'h1AA67,4);
TASK_PP(16'h1AA68,4);
TASK_PP(16'h1AA69,4);
TASK_PP(16'h1AA6A,4);
TASK_PP(16'h1AA6B,4);
TASK_PP(16'h1AA6C,4);
TASK_PP(16'h1AA6D,4);
TASK_PP(16'h1AA6E,4);
TASK_PP(16'h1AA6F,4);
TASK_PP(16'h1AA70,4);
TASK_PP(16'h1AA71,4);
TASK_PP(16'h1AA72,4);
TASK_PP(16'h1AA73,4);
TASK_PP(16'h1AA74,4);
TASK_PP(16'h1AA75,4);
TASK_PP(16'h1AA76,4);
TASK_PP(16'h1AA77,4);
TASK_PP(16'h1AA78,4);
TASK_PP(16'h1AA79,4);
TASK_PP(16'h1AA7A,4);
TASK_PP(16'h1AA7B,4);
TASK_PP(16'h1AA7C,4);
TASK_PP(16'h1AA7D,4);
TASK_PP(16'h1AA7E,4);
TASK_PP(16'h1AA7F,4);
TASK_PP(16'h1AA80,4);
TASK_PP(16'h1AA81,4);
TASK_PP(16'h1AA82,4);
TASK_PP(16'h1AA83,4);
TASK_PP(16'h1AA84,4);
TASK_PP(16'h1AA85,4);
TASK_PP(16'h1AA86,4);
TASK_PP(16'h1AA87,4);
TASK_PP(16'h1AA88,4);
TASK_PP(16'h1AA89,4);
TASK_PP(16'h1AA8A,4);
TASK_PP(16'h1AA8B,4);
TASK_PP(16'h1AA8C,4);
TASK_PP(16'h1AA8D,4);
TASK_PP(16'h1AA8E,4);
TASK_PP(16'h1AA8F,4);
TASK_PP(16'h1AA90,4);
TASK_PP(16'h1AA91,4);
TASK_PP(16'h1AA92,4);
TASK_PP(16'h1AA93,4);
TASK_PP(16'h1AA94,4);
TASK_PP(16'h1AA95,4);
TASK_PP(16'h1AA96,4);
TASK_PP(16'h1AA97,4);
TASK_PP(16'h1AA98,4);
TASK_PP(16'h1AA99,4);
TASK_PP(16'h1AA9A,4);
TASK_PP(16'h1AA9B,4);
TASK_PP(16'h1AA9C,4);
TASK_PP(16'h1AA9D,4);
TASK_PP(16'h1AA9E,4);
TASK_PP(16'h1AA9F,4);
TASK_PP(16'h1AAA0,4);
TASK_PP(16'h1AAA1,4);
TASK_PP(16'h1AAA2,4);
TASK_PP(16'h1AAA3,4);
TASK_PP(16'h1AAA4,4);
TASK_PP(16'h1AAA5,4);
TASK_PP(16'h1AAA6,4);
TASK_PP(16'h1AAA7,4);
TASK_PP(16'h1AAA8,4);
TASK_PP(16'h1AAA9,4);
TASK_PP(16'h1AAAA,4);
TASK_PP(16'h1AAAB,4);
TASK_PP(16'h1AAAC,4);
TASK_PP(16'h1AAAD,4);
TASK_PP(16'h1AAAE,4);
TASK_PP(16'h1AAAF,4);
TASK_PP(16'h1AAB0,4);
TASK_PP(16'h1AAB1,4);
TASK_PP(16'h1AAB2,4);
TASK_PP(16'h1AAB3,4);
TASK_PP(16'h1AAB4,4);
TASK_PP(16'h1AAB5,4);
TASK_PP(16'h1AAB6,4);
TASK_PP(16'h1AAB7,4);
TASK_PP(16'h1AAB8,4);
TASK_PP(16'h1AAB9,4);
TASK_PP(16'h1AABA,4);
TASK_PP(16'h1AABB,4);
TASK_PP(16'h1AABC,4);
TASK_PP(16'h1AABD,4);
TASK_PP(16'h1AABE,4);
TASK_PP(16'h1AABF,4);
TASK_PP(16'h1AAC0,4);
TASK_PP(16'h1AAC1,4);
TASK_PP(16'h1AAC2,4);
TASK_PP(16'h1AAC3,4);
TASK_PP(16'h1AAC4,4);
TASK_PP(16'h1AAC5,4);
TASK_PP(16'h1AAC6,4);
TASK_PP(16'h1AAC7,4);
TASK_PP(16'h1AAC8,4);
TASK_PP(16'h1AAC9,4);
TASK_PP(16'h1AACA,4);
TASK_PP(16'h1AACB,4);
TASK_PP(16'h1AACC,4);
TASK_PP(16'h1AACD,4);
TASK_PP(16'h1AACE,4);
TASK_PP(16'h1AACF,4);
TASK_PP(16'h1AAD0,4);
TASK_PP(16'h1AAD1,4);
TASK_PP(16'h1AAD2,4);
TASK_PP(16'h1AAD3,4);
TASK_PP(16'h1AAD4,4);
TASK_PP(16'h1AAD5,4);
TASK_PP(16'h1AAD6,4);
TASK_PP(16'h1AAD7,4);
TASK_PP(16'h1AAD8,4);
TASK_PP(16'h1AAD9,4);
TASK_PP(16'h1AADA,4);
TASK_PP(16'h1AADB,4);
TASK_PP(16'h1AADC,4);
TASK_PP(16'h1AADD,4);
TASK_PP(16'h1AADE,4);
TASK_PP(16'h1AADF,4);
TASK_PP(16'h1AAE0,4);
TASK_PP(16'h1AAE1,4);
TASK_PP(16'h1AAE2,4);
TASK_PP(16'h1AAE3,4);
TASK_PP(16'h1AAE4,4);
TASK_PP(16'h1AAE5,4);
TASK_PP(16'h1AAE6,4);
TASK_PP(16'h1AAE7,4);
TASK_PP(16'h1AAE8,4);
TASK_PP(16'h1AAE9,4);
TASK_PP(16'h1AAEA,4);
TASK_PP(16'h1AAEB,4);
TASK_PP(16'h1AAEC,4);
TASK_PP(16'h1AAED,4);
TASK_PP(16'h1AAEE,4);
TASK_PP(16'h1AAEF,4);
TASK_PP(16'h1AAF0,4);
TASK_PP(16'h1AAF1,4);
TASK_PP(16'h1AAF2,4);
TASK_PP(16'h1AAF3,4);
TASK_PP(16'h1AAF4,4);
TASK_PP(16'h1AAF5,4);
TASK_PP(16'h1AAF6,4);
TASK_PP(16'h1AAF7,4);
TASK_PP(16'h1AAF8,4);
TASK_PP(16'h1AAF9,4);
TASK_PP(16'h1AAFA,4);
TASK_PP(16'h1AAFB,4);
TASK_PP(16'h1AAFC,4);
TASK_PP(16'h1AAFD,4);
TASK_PP(16'h1AAFE,4);
TASK_PP(16'h1AAFF,4);
TASK_PP(16'h1AB00,4);
TASK_PP(16'h1AB01,4);
TASK_PP(16'h1AB02,4);
TASK_PP(16'h1AB03,4);
TASK_PP(16'h1AB04,4);
TASK_PP(16'h1AB05,4);
TASK_PP(16'h1AB06,4);
TASK_PP(16'h1AB07,4);
TASK_PP(16'h1AB08,4);
TASK_PP(16'h1AB09,4);
TASK_PP(16'h1AB0A,4);
TASK_PP(16'h1AB0B,4);
TASK_PP(16'h1AB0C,4);
TASK_PP(16'h1AB0D,4);
TASK_PP(16'h1AB0E,4);
TASK_PP(16'h1AB0F,4);
TASK_PP(16'h1AB10,4);
TASK_PP(16'h1AB11,4);
TASK_PP(16'h1AB12,4);
TASK_PP(16'h1AB13,4);
TASK_PP(16'h1AB14,4);
TASK_PP(16'h1AB15,4);
TASK_PP(16'h1AB16,4);
TASK_PP(16'h1AB17,4);
TASK_PP(16'h1AB18,4);
TASK_PP(16'h1AB19,4);
TASK_PP(16'h1AB1A,4);
TASK_PP(16'h1AB1B,4);
TASK_PP(16'h1AB1C,4);
TASK_PP(16'h1AB1D,4);
TASK_PP(16'h1AB1E,4);
TASK_PP(16'h1AB1F,4);
TASK_PP(16'h1AB20,4);
TASK_PP(16'h1AB21,4);
TASK_PP(16'h1AB22,4);
TASK_PP(16'h1AB23,4);
TASK_PP(16'h1AB24,4);
TASK_PP(16'h1AB25,4);
TASK_PP(16'h1AB26,4);
TASK_PP(16'h1AB27,4);
TASK_PP(16'h1AB28,4);
TASK_PP(16'h1AB29,4);
TASK_PP(16'h1AB2A,4);
TASK_PP(16'h1AB2B,4);
TASK_PP(16'h1AB2C,4);
TASK_PP(16'h1AB2D,4);
TASK_PP(16'h1AB2E,4);
TASK_PP(16'h1AB2F,4);
TASK_PP(16'h1AB30,4);
TASK_PP(16'h1AB31,4);
TASK_PP(16'h1AB32,4);
TASK_PP(16'h1AB33,4);
TASK_PP(16'h1AB34,4);
TASK_PP(16'h1AB35,4);
TASK_PP(16'h1AB36,4);
TASK_PP(16'h1AB37,4);
TASK_PP(16'h1AB38,4);
TASK_PP(16'h1AB39,4);
TASK_PP(16'h1AB3A,4);
TASK_PP(16'h1AB3B,4);
TASK_PP(16'h1AB3C,4);
TASK_PP(16'h1AB3D,4);
TASK_PP(16'h1AB3E,4);
TASK_PP(16'h1AB3F,4);
TASK_PP(16'h1AB40,4);
TASK_PP(16'h1AB41,4);
TASK_PP(16'h1AB42,4);
TASK_PP(16'h1AB43,4);
TASK_PP(16'h1AB44,4);
TASK_PP(16'h1AB45,4);
TASK_PP(16'h1AB46,4);
TASK_PP(16'h1AB47,4);
TASK_PP(16'h1AB48,4);
TASK_PP(16'h1AB49,4);
TASK_PP(16'h1AB4A,4);
TASK_PP(16'h1AB4B,4);
TASK_PP(16'h1AB4C,4);
TASK_PP(16'h1AB4D,4);
TASK_PP(16'h1AB4E,4);
TASK_PP(16'h1AB4F,4);
TASK_PP(16'h1AB50,4);
TASK_PP(16'h1AB51,4);
TASK_PP(16'h1AB52,4);
TASK_PP(16'h1AB53,4);
TASK_PP(16'h1AB54,4);
TASK_PP(16'h1AB55,4);
TASK_PP(16'h1AB56,4);
TASK_PP(16'h1AB57,4);
TASK_PP(16'h1AB58,4);
TASK_PP(16'h1AB59,4);
TASK_PP(16'h1AB5A,4);
TASK_PP(16'h1AB5B,4);
TASK_PP(16'h1AB5C,4);
TASK_PP(16'h1AB5D,4);
TASK_PP(16'h1AB5E,4);
TASK_PP(16'h1AB5F,4);
TASK_PP(16'h1AB60,4);
TASK_PP(16'h1AB61,4);
TASK_PP(16'h1AB62,4);
TASK_PP(16'h1AB63,4);
TASK_PP(16'h1AB64,4);
TASK_PP(16'h1AB65,4);
TASK_PP(16'h1AB66,4);
TASK_PP(16'h1AB67,4);
TASK_PP(16'h1AB68,4);
TASK_PP(16'h1AB69,4);
TASK_PP(16'h1AB6A,4);
TASK_PP(16'h1AB6B,4);
TASK_PP(16'h1AB6C,4);
TASK_PP(16'h1AB6D,4);
TASK_PP(16'h1AB6E,4);
TASK_PP(16'h1AB6F,4);
TASK_PP(16'h1AB70,4);
TASK_PP(16'h1AB71,4);
TASK_PP(16'h1AB72,4);
TASK_PP(16'h1AB73,4);
TASK_PP(16'h1AB74,4);
TASK_PP(16'h1AB75,4);
TASK_PP(16'h1AB76,4);
TASK_PP(16'h1AB77,4);
TASK_PP(16'h1AB78,4);
TASK_PP(16'h1AB79,4);
TASK_PP(16'h1AB7A,4);
TASK_PP(16'h1AB7B,4);
TASK_PP(16'h1AB7C,4);
TASK_PP(16'h1AB7D,4);
TASK_PP(16'h1AB7E,4);
TASK_PP(16'h1AB7F,4);
TASK_PP(16'h1AB80,4);
TASK_PP(16'h1AB81,4);
TASK_PP(16'h1AB82,4);
TASK_PP(16'h1AB83,4);
TASK_PP(16'h1AB84,4);
TASK_PP(16'h1AB85,4);
TASK_PP(16'h1AB86,4);
TASK_PP(16'h1AB87,4);
TASK_PP(16'h1AB88,4);
TASK_PP(16'h1AB89,4);
TASK_PP(16'h1AB8A,4);
TASK_PP(16'h1AB8B,4);
TASK_PP(16'h1AB8C,4);
TASK_PP(16'h1AB8D,4);
TASK_PP(16'h1AB8E,4);
TASK_PP(16'h1AB8F,4);
TASK_PP(16'h1AB90,4);
TASK_PP(16'h1AB91,4);
TASK_PP(16'h1AB92,4);
TASK_PP(16'h1AB93,4);
TASK_PP(16'h1AB94,4);
TASK_PP(16'h1AB95,4);
TASK_PP(16'h1AB96,4);
TASK_PP(16'h1AB97,4);
TASK_PP(16'h1AB98,4);
TASK_PP(16'h1AB99,4);
TASK_PP(16'h1AB9A,4);
TASK_PP(16'h1AB9B,4);
TASK_PP(16'h1AB9C,4);
TASK_PP(16'h1AB9D,4);
TASK_PP(16'h1AB9E,4);
TASK_PP(16'h1AB9F,4);
TASK_PP(16'h1ABA0,4);
TASK_PP(16'h1ABA1,4);
TASK_PP(16'h1ABA2,4);
TASK_PP(16'h1ABA3,4);
TASK_PP(16'h1ABA4,4);
TASK_PP(16'h1ABA5,4);
TASK_PP(16'h1ABA6,4);
TASK_PP(16'h1ABA7,4);
TASK_PP(16'h1ABA8,4);
TASK_PP(16'h1ABA9,4);
TASK_PP(16'h1ABAA,4);
TASK_PP(16'h1ABAB,4);
TASK_PP(16'h1ABAC,4);
TASK_PP(16'h1ABAD,4);
TASK_PP(16'h1ABAE,4);
TASK_PP(16'h1ABAF,4);
TASK_PP(16'h1ABB0,4);
TASK_PP(16'h1ABB1,4);
TASK_PP(16'h1ABB2,4);
TASK_PP(16'h1ABB3,4);
TASK_PP(16'h1ABB4,4);
TASK_PP(16'h1ABB5,4);
TASK_PP(16'h1ABB6,4);
TASK_PP(16'h1ABB7,4);
TASK_PP(16'h1ABB8,4);
TASK_PP(16'h1ABB9,4);
TASK_PP(16'h1ABBA,4);
TASK_PP(16'h1ABBB,4);
TASK_PP(16'h1ABBC,4);
TASK_PP(16'h1ABBD,4);
TASK_PP(16'h1ABBE,4);
TASK_PP(16'h1ABBF,4);
TASK_PP(16'h1ABC0,4);
TASK_PP(16'h1ABC1,4);
TASK_PP(16'h1ABC2,4);
TASK_PP(16'h1ABC3,4);
TASK_PP(16'h1ABC4,4);
TASK_PP(16'h1ABC5,4);
TASK_PP(16'h1ABC6,4);
TASK_PP(16'h1ABC7,4);
TASK_PP(16'h1ABC8,4);
TASK_PP(16'h1ABC9,4);
TASK_PP(16'h1ABCA,4);
TASK_PP(16'h1ABCB,4);
TASK_PP(16'h1ABCC,4);
TASK_PP(16'h1ABCD,4);
TASK_PP(16'h1ABCE,4);
TASK_PP(16'h1ABCF,4);
TASK_PP(16'h1ABD0,4);
TASK_PP(16'h1ABD1,4);
TASK_PP(16'h1ABD2,4);
TASK_PP(16'h1ABD3,4);
TASK_PP(16'h1ABD4,4);
TASK_PP(16'h1ABD5,4);
TASK_PP(16'h1ABD6,4);
TASK_PP(16'h1ABD7,4);
TASK_PP(16'h1ABD8,4);
TASK_PP(16'h1ABD9,4);
TASK_PP(16'h1ABDA,4);
TASK_PP(16'h1ABDB,4);
TASK_PP(16'h1ABDC,4);
TASK_PP(16'h1ABDD,4);
TASK_PP(16'h1ABDE,4);
TASK_PP(16'h1ABDF,4);
TASK_PP(16'h1ABE0,4);
TASK_PP(16'h1ABE1,4);
TASK_PP(16'h1ABE2,4);
TASK_PP(16'h1ABE3,4);
TASK_PP(16'h1ABE4,4);
TASK_PP(16'h1ABE5,4);
TASK_PP(16'h1ABE6,4);
TASK_PP(16'h1ABE7,4);
TASK_PP(16'h1ABE8,4);
TASK_PP(16'h1ABE9,4);
TASK_PP(16'h1ABEA,4);
TASK_PP(16'h1ABEB,4);
TASK_PP(16'h1ABEC,4);
TASK_PP(16'h1ABED,4);
TASK_PP(16'h1ABEE,4);
TASK_PP(16'h1ABEF,4);
TASK_PP(16'h1ABF0,4);
TASK_PP(16'h1ABF1,4);
TASK_PP(16'h1ABF2,4);
TASK_PP(16'h1ABF3,4);
TASK_PP(16'h1ABF4,4);
TASK_PP(16'h1ABF5,4);
TASK_PP(16'h1ABF6,4);
TASK_PP(16'h1ABF7,4);
TASK_PP(16'h1ABF8,4);
TASK_PP(16'h1ABF9,4);
TASK_PP(16'h1ABFA,4);
TASK_PP(16'h1ABFB,4);
TASK_PP(16'h1ABFC,4);
TASK_PP(16'h1ABFD,4);
TASK_PP(16'h1ABFE,4);
TASK_PP(16'h1ABFF,4);
TASK_PP(16'h1AC00,4);
TASK_PP(16'h1AC01,4);
TASK_PP(16'h1AC02,4);
TASK_PP(16'h1AC03,4);
TASK_PP(16'h1AC04,4);
TASK_PP(16'h1AC05,4);
TASK_PP(16'h1AC06,4);
TASK_PP(16'h1AC07,4);
TASK_PP(16'h1AC08,4);
TASK_PP(16'h1AC09,4);
TASK_PP(16'h1AC0A,4);
TASK_PP(16'h1AC0B,4);
TASK_PP(16'h1AC0C,4);
TASK_PP(16'h1AC0D,4);
TASK_PP(16'h1AC0E,4);
TASK_PP(16'h1AC0F,4);
TASK_PP(16'h1AC10,4);
TASK_PP(16'h1AC11,4);
TASK_PP(16'h1AC12,4);
TASK_PP(16'h1AC13,4);
TASK_PP(16'h1AC14,4);
TASK_PP(16'h1AC15,4);
TASK_PP(16'h1AC16,4);
TASK_PP(16'h1AC17,4);
TASK_PP(16'h1AC18,4);
TASK_PP(16'h1AC19,4);
TASK_PP(16'h1AC1A,4);
TASK_PP(16'h1AC1B,4);
TASK_PP(16'h1AC1C,4);
TASK_PP(16'h1AC1D,4);
TASK_PP(16'h1AC1E,4);
TASK_PP(16'h1AC1F,4);
TASK_PP(16'h1AC20,4);
TASK_PP(16'h1AC21,4);
TASK_PP(16'h1AC22,4);
TASK_PP(16'h1AC23,4);
TASK_PP(16'h1AC24,4);
TASK_PP(16'h1AC25,4);
TASK_PP(16'h1AC26,4);
TASK_PP(16'h1AC27,4);
TASK_PP(16'h1AC28,4);
TASK_PP(16'h1AC29,4);
TASK_PP(16'h1AC2A,4);
TASK_PP(16'h1AC2B,4);
TASK_PP(16'h1AC2C,4);
TASK_PP(16'h1AC2D,4);
TASK_PP(16'h1AC2E,4);
TASK_PP(16'h1AC2F,4);
TASK_PP(16'h1AC30,4);
TASK_PP(16'h1AC31,4);
TASK_PP(16'h1AC32,4);
TASK_PP(16'h1AC33,4);
TASK_PP(16'h1AC34,4);
TASK_PP(16'h1AC35,4);
TASK_PP(16'h1AC36,4);
TASK_PP(16'h1AC37,4);
TASK_PP(16'h1AC38,4);
TASK_PP(16'h1AC39,4);
TASK_PP(16'h1AC3A,4);
TASK_PP(16'h1AC3B,4);
TASK_PP(16'h1AC3C,4);
TASK_PP(16'h1AC3D,4);
TASK_PP(16'h1AC3E,4);
TASK_PP(16'h1AC3F,4);
TASK_PP(16'h1AC40,4);
TASK_PP(16'h1AC41,4);
TASK_PP(16'h1AC42,4);
TASK_PP(16'h1AC43,4);
TASK_PP(16'h1AC44,4);
TASK_PP(16'h1AC45,4);
TASK_PP(16'h1AC46,4);
TASK_PP(16'h1AC47,4);
TASK_PP(16'h1AC48,4);
TASK_PP(16'h1AC49,4);
TASK_PP(16'h1AC4A,4);
TASK_PP(16'h1AC4B,4);
TASK_PP(16'h1AC4C,4);
TASK_PP(16'h1AC4D,4);
TASK_PP(16'h1AC4E,4);
TASK_PP(16'h1AC4F,4);
TASK_PP(16'h1AC50,4);
TASK_PP(16'h1AC51,4);
TASK_PP(16'h1AC52,4);
TASK_PP(16'h1AC53,4);
TASK_PP(16'h1AC54,4);
TASK_PP(16'h1AC55,4);
TASK_PP(16'h1AC56,4);
TASK_PP(16'h1AC57,4);
TASK_PP(16'h1AC58,4);
TASK_PP(16'h1AC59,4);
TASK_PP(16'h1AC5A,4);
TASK_PP(16'h1AC5B,4);
TASK_PP(16'h1AC5C,4);
TASK_PP(16'h1AC5D,4);
TASK_PP(16'h1AC5E,4);
TASK_PP(16'h1AC5F,4);
TASK_PP(16'h1AC60,4);
TASK_PP(16'h1AC61,4);
TASK_PP(16'h1AC62,4);
TASK_PP(16'h1AC63,4);
TASK_PP(16'h1AC64,4);
TASK_PP(16'h1AC65,4);
TASK_PP(16'h1AC66,4);
TASK_PP(16'h1AC67,4);
TASK_PP(16'h1AC68,4);
TASK_PP(16'h1AC69,4);
TASK_PP(16'h1AC6A,4);
TASK_PP(16'h1AC6B,4);
TASK_PP(16'h1AC6C,4);
TASK_PP(16'h1AC6D,4);
TASK_PP(16'h1AC6E,4);
TASK_PP(16'h1AC6F,4);
TASK_PP(16'h1AC70,4);
TASK_PP(16'h1AC71,4);
TASK_PP(16'h1AC72,4);
TASK_PP(16'h1AC73,4);
TASK_PP(16'h1AC74,4);
TASK_PP(16'h1AC75,4);
TASK_PP(16'h1AC76,4);
TASK_PP(16'h1AC77,4);
TASK_PP(16'h1AC78,4);
TASK_PP(16'h1AC79,4);
TASK_PP(16'h1AC7A,4);
TASK_PP(16'h1AC7B,4);
TASK_PP(16'h1AC7C,4);
TASK_PP(16'h1AC7D,4);
TASK_PP(16'h1AC7E,4);
TASK_PP(16'h1AC7F,4);
TASK_PP(16'h1AC80,4);
TASK_PP(16'h1AC81,4);
TASK_PP(16'h1AC82,4);
TASK_PP(16'h1AC83,4);
TASK_PP(16'h1AC84,4);
TASK_PP(16'h1AC85,4);
TASK_PP(16'h1AC86,4);
TASK_PP(16'h1AC87,4);
TASK_PP(16'h1AC88,4);
TASK_PP(16'h1AC89,4);
TASK_PP(16'h1AC8A,4);
TASK_PP(16'h1AC8B,4);
TASK_PP(16'h1AC8C,4);
TASK_PP(16'h1AC8D,4);
TASK_PP(16'h1AC8E,4);
TASK_PP(16'h1AC8F,4);
TASK_PP(16'h1AC90,4);
TASK_PP(16'h1AC91,4);
TASK_PP(16'h1AC92,4);
TASK_PP(16'h1AC93,4);
TASK_PP(16'h1AC94,4);
TASK_PP(16'h1AC95,4);
TASK_PP(16'h1AC96,4);
TASK_PP(16'h1AC97,4);
TASK_PP(16'h1AC98,4);
TASK_PP(16'h1AC99,4);
TASK_PP(16'h1AC9A,4);
TASK_PP(16'h1AC9B,4);
TASK_PP(16'h1AC9C,4);
TASK_PP(16'h1AC9D,4);
TASK_PP(16'h1AC9E,4);
TASK_PP(16'h1AC9F,4);
TASK_PP(16'h1ACA0,4);
TASK_PP(16'h1ACA1,4);
TASK_PP(16'h1ACA2,4);
TASK_PP(16'h1ACA3,4);
TASK_PP(16'h1ACA4,4);
TASK_PP(16'h1ACA5,4);
TASK_PP(16'h1ACA6,4);
TASK_PP(16'h1ACA7,4);
TASK_PP(16'h1ACA8,4);
TASK_PP(16'h1ACA9,4);
TASK_PP(16'h1ACAA,4);
TASK_PP(16'h1ACAB,4);
TASK_PP(16'h1ACAC,4);
TASK_PP(16'h1ACAD,4);
TASK_PP(16'h1ACAE,4);
TASK_PP(16'h1ACAF,4);
TASK_PP(16'h1ACB0,4);
TASK_PP(16'h1ACB1,4);
TASK_PP(16'h1ACB2,4);
TASK_PP(16'h1ACB3,4);
TASK_PP(16'h1ACB4,4);
TASK_PP(16'h1ACB5,4);
TASK_PP(16'h1ACB6,4);
TASK_PP(16'h1ACB7,4);
TASK_PP(16'h1ACB8,4);
TASK_PP(16'h1ACB9,4);
TASK_PP(16'h1ACBA,4);
TASK_PP(16'h1ACBB,4);
TASK_PP(16'h1ACBC,4);
TASK_PP(16'h1ACBD,4);
TASK_PP(16'h1ACBE,4);
TASK_PP(16'h1ACBF,4);
TASK_PP(16'h1ACC0,4);
TASK_PP(16'h1ACC1,4);
TASK_PP(16'h1ACC2,4);
TASK_PP(16'h1ACC3,4);
TASK_PP(16'h1ACC4,4);
TASK_PP(16'h1ACC5,4);
TASK_PP(16'h1ACC6,4);
TASK_PP(16'h1ACC7,4);
TASK_PP(16'h1ACC8,4);
TASK_PP(16'h1ACC9,4);
TASK_PP(16'h1ACCA,4);
TASK_PP(16'h1ACCB,4);
TASK_PP(16'h1ACCC,4);
TASK_PP(16'h1ACCD,4);
TASK_PP(16'h1ACCE,4);
TASK_PP(16'h1ACCF,4);
TASK_PP(16'h1ACD0,4);
TASK_PP(16'h1ACD1,4);
TASK_PP(16'h1ACD2,4);
TASK_PP(16'h1ACD3,4);
TASK_PP(16'h1ACD4,4);
TASK_PP(16'h1ACD5,4);
TASK_PP(16'h1ACD6,4);
TASK_PP(16'h1ACD7,4);
TASK_PP(16'h1ACD8,4);
TASK_PP(16'h1ACD9,4);
TASK_PP(16'h1ACDA,4);
TASK_PP(16'h1ACDB,4);
TASK_PP(16'h1ACDC,4);
TASK_PP(16'h1ACDD,4);
TASK_PP(16'h1ACDE,4);
TASK_PP(16'h1ACDF,4);
TASK_PP(16'h1ACE0,4);
TASK_PP(16'h1ACE1,4);
TASK_PP(16'h1ACE2,4);
TASK_PP(16'h1ACE3,4);
TASK_PP(16'h1ACE4,4);
TASK_PP(16'h1ACE5,4);
TASK_PP(16'h1ACE6,4);
TASK_PP(16'h1ACE7,4);
TASK_PP(16'h1ACE8,4);
TASK_PP(16'h1ACE9,4);
TASK_PP(16'h1ACEA,4);
TASK_PP(16'h1ACEB,4);
TASK_PP(16'h1ACEC,4);
TASK_PP(16'h1ACED,4);
TASK_PP(16'h1ACEE,4);
TASK_PP(16'h1ACEF,4);
TASK_PP(16'h1ACF0,4);
TASK_PP(16'h1ACF1,4);
TASK_PP(16'h1ACF2,4);
TASK_PP(16'h1ACF3,4);
TASK_PP(16'h1ACF4,4);
TASK_PP(16'h1ACF5,4);
TASK_PP(16'h1ACF6,4);
TASK_PP(16'h1ACF7,4);
TASK_PP(16'h1ACF8,4);
TASK_PP(16'h1ACF9,4);
TASK_PP(16'h1ACFA,4);
TASK_PP(16'h1ACFB,4);
TASK_PP(16'h1ACFC,4);
TASK_PP(16'h1ACFD,4);
TASK_PP(16'h1ACFE,4);
TASK_PP(16'h1ACFF,4);
TASK_PP(16'h1AD00,4);
TASK_PP(16'h1AD01,4);
TASK_PP(16'h1AD02,4);
TASK_PP(16'h1AD03,4);
TASK_PP(16'h1AD04,4);
TASK_PP(16'h1AD05,4);
TASK_PP(16'h1AD06,4);
TASK_PP(16'h1AD07,4);
TASK_PP(16'h1AD08,4);
TASK_PP(16'h1AD09,4);
TASK_PP(16'h1AD0A,4);
TASK_PP(16'h1AD0B,4);
TASK_PP(16'h1AD0C,4);
TASK_PP(16'h1AD0D,4);
TASK_PP(16'h1AD0E,4);
TASK_PP(16'h1AD0F,4);
TASK_PP(16'h1AD10,4);
TASK_PP(16'h1AD11,4);
TASK_PP(16'h1AD12,4);
TASK_PP(16'h1AD13,4);
TASK_PP(16'h1AD14,4);
TASK_PP(16'h1AD15,4);
TASK_PP(16'h1AD16,4);
TASK_PP(16'h1AD17,4);
TASK_PP(16'h1AD18,4);
TASK_PP(16'h1AD19,4);
TASK_PP(16'h1AD1A,4);
TASK_PP(16'h1AD1B,4);
TASK_PP(16'h1AD1C,4);
TASK_PP(16'h1AD1D,4);
TASK_PP(16'h1AD1E,4);
TASK_PP(16'h1AD1F,4);
TASK_PP(16'h1AD20,4);
TASK_PP(16'h1AD21,4);
TASK_PP(16'h1AD22,4);
TASK_PP(16'h1AD23,4);
TASK_PP(16'h1AD24,4);
TASK_PP(16'h1AD25,4);
TASK_PP(16'h1AD26,4);
TASK_PP(16'h1AD27,4);
TASK_PP(16'h1AD28,4);
TASK_PP(16'h1AD29,4);
TASK_PP(16'h1AD2A,4);
TASK_PP(16'h1AD2B,4);
TASK_PP(16'h1AD2C,4);
TASK_PP(16'h1AD2D,4);
TASK_PP(16'h1AD2E,4);
TASK_PP(16'h1AD2F,4);
TASK_PP(16'h1AD30,4);
TASK_PP(16'h1AD31,4);
TASK_PP(16'h1AD32,4);
TASK_PP(16'h1AD33,4);
TASK_PP(16'h1AD34,4);
TASK_PP(16'h1AD35,4);
TASK_PP(16'h1AD36,4);
TASK_PP(16'h1AD37,4);
TASK_PP(16'h1AD38,4);
TASK_PP(16'h1AD39,4);
TASK_PP(16'h1AD3A,4);
TASK_PP(16'h1AD3B,4);
TASK_PP(16'h1AD3C,4);
TASK_PP(16'h1AD3D,4);
TASK_PP(16'h1AD3E,4);
TASK_PP(16'h1AD3F,4);
TASK_PP(16'h1AD40,4);
TASK_PP(16'h1AD41,4);
TASK_PP(16'h1AD42,4);
TASK_PP(16'h1AD43,4);
TASK_PP(16'h1AD44,4);
TASK_PP(16'h1AD45,4);
TASK_PP(16'h1AD46,4);
TASK_PP(16'h1AD47,4);
TASK_PP(16'h1AD48,4);
TASK_PP(16'h1AD49,4);
TASK_PP(16'h1AD4A,4);
TASK_PP(16'h1AD4B,4);
TASK_PP(16'h1AD4C,4);
TASK_PP(16'h1AD4D,4);
TASK_PP(16'h1AD4E,4);
TASK_PP(16'h1AD4F,4);
TASK_PP(16'h1AD50,4);
TASK_PP(16'h1AD51,4);
TASK_PP(16'h1AD52,4);
TASK_PP(16'h1AD53,4);
TASK_PP(16'h1AD54,4);
TASK_PP(16'h1AD55,4);
TASK_PP(16'h1AD56,4);
TASK_PP(16'h1AD57,4);
TASK_PP(16'h1AD58,4);
TASK_PP(16'h1AD59,4);
TASK_PP(16'h1AD5A,4);
TASK_PP(16'h1AD5B,4);
TASK_PP(16'h1AD5C,4);
TASK_PP(16'h1AD5D,4);
TASK_PP(16'h1AD5E,4);
TASK_PP(16'h1AD5F,4);
TASK_PP(16'h1AD60,4);
TASK_PP(16'h1AD61,4);
TASK_PP(16'h1AD62,4);
TASK_PP(16'h1AD63,4);
TASK_PP(16'h1AD64,4);
TASK_PP(16'h1AD65,4);
TASK_PP(16'h1AD66,4);
TASK_PP(16'h1AD67,4);
TASK_PP(16'h1AD68,4);
TASK_PP(16'h1AD69,4);
TASK_PP(16'h1AD6A,4);
TASK_PP(16'h1AD6B,4);
TASK_PP(16'h1AD6C,4);
TASK_PP(16'h1AD6D,4);
TASK_PP(16'h1AD6E,4);
TASK_PP(16'h1AD6F,4);
TASK_PP(16'h1AD70,4);
TASK_PP(16'h1AD71,4);
TASK_PP(16'h1AD72,4);
TASK_PP(16'h1AD73,4);
TASK_PP(16'h1AD74,4);
TASK_PP(16'h1AD75,4);
TASK_PP(16'h1AD76,4);
TASK_PP(16'h1AD77,4);
TASK_PP(16'h1AD78,4);
TASK_PP(16'h1AD79,4);
TASK_PP(16'h1AD7A,4);
TASK_PP(16'h1AD7B,4);
TASK_PP(16'h1AD7C,4);
TASK_PP(16'h1AD7D,4);
TASK_PP(16'h1AD7E,4);
TASK_PP(16'h1AD7F,4);
TASK_PP(16'h1AD80,4);
TASK_PP(16'h1AD81,4);
TASK_PP(16'h1AD82,4);
TASK_PP(16'h1AD83,4);
TASK_PP(16'h1AD84,4);
TASK_PP(16'h1AD85,4);
TASK_PP(16'h1AD86,4);
TASK_PP(16'h1AD87,4);
TASK_PP(16'h1AD88,4);
TASK_PP(16'h1AD89,4);
TASK_PP(16'h1AD8A,4);
TASK_PP(16'h1AD8B,4);
TASK_PP(16'h1AD8C,4);
TASK_PP(16'h1AD8D,4);
TASK_PP(16'h1AD8E,4);
TASK_PP(16'h1AD8F,4);
TASK_PP(16'h1AD90,4);
TASK_PP(16'h1AD91,4);
TASK_PP(16'h1AD92,4);
TASK_PP(16'h1AD93,4);
TASK_PP(16'h1AD94,4);
TASK_PP(16'h1AD95,4);
TASK_PP(16'h1AD96,4);
TASK_PP(16'h1AD97,4);
TASK_PP(16'h1AD98,4);
TASK_PP(16'h1AD99,4);
TASK_PP(16'h1AD9A,4);
TASK_PP(16'h1AD9B,4);
TASK_PP(16'h1AD9C,4);
TASK_PP(16'h1AD9D,4);
TASK_PP(16'h1AD9E,4);
TASK_PP(16'h1AD9F,4);
TASK_PP(16'h1ADA0,4);
TASK_PP(16'h1ADA1,4);
TASK_PP(16'h1ADA2,4);
TASK_PP(16'h1ADA3,4);
TASK_PP(16'h1ADA4,4);
TASK_PP(16'h1ADA5,4);
TASK_PP(16'h1ADA6,4);
TASK_PP(16'h1ADA7,4);
TASK_PP(16'h1ADA8,4);
TASK_PP(16'h1ADA9,4);
TASK_PP(16'h1ADAA,4);
TASK_PP(16'h1ADAB,4);
TASK_PP(16'h1ADAC,4);
TASK_PP(16'h1ADAD,4);
TASK_PP(16'h1ADAE,4);
TASK_PP(16'h1ADAF,4);
TASK_PP(16'h1ADB0,4);
TASK_PP(16'h1ADB1,4);
TASK_PP(16'h1ADB2,4);
TASK_PP(16'h1ADB3,4);
TASK_PP(16'h1ADB4,4);
TASK_PP(16'h1ADB5,4);
TASK_PP(16'h1ADB6,4);
TASK_PP(16'h1ADB7,4);
TASK_PP(16'h1ADB8,4);
TASK_PP(16'h1ADB9,4);
TASK_PP(16'h1ADBA,4);
TASK_PP(16'h1ADBB,4);
TASK_PP(16'h1ADBC,4);
TASK_PP(16'h1ADBD,4);
TASK_PP(16'h1ADBE,4);
TASK_PP(16'h1ADBF,4);
TASK_PP(16'h1ADC0,4);
TASK_PP(16'h1ADC1,4);
TASK_PP(16'h1ADC2,4);
TASK_PP(16'h1ADC3,4);
TASK_PP(16'h1ADC4,4);
TASK_PP(16'h1ADC5,4);
TASK_PP(16'h1ADC6,4);
TASK_PP(16'h1ADC7,4);
TASK_PP(16'h1ADC8,4);
TASK_PP(16'h1ADC9,4);
TASK_PP(16'h1ADCA,4);
TASK_PP(16'h1ADCB,4);
TASK_PP(16'h1ADCC,4);
TASK_PP(16'h1ADCD,4);
TASK_PP(16'h1ADCE,4);
TASK_PP(16'h1ADCF,4);
TASK_PP(16'h1ADD0,4);
TASK_PP(16'h1ADD1,4);
TASK_PP(16'h1ADD2,4);
TASK_PP(16'h1ADD3,4);
TASK_PP(16'h1ADD4,4);
TASK_PP(16'h1ADD5,4);
TASK_PP(16'h1ADD6,4);
TASK_PP(16'h1ADD7,4);
TASK_PP(16'h1ADD8,4);
TASK_PP(16'h1ADD9,4);
TASK_PP(16'h1ADDA,4);
TASK_PP(16'h1ADDB,4);
TASK_PP(16'h1ADDC,4);
TASK_PP(16'h1ADDD,4);
TASK_PP(16'h1ADDE,4);
TASK_PP(16'h1ADDF,4);
TASK_PP(16'h1ADE0,4);
TASK_PP(16'h1ADE1,4);
TASK_PP(16'h1ADE2,4);
TASK_PP(16'h1ADE3,4);
TASK_PP(16'h1ADE4,4);
TASK_PP(16'h1ADE5,4);
TASK_PP(16'h1ADE6,4);
TASK_PP(16'h1ADE7,4);
TASK_PP(16'h1ADE8,4);
TASK_PP(16'h1ADE9,4);
TASK_PP(16'h1ADEA,4);
TASK_PP(16'h1ADEB,4);
TASK_PP(16'h1ADEC,4);
TASK_PP(16'h1ADED,4);
TASK_PP(16'h1ADEE,4);
TASK_PP(16'h1ADEF,4);
TASK_PP(16'h1ADF0,4);
TASK_PP(16'h1ADF1,4);
TASK_PP(16'h1ADF2,4);
TASK_PP(16'h1ADF3,4);
TASK_PP(16'h1ADF4,4);
TASK_PP(16'h1ADF5,4);
TASK_PP(16'h1ADF6,4);
TASK_PP(16'h1ADF7,4);
TASK_PP(16'h1ADF8,4);
TASK_PP(16'h1ADF9,4);
TASK_PP(16'h1ADFA,4);
TASK_PP(16'h1ADFB,4);
TASK_PP(16'h1ADFC,4);
TASK_PP(16'h1ADFD,4);
TASK_PP(16'h1ADFE,4);
TASK_PP(16'h1ADFF,4);
TASK_PP(16'h1AE00,4);
TASK_PP(16'h1AE01,4);
TASK_PP(16'h1AE02,4);
TASK_PP(16'h1AE03,4);
TASK_PP(16'h1AE04,4);
TASK_PP(16'h1AE05,4);
TASK_PP(16'h1AE06,4);
TASK_PP(16'h1AE07,4);
TASK_PP(16'h1AE08,4);
TASK_PP(16'h1AE09,4);
TASK_PP(16'h1AE0A,4);
TASK_PP(16'h1AE0B,4);
TASK_PP(16'h1AE0C,4);
TASK_PP(16'h1AE0D,4);
TASK_PP(16'h1AE0E,4);
TASK_PP(16'h1AE0F,4);
TASK_PP(16'h1AE10,4);
TASK_PP(16'h1AE11,4);
TASK_PP(16'h1AE12,4);
TASK_PP(16'h1AE13,4);
TASK_PP(16'h1AE14,4);
TASK_PP(16'h1AE15,4);
TASK_PP(16'h1AE16,4);
TASK_PP(16'h1AE17,4);
TASK_PP(16'h1AE18,4);
TASK_PP(16'h1AE19,4);
TASK_PP(16'h1AE1A,4);
TASK_PP(16'h1AE1B,4);
TASK_PP(16'h1AE1C,4);
TASK_PP(16'h1AE1D,4);
TASK_PP(16'h1AE1E,4);
TASK_PP(16'h1AE1F,4);
TASK_PP(16'h1AE20,4);
TASK_PP(16'h1AE21,4);
TASK_PP(16'h1AE22,4);
TASK_PP(16'h1AE23,4);
TASK_PP(16'h1AE24,4);
TASK_PP(16'h1AE25,4);
TASK_PP(16'h1AE26,4);
TASK_PP(16'h1AE27,4);
TASK_PP(16'h1AE28,4);
TASK_PP(16'h1AE29,4);
TASK_PP(16'h1AE2A,4);
TASK_PP(16'h1AE2B,4);
TASK_PP(16'h1AE2C,4);
TASK_PP(16'h1AE2D,4);
TASK_PP(16'h1AE2E,4);
TASK_PP(16'h1AE2F,4);
TASK_PP(16'h1AE30,4);
TASK_PP(16'h1AE31,4);
TASK_PP(16'h1AE32,4);
TASK_PP(16'h1AE33,4);
TASK_PP(16'h1AE34,4);
TASK_PP(16'h1AE35,4);
TASK_PP(16'h1AE36,4);
TASK_PP(16'h1AE37,4);
TASK_PP(16'h1AE38,4);
TASK_PP(16'h1AE39,4);
TASK_PP(16'h1AE3A,4);
TASK_PP(16'h1AE3B,4);
TASK_PP(16'h1AE3C,4);
TASK_PP(16'h1AE3D,4);
TASK_PP(16'h1AE3E,4);
TASK_PP(16'h1AE3F,4);
TASK_PP(16'h1AE40,4);
TASK_PP(16'h1AE41,4);
TASK_PP(16'h1AE42,4);
TASK_PP(16'h1AE43,4);
TASK_PP(16'h1AE44,4);
TASK_PP(16'h1AE45,4);
TASK_PP(16'h1AE46,4);
TASK_PP(16'h1AE47,4);
TASK_PP(16'h1AE48,4);
TASK_PP(16'h1AE49,4);
TASK_PP(16'h1AE4A,4);
TASK_PP(16'h1AE4B,4);
TASK_PP(16'h1AE4C,4);
TASK_PP(16'h1AE4D,4);
TASK_PP(16'h1AE4E,4);
TASK_PP(16'h1AE4F,4);
TASK_PP(16'h1AE50,4);
TASK_PP(16'h1AE51,4);
TASK_PP(16'h1AE52,4);
TASK_PP(16'h1AE53,4);
TASK_PP(16'h1AE54,4);
TASK_PP(16'h1AE55,4);
TASK_PP(16'h1AE56,4);
TASK_PP(16'h1AE57,4);
TASK_PP(16'h1AE58,4);
TASK_PP(16'h1AE59,4);
TASK_PP(16'h1AE5A,4);
TASK_PP(16'h1AE5B,4);
TASK_PP(16'h1AE5C,4);
TASK_PP(16'h1AE5D,4);
TASK_PP(16'h1AE5E,4);
TASK_PP(16'h1AE5F,4);
TASK_PP(16'h1AE60,4);
TASK_PP(16'h1AE61,4);
TASK_PP(16'h1AE62,4);
TASK_PP(16'h1AE63,4);
TASK_PP(16'h1AE64,4);
TASK_PP(16'h1AE65,4);
TASK_PP(16'h1AE66,4);
TASK_PP(16'h1AE67,4);
TASK_PP(16'h1AE68,4);
TASK_PP(16'h1AE69,4);
TASK_PP(16'h1AE6A,4);
TASK_PP(16'h1AE6B,4);
TASK_PP(16'h1AE6C,4);
TASK_PP(16'h1AE6D,4);
TASK_PP(16'h1AE6E,4);
TASK_PP(16'h1AE6F,4);
TASK_PP(16'h1AE70,4);
TASK_PP(16'h1AE71,4);
TASK_PP(16'h1AE72,4);
TASK_PP(16'h1AE73,4);
TASK_PP(16'h1AE74,4);
TASK_PP(16'h1AE75,4);
TASK_PP(16'h1AE76,4);
TASK_PP(16'h1AE77,4);
TASK_PP(16'h1AE78,4);
TASK_PP(16'h1AE79,4);
TASK_PP(16'h1AE7A,4);
TASK_PP(16'h1AE7B,4);
TASK_PP(16'h1AE7C,4);
TASK_PP(16'h1AE7D,4);
TASK_PP(16'h1AE7E,4);
TASK_PP(16'h1AE7F,4);
TASK_PP(16'h1AE80,4);
TASK_PP(16'h1AE81,4);
TASK_PP(16'h1AE82,4);
TASK_PP(16'h1AE83,4);
TASK_PP(16'h1AE84,4);
TASK_PP(16'h1AE85,4);
TASK_PP(16'h1AE86,4);
TASK_PP(16'h1AE87,4);
TASK_PP(16'h1AE88,4);
TASK_PP(16'h1AE89,4);
TASK_PP(16'h1AE8A,4);
TASK_PP(16'h1AE8B,4);
TASK_PP(16'h1AE8C,4);
TASK_PP(16'h1AE8D,4);
TASK_PP(16'h1AE8E,4);
TASK_PP(16'h1AE8F,4);
TASK_PP(16'h1AE90,4);
TASK_PP(16'h1AE91,4);
TASK_PP(16'h1AE92,4);
TASK_PP(16'h1AE93,4);
TASK_PP(16'h1AE94,4);
TASK_PP(16'h1AE95,4);
TASK_PP(16'h1AE96,4);
TASK_PP(16'h1AE97,4);
TASK_PP(16'h1AE98,4);
TASK_PP(16'h1AE99,4);
TASK_PP(16'h1AE9A,4);
TASK_PP(16'h1AE9B,4);
TASK_PP(16'h1AE9C,4);
TASK_PP(16'h1AE9D,4);
TASK_PP(16'h1AE9E,4);
TASK_PP(16'h1AE9F,4);
TASK_PP(16'h1AEA0,4);
TASK_PP(16'h1AEA1,4);
TASK_PP(16'h1AEA2,4);
TASK_PP(16'h1AEA3,4);
TASK_PP(16'h1AEA4,4);
TASK_PP(16'h1AEA5,4);
TASK_PP(16'h1AEA6,4);
TASK_PP(16'h1AEA7,4);
TASK_PP(16'h1AEA8,4);
TASK_PP(16'h1AEA9,4);
TASK_PP(16'h1AEAA,4);
TASK_PP(16'h1AEAB,4);
TASK_PP(16'h1AEAC,4);
TASK_PP(16'h1AEAD,4);
TASK_PP(16'h1AEAE,4);
TASK_PP(16'h1AEAF,4);
TASK_PP(16'h1AEB0,4);
TASK_PP(16'h1AEB1,4);
TASK_PP(16'h1AEB2,4);
TASK_PP(16'h1AEB3,4);
TASK_PP(16'h1AEB4,4);
TASK_PP(16'h1AEB5,4);
TASK_PP(16'h1AEB6,4);
TASK_PP(16'h1AEB7,4);
TASK_PP(16'h1AEB8,4);
TASK_PP(16'h1AEB9,4);
TASK_PP(16'h1AEBA,4);
TASK_PP(16'h1AEBB,4);
TASK_PP(16'h1AEBC,4);
TASK_PP(16'h1AEBD,4);
TASK_PP(16'h1AEBE,4);
TASK_PP(16'h1AEBF,4);
TASK_PP(16'h1AEC0,4);
TASK_PP(16'h1AEC1,4);
TASK_PP(16'h1AEC2,4);
TASK_PP(16'h1AEC3,4);
TASK_PP(16'h1AEC4,4);
TASK_PP(16'h1AEC5,4);
TASK_PP(16'h1AEC6,4);
TASK_PP(16'h1AEC7,4);
TASK_PP(16'h1AEC8,4);
TASK_PP(16'h1AEC9,4);
TASK_PP(16'h1AECA,4);
TASK_PP(16'h1AECB,4);
TASK_PP(16'h1AECC,4);
TASK_PP(16'h1AECD,4);
TASK_PP(16'h1AECE,4);
TASK_PP(16'h1AECF,4);
TASK_PP(16'h1AED0,4);
TASK_PP(16'h1AED1,4);
TASK_PP(16'h1AED2,4);
TASK_PP(16'h1AED3,4);
TASK_PP(16'h1AED4,4);
TASK_PP(16'h1AED5,4);
TASK_PP(16'h1AED6,4);
TASK_PP(16'h1AED7,4);
TASK_PP(16'h1AED8,4);
TASK_PP(16'h1AED9,4);
TASK_PP(16'h1AEDA,4);
TASK_PP(16'h1AEDB,4);
TASK_PP(16'h1AEDC,4);
TASK_PP(16'h1AEDD,4);
TASK_PP(16'h1AEDE,4);
TASK_PP(16'h1AEDF,4);
TASK_PP(16'h1AEE0,4);
TASK_PP(16'h1AEE1,4);
TASK_PP(16'h1AEE2,4);
TASK_PP(16'h1AEE3,4);
TASK_PP(16'h1AEE4,4);
TASK_PP(16'h1AEE5,4);
TASK_PP(16'h1AEE6,4);
TASK_PP(16'h1AEE7,4);
TASK_PP(16'h1AEE8,4);
TASK_PP(16'h1AEE9,4);
TASK_PP(16'h1AEEA,4);
TASK_PP(16'h1AEEB,4);
TASK_PP(16'h1AEEC,4);
TASK_PP(16'h1AEED,4);
TASK_PP(16'h1AEEE,4);
TASK_PP(16'h1AEEF,4);
TASK_PP(16'h1AEF0,4);
TASK_PP(16'h1AEF1,4);
TASK_PP(16'h1AEF2,4);
TASK_PP(16'h1AEF3,4);
TASK_PP(16'h1AEF4,4);
TASK_PP(16'h1AEF5,4);
TASK_PP(16'h1AEF6,4);
TASK_PP(16'h1AEF7,4);
TASK_PP(16'h1AEF8,4);
TASK_PP(16'h1AEF9,4);
TASK_PP(16'h1AEFA,4);
TASK_PP(16'h1AEFB,4);
TASK_PP(16'h1AEFC,4);
TASK_PP(16'h1AEFD,4);
TASK_PP(16'h1AEFE,4);
TASK_PP(16'h1AEFF,4);
TASK_PP(16'h1AF00,4);
TASK_PP(16'h1AF01,4);
TASK_PP(16'h1AF02,4);
TASK_PP(16'h1AF03,4);
TASK_PP(16'h1AF04,4);
TASK_PP(16'h1AF05,4);
TASK_PP(16'h1AF06,4);
TASK_PP(16'h1AF07,4);
TASK_PP(16'h1AF08,4);
TASK_PP(16'h1AF09,4);
TASK_PP(16'h1AF0A,4);
TASK_PP(16'h1AF0B,4);
TASK_PP(16'h1AF0C,4);
TASK_PP(16'h1AF0D,4);
TASK_PP(16'h1AF0E,4);
TASK_PP(16'h1AF0F,4);
TASK_PP(16'h1AF10,4);
TASK_PP(16'h1AF11,4);
TASK_PP(16'h1AF12,4);
TASK_PP(16'h1AF13,4);
TASK_PP(16'h1AF14,4);
TASK_PP(16'h1AF15,4);
TASK_PP(16'h1AF16,4);
TASK_PP(16'h1AF17,4);
TASK_PP(16'h1AF18,4);
TASK_PP(16'h1AF19,4);
TASK_PP(16'h1AF1A,4);
TASK_PP(16'h1AF1B,4);
TASK_PP(16'h1AF1C,4);
TASK_PP(16'h1AF1D,4);
TASK_PP(16'h1AF1E,4);
TASK_PP(16'h1AF1F,4);
TASK_PP(16'h1AF20,4);
TASK_PP(16'h1AF21,4);
TASK_PP(16'h1AF22,4);
TASK_PP(16'h1AF23,4);
TASK_PP(16'h1AF24,4);
TASK_PP(16'h1AF25,4);
TASK_PP(16'h1AF26,4);
TASK_PP(16'h1AF27,4);
TASK_PP(16'h1AF28,4);
TASK_PP(16'h1AF29,4);
TASK_PP(16'h1AF2A,4);
TASK_PP(16'h1AF2B,4);
TASK_PP(16'h1AF2C,4);
TASK_PP(16'h1AF2D,4);
TASK_PP(16'h1AF2E,4);
TASK_PP(16'h1AF2F,4);
TASK_PP(16'h1AF30,4);
TASK_PP(16'h1AF31,4);
TASK_PP(16'h1AF32,4);
TASK_PP(16'h1AF33,4);
TASK_PP(16'h1AF34,4);
TASK_PP(16'h1AF35,4);
TASK_PP(16'h1AF36,4);
TASK_PP(16'h1AF37,4);
TASK_PP(16'h1AF38,4);
TASK_PP(16'h1AF39,4);
TASK_PP(16'h1AF3A,4);
TASK_PP(16'h1AF3B,4);
TASK_PP(16'h1AF3C,4);
TASK_PP(16'h1AF3D,4);
TASK_PP(16'h1AF3E,4);
TASK_PP(16'h1AF3F,4);
TASK_PP(16'h1AF40,4);
TASK_PP(16'h1AF41,4);
TASK_PP(16'h1AF42,4);
TASK_PP(16'h1AF43,4);
TASK_PP(16'h1AF44,4);
TASK_PP(16'h1AF45,4);
TASK_PP(16'h1AF46,4);
TASK_PP(16'h1AF47,4);
TASK_PP(16'h1AF48,4);
TASK_PP(16'h1AF49,4);
TASK_PP(16'h1AF4A,4);
TASK_PP(16'h1AF4B,4);
TASK_PP(16'h1AF4C,4);
TASK_PP(16'h1AF4D,4);
TASK_PP(16'h1AF4E,4);
TASK_PP(16'h1AF4F,4);
TASK_PP(16'h1AF50,4);
TASK_PP(16'h1AF51,4);
TASK_PP(16'h1AF52,4);
TASK_PP(16'h1AF53,4);
TASK_PP(16'h1AF54,4);
TASK_PP(16'h1AF55,4);
TASK_PP(16'h1AF56,4);
TASK_PP(16'h1AF57,4);
TASK_PP(16'h1AF58,4);
TASK_PP(16'h1AF59,4);
TASK_PP(16'h1AF5A,4);
TASK_PP(16'h1AF5B,4);
TASK_PP(16'h1AF5C,4);
TASK_PP(16'h1AF5D,4);
TASK_PP(16'h1AF5E,4);
TASK_PP(16'h1AF5F,4);
TASK_PP(16'h1AF60,4);
TASK_PP(16'h1AF61,4);
TASK_PP(16'h1AF62,4);
TASK_PP(16'h1AF63,4);
TASK_PP(16'h1AF64,4);
TASK_PP(16'h1AF65,4);
TASK_PP(16'h1AF66,4);
TASK_PP(16'h1AF67,4);
TASK_PP(16'h1AF68,4);
TASK_PP(16'h1AF69,4);
TASK_PP(16'h1AF6A,4);
TASK_PP(16'h1AF6B,4);
TASK_PP(16'h1AF6C,4);
TASK_PP(16'h1AF6D,4);
TASK_PP(16'h1AF6E,4);
TASK_PP(16'h1AF6F,4);
TASK_PP(16'h1AF70,4);
TASK_PP(16'h1AF71,4);
TASK_PP(16'h1AF72,4);
TASK_PP(16'h1AF73,4);
TASK_PP(16'h1AF74,4);
TASK_PP(16'h1AF75,4);
TASK_PP(16'h1AF76,4);
TASK_PP(16'h1AF77,4);
TASK_PP(16'h1AF78,4);
TASK_PP(16'h1AF79,4);
TASK_PP(16'h1AF7A,4);
TASK_PP(16'h1AF7B,4);
TASK_PP(16'h1AF7C,4);
TASK_PP(16'h1AF7D,4);
TASK_PP(16'h1AF7E,4);
TASK_PP(16'h1AF7F,4);
TASK_PP(16'h1AF80,4);
TASK_PP(16'h1AF81,4);
TASK_PP(16'h1AF82,4);
TASK_PP(16'h1AF83,4);
TASK_PP(16'h1AF84,4);
TASK_PP(16'h1AF85,4);
TASK_PP(16'h1AF86,4);
TASK_PP(16'h1AF87,4);
TASK_PP(16'h1AF88,4);
TASK_PP(16'h1AF89,4);
TASK_PP(16'h1AF8A,4);
TASK_PP(16'h1AF8B,4);
TASK_PP(16'h1AF8C,4);
TASK_PP(16'h1AF8D,4);
TASK_PP(16'h1AF8E,4);
TASK_PP(16'h1AF8F,4);
TASK_PP(16'h1AF90,4);
TASK_PP(16'h1AF91,4);
TASK_PP(16'h1AF92,4);
TASK_PP(16'h1AF93,4);
TASK_PP(16'h1AF94,4);
TASK_PP(16'h1AF95,4);
TASK_PP(16'h1AF96,4);
TASK_PP(16'h1AF97,4);
TASK_PP(16'h1AF98,4);
TASK_PP(16'h1AF99,4);
TASK_PP(16'h1AF9A,4);
TASK_PP(16'h1AF9B,4);
TASK_PP(16'h1AF9C,4);
TASK_PP(16'h1AF9D,4);
TASK_PP(16'h1AF9E,4);
TASK_PP(16'h1AF9F,4);
TASK_PP(16'h1AFA0,4);
TASK_PP(16'h1AFA1,4);
TASK_PP(16'h1AFA2,4);
TASK_PP(16'h1AFA3,4);
TASK_PP(16'h1AFA4,4);
TASK_PP(16'h1AFA5,4);
TASK_PP(16'h1AFA6,4);
TASK_PP(16'h1AFA7,4);
TASK_PP(16'h1AFA8,4);
TASK_PP(16'h1AFA9,4);
TASK_PP(16'h1AFAA,4);
TASK_PP(16'h1AFAB,4);
TASK_PP(16'h1AFAC,4);
TASK_PP(16'h1AFAD,4);
TASK_PP(16'h1AFAE,4);
TASK_PP(16'h1AFAF,4);
TASK_PP(16'h1AFB0,4);
TASK_PP(16'h1AFB1,4);
TASK_PP(16'h1AFB2,4);
TASK_PP(16'h1AFB3,4);
TASK_PP(16'h1AFB4,4);
TASK_PP(16'h1AFB5,4);
TASK_PP(16'h1AFB6,4);
TASK_PP(16'h1AFB7,4);
TASK_PP(16'h1AFB8,4);
TASK_PP(16'h1AFB9,4);
TASK_PP(16'h1AFBA,4);
TASK_PP(16'h1AFBB,4);
TASK_PP(16'h1AFBC,4);
TASK_PP(16'h1AFBD,4);
TASK_PP(16'h1AFBE,4);
TASK_PP(16'h1AFBF,4);
TASK_PP(16'h1AFC0,4);
TASK_PP(16'h1AFC1,4);
TASK_PP(16'h1AFC2,4);
TASK_PP(16'h1AFC3,4);
TASK_PP(16'h1AFC4,4);
TASK_PP(16'h1AFC5,4);
TASK_PP(16'h1AFC6,4);
TASK_PP(16'h1AFC7,4);
TASK_PP(16'h1AFC8,4);
TASK_PP(16'h1AFC9,4);
TASK_PP(16'h1AFCA,4);
TASK_PP(16'h1AFCB,4);
TASK_PP(16'h1AFCC,4);
TASK_PP(16'h1AFCD,4);
TASK_PP(16'h1AFCE,4);
TASK_PP(16'h1AFCF,4);
TASK_PP(16'h1AFD0,4);
TASK_PP(16'h1AFD1,4);
TASK_PP(16'h1AFD2,4);
TASK_PP(16'h1AFD3,4);
TASK_PP(16'h1AFD4,4);
TASK_PP(16'h1AFD5,4);
TASK_PP(16'h1AFD6,4);
TASK_PP(16'h1AFD7,4);
TASK_PP(16'h1AFD8,4);
TASK_PP(16'h1AFD9,4);
TASK_PP(16'h1AFDA,4);
TASK_PP(16'h1AFDB,4);
TASK_PP(16'h1AFDC,4);
TASK_PP(16'h1AFDD,4);
TASK_PP(16'h1AFDE,4);
TASK_PP(16'h1AFDF,4);
TASK_PP(16'h1AFE0,4);
TASK_PP(16'h1AFE1,4);
TASK_PP(16'h1AFE2,4);
TASK_PP(16'h1AFE3,4);
TASK_PP(16'h1AFE4,4);
TASK_PP(16'h1AFE5,4);
TASK_PP(16'h1AFE6,4);
TASK_PP(16'h1AFE7,4);
TASK_PP(16'h1AFE8,4);
TASK_PP(16'h1AFE9,4);
TASK_PP(16'h1AFEA,4);
TASK_PP(16'h1AFEB,4);
TASK_PP(16'h1AFEC,4);
TASK_PP(16'h1AFED,4);
TASK_PP(16'h1AFEE,4);
TASK_PP(16'h1AFEF,4);
TASK_PP(16'h1AFF0,4);
TASK_PP(16'h1AFF1,4);
TASK_PP(16'h1AFF2,4);
TASK_PP(16'h1AFF3,4);
TASK_PP(16'h1AFF4,4);
TASK_PP(16'h1AFF5,4);
TASK_PP(16'h1AFF6,4);
TASK_PP(16'h1AFF7,4);
TASK_PP(16'h1AFF8,4);
TASK_PP(16'h1AFF9,4);
TASK_PP(16'h1AFFA,4);
TASK_PP(16'h1AFFB,4);
TASK_PP(16'h1AFFC,4);
TASK_PP(16'h1AFFD,4);
TASK_PP(16'h1AFFE,4);
TASK_PP(16'h1AFFF,4);
TASK_PP(16'h1B000,4);
TASK_PP(16'h1B001,4);
TASK_PP(16'h1B002,4);
TASK_PP(16'h1B003,4);
TASK_PP(16'h1B004,4);
TASK_PP(16'h1B005,4);
TASK_PP(16'h1B006,4);
TASK_PP(16'h1B007,4);
TASK_PP(16'h1B008,4);
TASK_PP(16'h1B009,4);
TASK_PP(16'h1B00A,4);
TASK_PP(16'h1B00B,4);
TASK_PP(16'h1B00C,4);
TASK_PP(16'h1B00D,4);
TASK_PP(16'h1B00E,4);
TASK_PP(16'h1B00F,4);
TASK_PP(16'h1B010,4);
TASK_PP(16'h1B011,4);
TASK_PP(16'h1B012,4);
TASK_PP(16'h1B013,4);
TASK_PP(16'h1B014,4);
TASK_PP(16'h1B015,4);
TASK_PP(16'h1B016,4);
TASK_PP(16'h1B017,4);
TASK_PP(16'h1B018,4);
TASK_PP(16'h1B019,4);
TASK_PP(16'h1B01A,4);
TASK_PP(16'h1B01B,4);
TASK_PP(16'h1B01C,4);
TASK_PP(16'h1B01D,4);
TASK_PP(16'h1B01E,4);
TASK_PP(16'h1B01F,4);
TASK_PP(16'h1B020,4);
TASK_PP(16'h1B021,4);
TASK_PP(16'h1B022,4);
TASK_PP(16'h1B023,4);
TASK_PP(16'h1B024,4);
TASK_PP(16'h1B025,4);
TASK_PP(16'h1B026,4);
TASK_PP(16'h1B027,4);
TASK_PP(16'h1B028,4);
TASK_PP(16'h1B029,4);
TASK_PP(16'h1B02A,4);
TASK_PP(16'h1B02B,4);
TASK_PP(16'h1B02C,4);
TASK_PP(16'h1B02D,4);
TASK_PP(16'h1B02E,4);
TASK_PP(16'h1B02F,4);
TASK_PP(16'h1B030,4);
TASK_PP(16'h1B031,4);
TASK_PP(16'h1B032,4);
TASK_PP(16'h1B033,4);
TASK_PP(16'h1B034,4);
TASK_PP(16'h1B035,4);
TASK_PP(16'h1B036,4);
TASK_PP(16'h1B037,4);
TASK_PP(16'h1B038,4);
TASK_PP(16'h1B039,4);
TASK_PP(16'h1B03A,4);
TASK_PP(16'h1B03B,4);
TASK_PP(16'h1B03C,4);
TASK_PP(16'h1B03D,4);
TASK_PP(16'h1B03E,4);
TASK_PP(16'h1B03F,4);
TASK_PP(16'h1B040,4);
TASK_PP(16'h1B041,4);
TASK_PP(16'h1B042,4);
TASK_PP(16'h1B043,4);
TASK_PP(16'h1B044,4);
TASK_PP(16'h1B045,4);
TASK_PP(16'h1B046,4);
TASK_PP(16'h1B047,4);
TASK_PP(16'h1B048,4);
TASK_PP(16'h1B049,4);
TASK_PP(16'h1B04A,4);
TASK_PP(16'h1B04B,4);
TASK_PP(16'h1B04C,4);
TASK_PP(16'h1B04D,4);
TASK_PP(16'h1B04E,4);
TASK_PP(16'h1B04F,4);
TASK_PP(16'h1B050,4);
TASK_PP(16'h1B051,4);
TASK_PP(16'h1B052,4);
TASK_PP(16'h1B053,4);
TASK_PP(16'h1B054,4);
TASK_PP(16'h1B055,4);
TASK_PP(16'h1B056,4);
TASK_PP(16'h1B057,4);
TASK_PP(16'h1B058,4);
TASK_PP(16'h1B059,4);
TASK_PP(16'h1B05A,4);
TASK_PP(16'h1B05B,4);
TASK_PP(16'h1B05C,4);
TASK_PP(16'h1B05D,4);
TASK_PP(16'h1B05E,4);
TASK_PP(16'h1B05F,4);
TASK_PP(16'h1B060,4);
TASK_PP(16'h1B061,4);
TASK_PP(16'h1B062,4);
TASK_PP(16'h1B063,4);
TASK_PP(16'h1B064,4);
TASK_PP(16'h1B065,4);
TASK_PP(16'h1B066,4);
TASK_PP(16'h1B067,4);
TASK_PP(16'h1B068,4);
TASK_PP(16'h1B069,4);
TASK_PP(16'h1B06A,4);
TASK_PP(16'h1B06B,4);
TASK_PP(16'h1B06C,4);
TASK_PP(16'h1B06D,4);
TASK_PP(16'h1B06E,4);
TASK_PP(16'h1B06F,4);
TASK_PP(16'h1B070,4);
TASK_PP(16'h1B071,4);
TASK_PP(16'h1B072,4);
TASK_PP(16'h1B073,4);
TASK_PP(16'h1B074,4);
TASK_PP(16'h1B075,4);
TASK_PP(16'h1B076,4);
TASK_PP(16'h1B077,4);
TASK_PP(16'h1B078,4);
TASK_PP(16'h1B079,4);
TASK_PP(16'h1B07A,4);
TASK_PP(16'h1B07B,4);
TASK_PP(16'h1B07C,4);
TASK_PP(16'h1B07D,4);
TASK_PP(16'h1B07E,4);
TASK_PP(16'h1B07F,4);
TASK_PP(16'h1B080,4);
TASK_PP(16'h1B081,4);
TASK_PP(16'h1B082,4);
TASK_PP(16'h1B083,4);
TASK_PP(16'h1B084,4);
TASK_PP(16'h1B085,4);
TASK_PP(16'h1B086,4);
TASK_PP(16'h1B087,4);
TASK_PP(16'h1B088,4);
TASK_PP(16'h1B089,4);
TASK_PP(16'h1B08A,4);
TASK_PP(16'h1B08B,4);
TASK_PP(16'h1B08C,4);
TASK_PP(16'h1B08D,4);
TASK_PP(16'h1B08E,4);
TASK_PP(16'h1B08F,4);
TASK_PP(16'h1B090,4);
TASK_PP(16'h1B091,4);
TASK_PP(16'h1B092,4);
TASK_PP(16'h1B093,4);
TASK_PP(16'h1B094,4);
TASK_PP(16'h1B095,4);
TASK_PP(16'h1B096,4);
TASK_PP(16'h1B097,4);
TASK_PP(16'h1B098,4);
TASK_PP(16'h1B099,4);
TASK_PP(16'h1B09A,4);
TASK_PP(16'h1B09B,4);
TASK_PP(16'h1B09C,4);
TASK_PP(16'h1B09D,4);
TASK_PP(16'h1B09E,4);
TASK_PP(16'h1B09F,4);
TASK_PP(16'h1B0A0,4);
TASK_PP(16'h1B0A1,4);
TASK_PP(16'h1B0A2,4);
TASK_PP(16'h1B0A3,4);
TASK_PP(16'h1B0A4,4);
TASK_PP(16'h1B0A5,4);
TASK_PP(16'h1B0A6,4);
TASK_PP(16'h1B0A7,4);
TASK_PP(16'h1B0A8,4);
TASK_PP(16'h1B0A9,4);
TASK_PP(16'h1B0AA,4);
TASK_PP(16'h1B0AB,4);
TASK_PP(16'h1B0AC,4);
TASK_PP(16'h1B0AD,4);
TASK_PP(16'h1B0AE,4);
TASK_PP(16'h1B0AF,4);
TASK_PP(16'h1B0B0,4);
TASK_PP(16'h1B0B1,4);
TASK_PP(16'h1B0B2,4);
TASK_PP(16'h1B0B3,4);
TASK_PP(16'h1B0B4,4);
TASK_PP(16'h1B0B5,4);
TASK_PP(16'h1B0B6,4);
TASK_PP(16'h1B0B7,4);
TASK_PP(16'h1B0B8,4);
TASK_PP(16'h1B0B9,4);
TASK_PP(16'h1B0BA,4);
TASK_PP(16'h1B0BB,4);
TASK_PP(16'h1B0BC,4);
TASK_PP(16'h1B0BD,4);
TASK_PP(16'h1B0BE,4);
TASK_PP(16'h1B0BF,4);
TASK_PP(16'h1B0C0,4);
TASK_PP(16'h1B0C1,4);
TASK_PP(16'h1B0C2,4);
TASK_PP(16'h1B0C3,4);
TASK_PP(16'h1B0C4,4);
TASK_PP(16'h1B0C5,4);
TASK_PP(16'h1B0C6,4);
TASK_PP(16'h1B0C7,4);
TASK_PP(16'h1B0C8,4);
TASK_PP(16'h1B0C9,4);
TASK_PP(16'h1B0CA,4);
TASK_PP(16'h1B0CB,4);
TASK_PP(16'h1B0CC,4);
TASK_PP(16'h1B0CD,4);
TASK_PP(16'h1B0CE,4);
TASK_PP(16'h1B0CF,4);
TASK_PP(16'h1B0D0,4);
TASK_PP(16'h1B0D1,4);
TASK_PP(16'h1B0D2,4);
TASK_PP(16'h1B0D3,4);
TASK_PP(16'h1B0D4,4);
TASK_PP(16'h1B0D5,4);
TASK_PP(16'h1B0D6,4);
TASK_PP(16'h1B0D7,4);
TASK_PP(16'h1B0D8,4);
TASK_PP(16'h1B0D9,4);
TASK_PP(16'h1B0DA,4);
TASK_PP(16'h1B0DB,4);
TASK_PP(16'h1B0DC,4);
TASK_PP(16'h1B0DD,4);
TASK_PP(16'h1B0DE,4);
TASK_PP(16'h1B0DF,4);
TASK_PP(16'h1B0E0,4);
TASK_PP(16'h1B0E1,4);
TASK_PP(16'h1B0E2,4);
TASK_PP(16'h1B0E3,4);
TASK_PP(16'h1B0E4,4);
TASK_PP(16'h1B0E5,4);
TASK_PP(16'h1B0E6,4);
TASK_PP(16'h1B0E7,4);
TASK_PP(16'h1B0E8,4);
TASK_PP(16'h1B0E9,4);
TASK_PP(16'h1B0EA,4);
TASK_PP(16'h1B0EB,4);
TASK_PP(16'h1B0EC,4);
TASK_PP(16'h1B0ED,4);
TASK_PP(16'h1B0EE,4);
TASK_PP(16'h1B0EF,4);
TASK_PP(16'h1B0F0,4);
TASK_PP(16'h1B0F1,4);
TASK_PP(16'h1B0F2,4);
TASK_PP(16'h1B0F3,4);
TASK_PP(16'h1B0F4,4);
TASK_PP(16'h1B0F5,4);
TASK_PP(16'h1B0F6,4);
TASK_PP(16'h1B0F7,4);
TASK_PP(16'h1B0F8,4);
TASK_PP(16'h1B0F9,4);
TASK_PP(16'h1B0FA,4);
TASK_PP(16'h1B0FB,4);
TASK_PP(16'h1B0FC,4);
TASK_PP(16'h1B0FD,4);
TASK_PP(16'h1B0FE,4);
TASK_PP(16'h1B0FF,4);
TASK_PP(16'h1B100,4);
TASK_PP(16'h1B101,4);
TASK_PP(16'h1B102,4);
TASK_PP(16'h1B103,4);
TASK_PP(16'h1B104,4);
TASK_PP(16'h1B105,4);
TASK_PP(16'h1B106,4);
TASK_PP(16'h1B107,4);
TASK_PP(16'h1B108,4);
TASK_PP(16'h1B109,4);
TASK_PP(16'h1B10A,4);
TASK_PP(16'h1B10B,4);
TASK_PP(16'h1B10C,4);
TASK_PP(16'h1B10D,4);
TASK_PP(16'h1B10E,4);
TASK_PP(16'h1B10F,4);
TASK_PP(16'h1B110,4);
TASK_PP(16'h1B111,4);
TASK_PP(16'h1B112,4);
TASK_PP(16'h1B113,4);
TASK_PP(16'h1B114,4);
TASK_PP(16'h1B115,4);
TASK_PP(16'h1B116,4);
TASK_PP(16'h1B117,4);
TASK_PP(16'h1B118,4);
TASK_PP(16'h1B119,4);
TASK_PP(16'h1B11A,4);
TASK_PP(16'h1B11B,4);
TASK_PP(16'h1B11C,4);
TASK_PP(16'h1B11D,4);
TASK_PP(16'h1B11E,4);
TASK_PP(16'h1B11F,4);
TASK_PP(16'h1B120,4);
TASK_PP(16'h1B121,4);
TASK_PP(16'h1B122,4);
TASK_PP(16'h1B123,4);
TASK_PP(16'h1B124,4);
TASK_PP(16'h1B125,4);
TASK_PP(16'h1B126,4);
TASK_PP(16'h1B127,4);
TASK_PP(16'h1B128,4);
TASK_PP(16'h1B129,4);
TASK_PP(16'h1B12A,4);
TASK_PP(16'h1B12B,4);
TASK_PP(16'h1B12C,4);
TASK_PP(16'h1B12D,4);
TASK_PP(16'h1B12E,4);
TASK_PP(16'h1B12F,4);
TASK_PP(16'h1B130,4);
TASK_PP(16'h1B131,4);
TASK_PP(16'h1B132,4);
TASK_PP(16'h1B133,4);
TASK_PP(16'h1B134,4);
TASK_PP(16'h1B135,4);
TASK_PP(16'h1B136,4);
TASK_PP(16'h1B137,4);
TASK_PP(16'h1B138,4);
TASK_PP(16'h1B139,4);
TASK_PP(16'h1B13A,4);
TASK_PP(16'h1B13B,4);
TASK_PP(16'h1B13C,4);
TASK_PP(16'h1B13D,4);
TASK_PP(16'h1B13E,4);
TASK_PP(16'h1B13F,4);
TASK_PP(16'h1B140,4);
TASK_PP(16'h1B141,4);
TASK_PP(16'h1B142,4);
TASK_PP(16'h1B143,4);
TASK_PP(16'h1B144,4);
TASK_PP(16'h1B145,4);
TASK_PP(16'h1B146,4);
TASK_PP(16'h1B147,4);
TASK_PP(16'h1B148,4);
TASK_PP(16'h1B149,4);
TASK_PP(16'h1B14A,4);
TASK_PP(16'h1B14B,4);
TASK_PP(16'h1B14C,4);
TASK_PP(16'h1B14D,4);
TASK_PP(16'h1B14E,4);
TASK_PP(16'h1B14F,4);
TASK_PP(16'h1B150,4);
TASK_PP(16'h1B151,4);
TASK_PP(16'h1B152,4);
TASK_PP(16'h1B153,4);
TASK_PP(16'h1B154,4);
TASK_PP(16'h1B155,4);
TASK_PP(16'h1B156,4);
TASK_PP(16'h1B157,4);
TASK_PP(16'h1B158,4);
TASK_PP(16'h1B159,4);
TASK_PP(16'h1B15A,4);
TASK_PP(16'h1B15B,4);
TASK_PP(16'h1B15C,4);
TASK_PP(16'h1B15D,4);
TASK_PP(16'h1B15E,4);
TASK_PP(16'h1B15F,4);
TASK_PP(16'h1B160,4);
TASK_PP(16'h1B161,4);
TASK_PP(16'h1B162,4);
TASK_PP(16'h1B163,4);
TASK_PP(16'h1B164,4);
TASK_PP(16'h1B165,4);
TASK_PP(16'h1B166,4);
TASK_PP(16'h1B167,4);
TASK_PP(16'h1B168,4);
TASK_PP(16'h1B169,4);
TASK_PP(16'h1B16A,4);
TASK_PP(16'h1B16B,4);
TASK_PP(16'h1B16C,4);
TASK_PP(16'h1B16D,4);
TASK_PP(16'h1B16E,4);
TASK_PP(16'h1B16F,4);
TASK_PP(16'h1B170,4);
TASK_PP(16'h1B171,4);
TASK_PP(16'h1B172,4);
TASK_PP(16'h1B173,4);
TASK_PP(16'h1B174,4);
TASK_PP(16'h1B175,4);
TASK_PP(16'h1B176,4);
TASK_PP(16'h1B177,4);
TASK_PP(16'h1B178,4);
TASK_PP(16'h1B179,4);
TASK_PP(16'h1B17A,4);
TASK_PP(16'h1B17B,4);
TASK_PP(16'h1B17C,4);
TASK_PP(16'h1B17D,4);
TASK_PP(16'h1B17E,4);
TASK_PP(16'h1B17F,4);
TASK_PP(16'h1B180,4);
TASK_PP(16'h1B181,4);
TASK_PP(16'h1B182,4);
TASK_PP(16'h1B183,4);
TASK_PP(16'h1B184,4);
TASK_PP(16'h1B185,4);
TASK_PP(16'h1B186,4);
TASK_PP(16'h1B187,4);
TASK_PP(16'h1B188,4);
TASK_PP(16'h1B189,4);
TASK_PP(16'h1B18A,4);
TASK_PP(16'h1B18B,4);
TASK_PP(16'h1B18C,4);
TASK_PP(16'h1B18D,4);
TASK_PP(16'h1B18E,4);
TASK_PP(16'h1B18F,4);
TASK_PP(16'h1B190,4);
TASK_PP(16'h1B191,4);
TASK_PP(16'h1B192,4);
TASK_PP(16'h1B193,4);
TASK_PP(16'h1B194,4);
TASK_PP(16'h1B195,4);
TASK_PP(16'h1B196,4);
TASK_PP(16'h1B197,4);
TASK_PP(16'h1B198,4);
TASK_PP(16'h1B199,4);
TASK_PP(16'h1B19A,4);
TASK_PP(16'h1B19B,4);
TASK_PP(16'h1B19C,4);
TASK_PP(16'h1B19D,4);
TASK_PP(16'h1B19E,4);
TASK_PP(16'h1B19F,4);
TASK_PP(16'h1B1A0,4);
TASK_PP(16'h1B1A1,4);
TASK_PP(16'h1B1A2,4);
TASK_PP(16'h1B1A3,4);
TASK_PP(16'h1B1A4,4);
TASK_PP(16'h1B1A5,4);
TASK_PP(16'h1B1A6,4);
TASK_PP(16'h1B1A7,4);
TASK_PP(16'h1B1A8,4);
TASK_PP(16'h1B1A9,4);
TASK_PP(16'h1B1AA,4);
TASK_PP(16'h1B1AB,4);
TASK_PP(16'h1B1AC,4);
TASK_PP(16'h1B1AD,4);
TASK_PP(16'h1B1AE,4);
TASK_PP(16'h1B1AF,4);
TASK_PP(16'h1B1B0,4);
TASK_PP(16'h1B1B1,4);
TASK_PP(16'h1B1B2,4);
TASK_PP(16'h1B1B3,4);
TASK_PP(16'h1B1B4,4);
TASK_PP(16'h1B1B5,4);
TASK_PP(16'h1B1B6,4);
TASK_PP(16'h1B1B7,4);
TASK_PP(16'h1B1B8,4);
TASK_PP(16'h1B1B9,4);
TASK_PP(16'h1B1BA,4);
TASK_PP(16'h1B1BB,4);
TASK_PP(16'h1B1BC,4);
TASK_PP(16'h1B1BD,4);
TASK_PP(16'h1B1BE,4);
TASK_PP(16'h1B1BF,4);
TASK_PP(16'h1B1C0,4);
TASK_PP(16'h1B1C1,4);
TASK_PP(16'h1B1C2,4);
TASK_PP(16'h1B1C3,4);
TASK_PP(16'h1B1C4,4);
TASK_PP(16'h1B1C5,4);
TASK_PP(16'h1B1C6,4);
TASK_PP(16'h1B1C7,4);
TASK_PP(16'h1B1C8,4);
TASK_PP(16'h1B1C9,4);
TASK_PP(16'h1B1CA,4);
TASK_PP(16'h1B1CB,4);
TASK_PP(16'h1B1CC,4);
TASK_PP(16'h1B1CD,4);
TASK_PP(16'h1B1CE,4);
TASK_PP(16'h1B1CF,4);
TASK_PP(16'h1B1D0,4);
TASK_PP(16'h1B1D1,4);
TASK_PP(16'h1B1D2,4);
TASK_PP(16'h1B1D3,4);
TASK_PP(16'h1B1D4,4);
TASK_PP(16'h1B1D5,4);
TASK_PP(16'h1B1D6,4);
TASK_PP(16'h1B1D7,4);
TASK_PP(16'h1B1D8,4);
TASK_PP(16'h1B1D9,4);
TASK_PP(16'h1B1DA,4);
TASK_PP(16'h1B1DB,4);
TASK_PP(16'h1B1DC,4);
TASK_PP(16'h1B1DD,4);
TASK_PP(16'h1B1DE,4);
TASK_PP(16'h1B1DF,4);
TASK_PP(16'h1B1E0,4);
TASK_PP(16'h1B1E1,4);
TASK_PP(16'h1B1E2,4);
TASK_PP(16'h1B1E3,4);
TASK_PP(16'h1B1E4,4);
TASK_PP(16'h1B1E5,4);
TASK_PP(16'h1B1E6,4);
TASK_PP(16'h1B1E7,4);
TASK_PP(16'h1B1E8,4);
TASK_PP(16'h1B1E9,4);
TASK_PP(16'h1B1EA,4);
TASK_PP(16'h1B1EB,4);
TASK_PP(16'h1B1EC,4);
TASK_PP(16'h1B1ED,4);
TASK_PP(16'h1B1EE,4);
TASK_PP(16'h1B1EF,4);
TASK_PP(16'h1B1F0,4);
TASK_PP(16'h1B1F1,4);
TASK_PP(16'h1B1F2,4);
TASK_PP(16'h1B1F3,4);
TASK_PP(16'h1B1F4,4);
TASK_PP(16'h1B1F5,4);
TASK_PP(16'h1B1F6,4);
TASK_PP(16'h1B1F7,4);
TASK_PP(16'h1B1F8,4);
TASK_PP(16'h1B1F9,4);
TASK_PP(16'h1B1FA,4);
TASK_PP(16'h1B1FB,4);
TASK_PP(16'h1B1FC,4);
TASK_PP(16'h1B1FD,4);
TASK_PP(16'h1B1FE,4);
TASK_PP(16'h1B1FF,4);
TASK_PP(16'h1B200,4);
TASK_PP(16'h1B201,4);
TASK_PP(16'h1B202,4);
TASK_PP(16'h1B203,4);
TASK_PP(16'h1B204,4);
TASK_PP(16'h1B205,4);
TASK_PP(16'h1B206,4);
TASK_PP(16'h1B207,4);
TASK_PP(16'h1B208,4);
TASK_PP(16'h1B209,4);
TASK_PP(16'h1B20A,4);
TASK_PP(16'h1B20B,4);
TASK_PP(16'h1B20C,4);
TASK_PP(16'h1B20D,4);
TASK_PP(16'h1B20E,4);
TASK_PP(16'h1B20F,4);
TASK_PP(16'h1B210,4);
TASK_PP(16'h1B211,4);
TASK_PP(16'h1B212,4);
TASK_PP(16'h1B213,4);
TASK_PP(16'h1B214,4);
TASK_PP(16'h1B215,4);
TASK_PP(16'h1B216,4);
TASK_PP(16'h1B217,4);
TASK_PP(16'h1B218,4);
TASK_PP(16'h1B219,4);
TASK_PP(16'h1B21A,4);
TASK_PP(16'h1B21B,4);
TASK_PP(16'h1B21C,4);
TASK_PP(16'h1B21D,4);
TASK_PP(16'h1B21E,4);
TASK_PP(16'h1B21F,4);
TASK_PP(16'h1B220,4);
TASK_PP(16'h1B221,4);
TASK_PP(16'h1B222,4);
TASK_PP(16'h1B223,4);
TASK_PP(16'h1B224,4);
TASK_PP(16'h1B225,4);
TASK_PP(16'h1B226,4);
TASK_PP(16'h1B227,4);
TASK_PP(16'h1B228,4);
TASK_PP(16'h1B229,4);
TASK_PP(16'h1B22A,4);
TASK_PP(16'h1B22B,4);
TASK_PP(16'h1B22C,4);
TASK_PP(16'h1B22D,4);
TASK_PP(16'h1B22E,4);
TASK_PP(16'h1B22F,4);
TASK_PP(16'h1B230,4);
TASK_PP(16'h1B231,4);
TASK_PP(16'h1B232,4);
TASK_PP(16'h1B233,4);
TASK_PP(16'h1B234,4);
TASK_PP(16'h1B235,4);
TASK_PP(16'h1B236,4);
TASK_PP(16'h1B237,4);
TASK_PP(16'h1B238,4);
TASK_PP(16'h1B239,4);
TASK_PP(16'h1B23A,4);
TASK_PP(16'h1B23B,4);
TASK_PP(16'h1B23C,4);
TASK_PP(16'h1B23D,4);
TASK_PP(16'h1B23E,4);
TASK_PP(16'h1B23F,4);
TASK_PP(16'h1B240,4);
TASK_PP(16'h1B241,4);
TASK_PP(16'h1B242,4);
TASK_PP(16'h1B243,4);
TASK_PP(16'h1B244,4);
TASK_PP(16'h1B245,4);
TASK_PP(16'h1B246,4);
TASK_PP(16'h1B247,4);
TASK_PP(16'h1B248,4);
TASK_PP(16'h1B249,4);
TASK_PP(16'h1B24A,4);
TASK_PP(16'h1B24B,4);
TASK_PP(16'h1B24C,4);
TASK_PP(16'h1B24D,4);
TASK_PP(16'h1B24E,4);
TASK_PP(16'h1B24F,4);
TASK_PP(16'h1B250,4);
TASK_PP(16'h1B251,4);
TASK_PP(16'h1B252,4);
TASK_PP(16'h1B253,4);
TASK_PP(16'h1B254,4);
TASK_PP(16'h1B255,4);
TASK_PP(16'h1B256,4);
TASK_PP(16'h1B257,4);
TASK_PP(16'h1B258,4);
TASK_PP(16'h1B259,4);
TASK_PP(16'h1B25A,4);
TASK_PP(16'h1B25B,4);
TASK_PP(16'h1B25C,4);
TASK_PP(16'h1B25D,4);
TASK_PP(16'h1B25E,4);
TASK_PP(16'h1B25F,4);
TASK_PP(16'h1B260,4);
TASK_PP(16'h1B261,4);
TASK_PP(16'h1B262,4);
TASK_PP(16'h1B263,4);
TASK_PP(16'h1B264,4);
TASK_PP(16'h1B265,4);
TASK_PP(16'h1B266,4);
TASK_PP(16'h1B267,4);
TASK_PP(16'h1B268,4);
TASK_PP(16'h1B269,4);
TASK_PP(16'h1B26A,4);
TASK_PP(16'h1B26B,4);
TASK_PP(16'h1B26C,4);
TASK_PP(16'h1B26D,4);
TASK_PP(16'h1B26E,4);
TASK_PP(16'h1B26F,4);
TASK_PP(16'h1B270,4);
TASK_PP(16'h1B271,4);
TASK_PP(16'h1B272,4);
TASK_PP(16'h1B273,4);
TASK_PP(16'h1B274,4);
TASK_PP(16'h1B275,4);
TASK_PP(16'h1B276,4);
TASK_PP(16'h1B277,4);
TASK_PP(16'h1B278,4);
TASK_PP(16'h1B279,4);
TASK_PP(16'h1B27A,4);
TASK_PP(16'h1B27B,4);
TASK_PP(16'h1B27C,4);
TASK_PP(16'h1B27D,4);
TASK_PP(16'h1B27E,4);
TASK_PP(16'h1B27F,4);
TASK_PP(16'h1B280,4);
TASK_PP(16'h1B281,4);
TASK_PP(16'h1B282,4);
TASK_PP(16'h1B283,4);
TASK_PP(16'h1B284,4);
TASK_PP(16'h1B285,4);
TASK_PP(16'h1B286,4);
TASK_PP(16'h1B287,4);
TASK_PP(16'h1B288,4);
TASK_PP(16'h1B289,4);
TASK_PP(16'h1B28A,4);
TASK_PP(16'h1B28B,4);
TASK_PP(16'h1B28C,4);
TASK_PP(16'h1B28D,4);
TASK_PP(16'h1B28E,4);
TASK_PP(16'h1B28F,4);
TASK_PP(16'h1B290,4);
TASK_PP(16'h1B291,4);
TASK_PP(16'h1B292,4);
TASK_PP(16'h1B293,4);
TASK_PP(16'h1B294,4);
TASK_PP(16'h1B295,4);
TASK_PP(16'h1B296,4);
TASK_PP(16'h1B297,4);
TASK_PP(16'h1B298,4);
TASK_PP(16'h1B299,4);
TASK_PP(16'h1B29A,4);
TASK_PP(16'h1B29B,4);
TASK_PP(16'h1B29C,4);
TASK_PP(16'h1B29D,4);
TASK_PP(16'h1B29E,4);
TASK_PP(16'h1B29F,4);
TASK_PP(16'h1B2A0,4);
TASK_PP(16'h1B2A1,4);
TASK_PP(16'h1B2A2,4);
TASK_PP(16'h1B2A3,4);
TASK_PP(16'h1B2A4,4);
TASK_PP(16'h1B2A5,4);
TASK_PP(16'h1B2A6,4);
TASK_PP(16'h1B2A7,4);
TASK_PP(16'h1B2A8,4);
TASK_PP(16'h1B2A9,4);
TASK_PP(16'h1B2AA,4);
TASK_PP(16'h1B2AB,4);
TASK_PP(16'h1B2AC,4);
TASK_PP(16'h1B2AD,4);
TASK_PP(16'h1B2AE,4);
TASK_PP(16'h1B2AF,4);
TASK_PP(16'h1B2B0,4);
TASK_PP(16'h1B2B1,4);
TASK_PP(16'h1B2B2,4);
TASK_PP(16'h1B2B3,4);
TASK_PP(16'h1B2B4,4);
TASK_PP(16'h1B2B5,4);
TASK_PP(16'h1B2B6,4);
TASK_PP(16'h1B2B7,4);
TASK_PP(16'h1B2B8,4);
TASK_PP(16'h1B2B9,4);
TASK_PP(16'h1B2BA,4);
TASK_PP(16'h1B2BB,4);
TASK_PP(16'h1B2BC,4);
TASK_PP(16'h1B2BD,4);
TASK_PP(16'h1B2BE,4);
TASK_PP(16'h1B2BF,4);
TASK_PP(16'h1B2C0,4);
TASK_PP(16'h1B2C1,4);
TASK_PP(16'h1B2C2,4);
TASK_PP(16'h1B2C3,4);
TASK_PP(16'h1B2C4,4);
TASK_PP(16'h1B2C5,4);
TASK_PP(16'h1B2C6,4);
TASK_PP(16'h1B2C7,4);
TASK_PP(16'h1B2C8,4);
TASK_PP(16'h1B2C9,4);
TASK_PP(16'h1B2CA,4);
TASK_PP(16'h1B2CB,4);
TASK_PP(16'h1B2CC,4);
TASK_PP(16'h1B2CD,4);
TASK_PP(16'h1B2CE,4);
TASK_PP(16'h1B2CF,4);
TASK_PP(16'h1B2D0,4);
TASK_PP(16'h1B2D1,4);
TASK_PP(16'h1B2D2,4);
TASK_PP(16'h1B2D3,4);
TASK_PP(16'h1B2D4,4);
TASK_PP(16'h1B2D5,4);
TASK_PP(16'h1B2D6,4);
TASK_PP(16'h1B2D7,4);
TASK_PP(16'h1B2D8,4);
TASK_PP(16'h1B2D9,4);
TASK_PP(16'h1B2DA,4);
TASK_PP(16'h1B2DB,4);
TASK_PP(16'h1B2DC,4);
TASK_PP(16'h1B2DD,4);
TASK_PP(16'h1B2DE,4);
TASK_PP(16'h1B2DF,4);
TASK_PP(16'h1B2E0,4);
TASK_PP(16'h1B2E1,4);
TASK_PP(16'h1B2E2,4);
TASK_PP(16'h1B2E3,4);
TASK_PP(16'h1B2E4,4);
TASK_PP(16'h1B2E5,4);
TASK_PP(16'h1B2E6,4);
TASK_PP(16'h1B2E7,4);
TASK_PP(16'h1B2E8,4);
TASK_PP(16'h1B2E9,4);
TASK_PP(16'h1B2EA,4);
TASK_PP(16'h1B2EB,4);
TASK_PP(16'h1B2EC,4);
TASK_PP(16'h1B2ED,4);
TASK_PP(16'h1B2EE,4);
TASK_PP(16'h1B2EF,4);
TASK_PP(16'h1B2F0,4);
TASK_PP(16'h1B2F1,4);
TASK_PP(16'h1B2F2,4);
TASK_PP(16'h1B2F3,4);
TASK_PP(16'h1B2F4,4);
TASK_PP(16'h1B2F5,4);
TASK_PP(16'h1B2F6,4);
TASK_PP(16'h1B2F7,4);
TASK_PP(16'h1B2F8,4);
TASK_PP(16'h1B2F9,4);
TASK_PP(16'h1B2FA,4);
TASK_PP(16'h1B2FB,4);
TASK_PP(16'h1B2FC,4);
TASK_PP(16'h1B2FD,4);
TASK_PP(16'h1B2FE,4);
TASK_PP(16'h1B2FF,4);
TASK_PP(16'h1B300,4);
TASK_PP(16'h1B301,4);
TASK_PP(16'h1B302,4);
TASK_PP(16'h1B303,4);
TASK_PP(16'h1B304,4);
TASK_PP(16'h1B305,4);
TASK_PP(16'h1B306,4);
TASK_PP(16'h1B307,4);
TASK_PP(16'h1B308,4);
TASK_PP(16'h1B309,4);
TASK_PP(16'h1B30A,4);
TASK_PP(16'h1B30B,4);
TASK_PP(16'h1B30C,4);
TASK_PP(16'h1B30D,4);
TASK_PP(16'h1B30E,4);
TASK_PP(16'h1B30F,4);
TASK_PP(16'h1B310,4);
TASK_PP(16'h1B311,4);
TASK_PP(16'h1B312,4);
TASK_PP(16'h1B313,4);
TASK_PP(16'h1B314,4);
TASK_PP(16'h1B315,4);
TASK_PP(16'h1B316,4);
TASK_PP(16'h1B317,4);
TASK_PP(16'h1B318,4);
TASK_PP(16'h1B319,4);
TASK_PP(16'h1B31A,4);
TASK_PP(16'h1B31B,4);
TASK_PP(16'h1B31C,4);
TASK_PP(16'h1B31D,4);
TASK_PP(16'h1B31E,4);
TASK_PP(16'h1B31F,4);
TASK_PP(16'h1B320,4);
TASK_PP(16'h1B321,4);
TASK_PP(16'h1B322,4);
TASK_PP(16'h1B323,4);
TASK_PP(16'h1B324,4);
TASK_PP(16'h1B325,4);
TASK_PP(16'h1B326,4);
TASK_PP(16'h1B327,4);
TASK_PP(16'h1B328,4);
TASK_PP(16'h1B329,4);
TASK_PP(16'h1B32A,4);
TASK_PP(16'h1B32B,4);
TASK_PP(16'h1B32C,4);
TASK_PP(16'h1B32D,4);
TASK_PP(16'h1B32E,4);
TASK_PP(16'h1B32F,4);
TASK_PP(16'h1B330,4);
TASK_PP(16'h1B331,4);
TASK_PP(16'h1B332,4);
TASK_PP(16'h1B333,4);
TASK_PP(16'h1B334,4);
TASK_PP(16'h1B335,4);
TASK_PP(16'h1B336,4);
TASK_PP(16'h1B337,4);
TASK_PP(16'h1B338,4);
TASK_PP(16'h1B339,4);
TASK_PP(16'h1B33A,4);
TASK_PP(16'h1B33B,4);
TASK_PP(16'h1B33C,4);
TASK_PP(16'h1B33D,4);
TASK_PP(16'h1B33E,4);
TASK_PP(16'h1B33F,4);
TASK_PP(16'h1B340,4);
TASK_PP(16'h1B341,4);
TASK_PP(16'h1B342,4);
TASK_PP(16'h1B343,4);
TASK_PP(16'h1B344,4);
TASK_PP(16'h1B345,4);
TASK_PP(16'h1B346,4);
TASK_PP(16'h1B347,4);
TASK_PP(16'h1B348,4);
TASK_PP(16'h1B349,4);
TASK_PP(16'h1B34A,4);
TASK_PP(16'h1B34B,4);
TASK_PP(16'h1B34C,4);
TASK_PP(16'h1B34D,4);
TASK_PP(16'h1B34E,4);
TASK_PP(16'h1B34F,4);
TASK_PP(16'h1B350,4);
TASK_PP(16'h1B351,4);
TASK_PP(16'h1B352,4);
TASK_PP(16'h1B353,4);
TASK_PP(16'h1B354,4);
TASK_PP(16'h1B355,4);
TASK_PP(16'h1B356,4);
TASK_PP(16'h1B357,4);
TASK_PP(16'h1B358,4);
TASK_PP(16'h1B359,4);
TASK_PP(16'h1B35A,4);
TASK_PP(16'h1B35B,4);
TASK_PP(16'h1B35C,4);
TASK_PP(16'h1B35D,4);
TASK_PP(16'h1B35E,4);
TASK_PP(16'h1B35F,4);
TASK_PP(16'h1B360,4);
TASK_PP(16'h1B361,4);
TASK_PP(16'h1B362,4);
TASK_PP(16'h1B363,4);
TASK_PP(16'h1B364,4);
TASK_PP(16'h1B365,4);
TASK_PP(16'h1B366,4);
TASK_PP(16'h1B367,4);
TASK_PP(16'h1B368,4);
TASK_PP(16'h1B369,4);
TASK_PP(16'h1B36A,4);
TASK_PP(16'h1B36B,4);
TASK_PP(16'h1B36C,4);
TASK_PP(16'h1B36D,4);
TASK_PP(16'h1B36E,4);
TASK_PP(16'h1B36F,4);
TASK_PP(16'h1B370,4);
TASK_PP(16'h1B371,4);
TASK_PP(16'h1B372,4);
TASK_PP(16'h1B373,4);
TASK_PP(16'h1B374,4);
TASK_PP(16'h1B375,4);
TASK_PP(16'h1B376,4);
TASK_PP(16'h1B377,4);
TASK_PP(16'h1B378,4);
TASK_PP(16'h1B379,4);
TASK_PP(16'h1B37A,4);
TASK_PP(16'h1B37B,4);
TASK_PP(16'h1B37C,4);
TASK_PP(16'h1B37D,4);
TASK_PP(16'h1B37E,4);
TASK_PP(16'h1B37F,4);
TASK_PP(16'h1B380,4);
TASK_PP(16'h1B381,4);
TASK_PP(16'h1B382,4);
TASK_PP(16'h1B383,4);
TASK_PP(16'h1B384,4);
TASK_PP(16'h1B385,4);
TASK_PP(16'h1B386,4);
TASK_PP(16'h1B387,4);
TASK_PP(16'h1B388,4);
TASK_PP(16'h1B389,4);
TASK_PP(16'h1B38A,4);
TASK_PP(16'h1B38B,4);
TASK_PP(16'h1B38C,4);
TASK_PP(16'h1B38D,4);
TASK_PP(16'h1B38E,4);
TASK_PP(16'h1B38F,4);
TASK_PP(16'h1B390,4);
TASK_PP(16'h1B391,4);
TASK_PP(16'h1B392,4);
TASK_PP(16'h1B393,4);
TASK_PP(16'h1B394,4);
TASK_PP(16'h1B395,4);
TASK_PP(16'h1B396,4);
TASK_PP(16'h1B397,4);
TASK_PP(16'h1B398,4);
TASK_PP(16'h1B399,4);
TASK_PP(16'h1B39A,4);
TASK_PP(16'h1B39B,4);
TASK_PP(16'h1B39C,4);
TASK_PP(16'h1B39D,4);
TASK_PP(16'h1B39E,4);
TASK_PP(16'h1B39F,4);
TASK_PP(16'h1B3A0,4);
TASK_PP(16'h1B3A1,4);
TASK_PP(16'h1B3A2,4);
TASK_PP(16'h1B3A3,4);
TASK_PP(16'h1B3A4,4);
TASK_PP(16'h1B3A5,4);
TASK_PP(16'h1B3A6,4);
TASK_PP(16'h1B3A7,4);
TASK_PP(16'h1B3A8,4);
TASK_PP(16'h1B3A9,4);
TASK_PP(16'h1B3AA,4);
TASK_PP(16'h1B3AB,4);
TASK_PP(16'h1B3AC,4);
TASK_PP(16'h1B3AD,4);
TASK_PP(16'h1B3AE,4);
TASK_PP(16'h1B3AF,4);
TASK_PP(16'h1B3B0,4);
TASK_PP(16'h1B3B1,4);
TASK_PP(16'h1B3B2,4);
TASK_PP(16'h1B3B3,4);
TASK_PP(16'h1B3B4,4);
TASK_PP(16'h1B3B5,4);
TASK_PP(16'h1B3B6,4);
TASK_PP(16'h1B3B7,4);
TASK_PP(16'h1B3B8,4);
TASK_PP(16'h1B3B9,4);
TASK_PP(16'h1B3BA,4);
TASK_PP(16'h1B3BB,4);
TASK_PP(16'h1B3BC,4);
TASK_PP(16'h1B3BD,4);
TASK_PP(16'h1B3BE,4);
TASK_PP(16'h1B3BF,4);
TASK_PP(16'h1B3C0,4);
TASK_PP(16'h1B3C1,4);
TASK_PP(16'h1B3C2,4);
TASK_PP(16'h1B3C3,4);
TASK_PP(16'h1B3C4,4);
TASK_PP(16'h1B3C5,4);
TASK_PP(16'h1B3C6,4);
TASK_PP(16'h1B3C7,4);
TASK_PP(16'h1B3C8,4);
TASK_PP(16'h1B3C9,4);
TASK_PP(16'h1B3CA,4);
TASK_PP(16'h1B3CB,4);
TASK_PP(16'h1B3CC,4);
TASK_PP(16'h1B3CD,4);
TASK_PP(16'h1B3CE,4);
TASK_PP(16'h1B3CF,4);
TASK_PP(16'h1B3D0,4);
TASK_PP(16'h1B3D1,4);
TASK_PP(16'h1B3D2,4);
TASK_PP(16'h1B3D3,4);
TASK_PP(16'h1B3D4,4);
TASK_PP(16'h1B3D5,4);
TASK_PP(16'h1B3D6,4);
TASK_PP(16'h1B3D7,4);
TASK_PP(16'h1B3D8,4);
TASK_PP(16'h1B3D9,4);
TASK_PP(16'h1B3DA,4);
TASK_PP(16'h1B3DB,4);
TASK_PP(16'h1B3DC,4);
TASK_PP(16'h1B3DD,4);
TASK_PP(16'h1B3DE,4);
TASK_PP(16'h1B3DF,4);
TASK_PP(16'h1B3E0,4);
TASK_PP(16'h1B3E1,4);
TASK_PP(16'h1B3E2,4);
TASK_PP(16'h1B3E3,4);
TASK_PP(16'h1B3E4,4);
TASK_PP(16'h1B3E5,4);
TASK_PP(16'h1B3E6,4);
TASK_PP(16'h1B3E7,4);
TASK_PP(16'h1B3E8,4);
TASK_PP(16'h1B3E9,4);
TASK_PP(16'h1B3EA,4);
TASK_PP(16'h1B3EB,4);
TASK_PP(16'h1B3EC,4);
TASK_PP(16'h1B3ED,4);
TASK_PP(16'h1B3EE,4);
TASK_PP(16'h1B3EF,4);
TASK_PP(16'h1B3F0,4);
TASK_PP(16'h1B3F1,4);
TASK_PP(16'h1B3F2,4);
TASK_PP(16'h1B3F3,4);
TASK_PP(16'h1B3F4,4);
TASK_PP(16'h1B3F5,4);
TASK_PP(16'h1B3F6,4);
TASK_PP(16'h1B3F7,4);
TASK_PP(16'h1B3F8,4);
TASK_PP(16'h1B3F9,4);
TASK_PP(16'h1B3FA,4);
TASK_PP(16'h1B3FB,4);
TASK_PP(16'h1B3FC,4);
TASK_PP(16'h1B3FD,4);
TASK_PP(16'h1B3FE,4);
TASK_PP(16'h1B3FF,4);
TASK_PP(16'h1B400,4);
TASK_PP(16'h1B401,4);
TASK_PP(16'h1B402,4);
TASK_PP(16'h1B403,4);
TASK_PP(16'h1B404,4);
TASK_PP(16'h1B405,4);
TASK_PP(16'h1B406,4);
TASK_PP(16'h1B407,4);
TASK_PP(16'h1B408,4);
TASK_PP(16'h1B409,4);
TASK_PP(16'h1B40A,4);
TASK_PP(16'h1B40B,4);
TASK_PP(16'h1B40C,4);
TASK_PP(16'h1B40D,4);
TASK_PP(16'h1B40E,4);
TASK_PP(16'h1B40F,4);
TASK_PP(16'h1B410,4);
TASK_PP(16'h1B411,4);
TASK_PP(16'h1B412,4);
TASK_PP(16'h1B413,4);
TASK_PP(16'h1B414,4);
TASK_PP(16'h1B415,4);
TASK_PP(16'h1B416,4);
TASK_PP(16'h1B417,4);
TASK_PP(16'h1B418,4);
TASK_PP(16'h1B419,4);
TASK_PP(16'h1B41A,4);
TASK_PP(16'h1B41B,4);
TASK_PP(16'h1B41C,4);
TASK_PP(16'h1B41D,4);
TASK_PP(16'h1B41E,4);
TASK_PP(16'h1B41F,4);
TASK_PP(16'h1B420,4);
TASK_PP(16'h1B421,4);
TASK_PP(16'h1B422,4);
TASK_PP(16'h1B423,4);
TASK_PP(16'h1B424,4);
TASK_PP(16'h1B425,4);
TASK_PP(16'h1B426,4);
TASK_PP(16'h1B427,4);
TASK_PP(16'h1B428,4);
TASK_PP(16'h1B429,4);
TASK_PP(16'h1B42A,4);
TASK_PP(16'h1B42B,4);
TASK_PP(16'h1B42C,4);
TASK_PP(16'h1B42D,4);
TASK_PP(16'h1B42E,4);
TASK_PP(16'h1B42F,4);
TASK_PP(16'h1B430,4);
TASK_PP(16'h1B431,4);
TASK_PP(16'h1B432,4);
TASK_PP(16'h1B433,4);
TASK_PP(16'h1B434,4);
TASK_PP(16'h1B435,4);
TASK_PP(16'h1B436,4);
TASK_PP(16'h1B437,4);
TASK_PP(16'h1B438,4);
TASK_PP(16'h1B439,4);
TASK_PP(16'h1B43A,4);
TASK_PP(16'h1B43B,4);
TASK_PP(16'h1B43C,4);
TASK_PP(16'h1B43D,4);
TASK_PP(16'h1B43E,4);
TASK_PP(16'h1B43F,4);
TASK_PP(16'h1B440,4);
TASK_PP(16'h1B441,4);
TASK_PP(16'h1B442,4);
TASK_PP(16'h1B443,4);
TASK_PP(16'h1B444,4);
TASK_PP(16'h1B445,4);
TASK_PP(16'h1B446,4);
TASK_PP(16'h1B447,4);
TASK_PP(16'h1B448,4);
TASK_PP(16'h1B449,4);
TASK_PP(16'h1B44A,4);
TASK_PP(16'h1B44B,4);
TASK_PP(16'h1B44C,4);
TASK_PP(16'h1B44D,4);
TASK_PP(16'h1B44E,4);
TASK_PP(16'h1B44F,4);
TASK_PP(16'h1B450,4);
TASK_PP(16'h1B451,4);
TASK_PP(16'h1B452,4);
TASK_PP(16'h1B453,4);
TASK_PP(16'h1B454,4);
TASK_PP(16'h1B455,4);
TASK_PP(16'h1B456,4);
TASK_PP(16'h1B457,4);
TASK_PP(16'h1B458,4);
TASK_PP(16'h1B459,4);
TASK_PP(16'h1B45A,4);
TASK_PP(16'h1B45B,4);
TASK_PP(16'h1B45C,4);
TASK_PP(16'h1B45D,4);
TASK_PP(16'h1B45E,4);
TASK_PP(16'h1B45F,4);
TASK_PP(16'h1B460,4);
TASK_PP(16'h1B461,4);
TASK_PP(16'h1B462,4);
TASK_PP(16'h1B463,4);
TASK_PP(16'h1B464,4);
TASK_PP(16'h1B465,4);
TASK_PP(16'h1B466,4);
TASK_PP(16'h1B467,4);
TASK_PP(16'h1B468,4);
TASK_PP(16'h1B469,4);
TASK_PP(16'h1B46A,4);
TASK_PP(16'h1B46B,4);
TASK_PP(16'h1B46C,4);
TASK_PP(16'h1B46D,4);
TASK_PP(16'h1B46E,4);
TASK_PP(16'h1B46F,4);
TASK_PP(16'h1B470,4);
TASK_PP(16'h1B471,4);
TASK_PP(16'h1B472,4);
TASK_PP(16'h1B473,4);
TASK_PP(16'h1B474,4);
TASK_PP(16'h1B475,4);
TASK_PP(16'h1B476,4);
TASK_PP(16'h1B477,4);
TASK_PP(16'h1B478,4);
TASK_PP(16'h1B479,4);
TASK_PP(16'h1B47A,4);
TASK_PP(16'h1B47B,4);
TASK_PP(16'h1B47C,4);
TASK_PP(16'h1B47D,4);
TASK_PP(16'h1B47E,4);
TASK_PP(16'h1B47F,4);
TASK_PP(16'h1B480,4);
TASK_PP(16'h1B481,4);
TASK_PP(16'h1B482,4);
TASK_PP(16'h1B483,4);
TASK_PP(16'h1B484,4);
TASK_PP(16'h1B485,4);
TASK_PP(16'h1B486,4);
TASK_PP(16'h1B487,4);
TASK_PP(16'h1B488,4);
TASK_PP(16'h1B489,4);
TASK_PP(16'h1B48A,4);
TASK_PP(16'h1B48B,4);
TASK_PP(16'h1B48C,4);
TASK_PP(16'h1B48D,4);
TASK_PP(16'h1B48E,4);
TASK_PP(16'h1B48F,4);
TASK_PP(16'h1B490,4);
TASK_PP(16'h1B491,4);
TASK_PP(16'h1B492,4);
TASK_PP(16'h1B493,4);
TASK_PP(16'h1B494,4);
TASK_PP(16'h1B495,4);
TASK_PP(16'h1B496,4);
TASK_PP(16'h1B497,4);
TASK_PP(16'h1B498,4);
TASK_PP(16'h1B499,4);
TASK_PP(16'h1B49A,4);
TASK_PP(16'h1B49B,4);
TASK_PP(16'h1B49C,4);
TASK_PP(16'h1B49D,4);
TASK_PP(16'h1B49E,4);
TASK_PP(16'h1B49F,4);
TASK_PP(16'h1B4A0,4);
TASK_PP(16'h1B4A1,4);
TASK_PP(16'h1B4A2,4);
TASK_PP(16'h1B4A3,4);
TASK_PP(16'h1B4A4,4);
TASK_PP(16'h1B4A5,4);
TASK_PP(16'h1B4A6,4);
TASK_PP(16'h1B4A7,4);
TASK_PP(16'h1B4A8,4);
TASK_PP(16'h1B4A9,4);
TASK_PP(16'h1B4AA,4);
TASK_PP(16'h1B4AB,4);
TASK_PP(16'h1B4AC,4);
TASK_PP(16'h1B4AD,4);
TASK_PP(16'h1B4AE,4);
TASK_PP(16'h1B4AF,4);
TASK_PP(16'h1B4B0,4);
TASK_PP(16'h1B4B1,4);
TASK_PP(16'h1B4B2,4);
TASK_PP(16'h1B4B3,4);
TASK_PP(16'h1B4B4,4);
TASK_PP(16'h1B4B5,4);
TASK_PP(16'h1B4B6,4);
TASK_PP(16'h1B4B7,4);
TASK_PP(16'h1B4B8,4);
TASK_PP(16'h1B4B9,4);
TASK_PP(16'h1B4BA,4);
TASK_PP(16'h1B4BB,4);
TASK_PP(16'h1B4BC,4);
TASK_PP(16'h1B4BD,4);
TASK_PP(16'h1B4BE,4);
TASK_PP(16'h1B4BF,4);
TASK_PP(16'h1B4C0,4);
TASK_PP(16'h1B4C1,4);
TASK_PP(16'h1B4C2,4);
TASK_PP(16'h1B4C3,4);
TASK_PP(16'h1B4C4,4);
TASK_PP(16'h1B4C5,4);
TASK_PP(16'h1B4C6,4);
TASK_PP(16'h1B4C7,4);
TASK_PP(16'h1B4C8,4);
TASK_PP(16'h1B4C9,4);
TASK_PP(16'h1B4CA,4);
TASK_PP(16'h1B4CB,4);
TASK_PP(16'h1B4CC,4);
TASK_PP(16'h1B4CD,4);
TASK_PP(16'h1B4CE,4);
TASK_PP(16'h1B4CF,4);
TASK_PP(16'h1B4D0,4);
TASK_PP(16'h1B4D1,4);
TASK_PP(16'h1B4D2,4);
TASK_PP(16'h1B4D3,4);
TASK_PP(16'h1B4D4,4);
TASK_PP(16'h1B4D5,4);
TASK_PP(16'h1B4D6,4);
TASK_PP(16'h1B4D7,4);
TASK_PP(16'h1B4D8,4);
TASK_PP(16'h1B4D9,4);
TASK_PP(16'h1B4DA,4);
TASK_PP(16'h1B4DB,4);
TASK_PP(16'h1B4DC,4);
TASK_PP(16'h1B4DD,4);
TASK_PP(16'h1B4DE,4);
TASK_PP(16'h1B4DF,4);
TASK_PP(16'h1B4E0,4);
TASK_PP(16'h1B4E1,4);
TASK_PP(16'h1B4E2,4);
TASK_PP(16'h1B4E3,4);
TASK_PP(16'h1B4E4,4);
TASK_PP(16'h1B4E5,4);
TASK_PP(16'h1B4E6,4);
TASK_PP(16'h1B4E7,4);
TASK_PP(16'h1B4E8,4);
TASK_PP(16'h1B4E9,4);
TASK_PP(16'h1B4EA,4);
TASK_PP(16'h1B4EB,4);
TASK_PP(16'h1B4EC,4);
TASK_PP(16'h1B4ED,4);
TASK_PP(16'h1B4EE,4);
TASK_PP(16'h1B4EF,4);
TASK_PP(16'h1B4F0,4);
TASK_PP(16'h1B4F1,4);
TASK_PP(16'h1B4F2,4);
TASK_PP(16'h1B4F3,4);
TASK_PP(16'h1B4F4,4);
TASK_PP(16'h1B4F5,4);
TASK_PP(16'h1B4F6,4);
TASK_PP(16'h1B4F7,4);
TASK_PP(16'h1B4F8,4);
TASK_PP(16'h1B4F9,4);
TASK_PP(16'h1B4FA,4);
TASK_PP(16'h1B4FB,4);
TASK_PP(16'h1B4FC,4);
TASK_PP(16'h1B4FD,4);
TASK_PP(16'h1B4FE,4);
TASK_PP(16'h1B4FF,4);
TASK_PP(16'h1B500,4);
TASK_PP(16'h1B501,4);
TASK_PP(16'h1B502,4);
TASK_PP(16'h1B503,4);
TASK_PP(16'h1B504,4);
TASK_PP(16'h1B505,4);
TASK_PP(16'h1B506,4);
TASK_PP(16'h1B507,4);
TASK_PP(16'h1B508,4);
TASK_PP(16'h1B509,4);
TASK_PP(16'h1B50A,4);
TASK_PP(16'h1B50B,4);
TASK_PP(16'h1B50C,4);
TASK_PP(16'h1B50D,4);
TASK_PP(16'h1B50E,4);
TASK_PP(16'h1B50F,4);
TASK_PP(16'h1B510,4);
TASK_PP(16'h1B511,4);
TASK_PP(16'h1B512,4);
TASK_PP(16'h1B513,4);
TASK_PP(16'h1B514,4);
TASK_PP(16'h1B515,4);
TASK_PP(16'h1B516,4);
TASK_PP(16'h1B517,4);
TASK_PP(16'h1B518,4);
TASK_PP(16'h1B519,4);
TASK_PP(16'h1B51A,4);
TASK_PP(16'h1B51B,4);
TASK_PP(16'h1B51C,4);
TASK_PP(16'h1B51D,4);
TASK_PP(16'h1B51E,4);
TASK_PP(16'h1B51F,4);
TASK_PP(16'h1B520,4);
TASK_PP(16'h1B521,4);
TASK_PP(16'h1B522,4);
TASK_PP(16'h1B523,4);
TASK_PP(16'h1B524,4);
TASK_PP(16'h1B525,4);
TASK_PP(16'h1B526,4);
TASK_PP(16'h1B527,4);
TASK_PP(16'h1B528,4);
TASK_PP(16'h1B529,4);
TASK_PP(16'h1B52A,4);
TASK_PP(16'h1B52B,4);
TASK_PP(16'h1B52C,4);
TASK_PP(16'h1B52D,4);
TASK_PP(16'h1B52E,4);
TASK_PP(16'h1B52F,4);
TASK_PP(16'h1B530,4);
TASK_PP(16'h1B531,4);
TASK_PP(16'h1B532,4);
TASK_PP(16'h1B533,4);
TASK_PP(16'h1B534,4);
TASK_PP(16'h1B535,4);
TASK_PP(16'h1B536,4);
TASK_PP(16'h1B537,4);
TASK_PP(16'h1B538,4);
TASK_PP(16'h1B539,4);
TASK_PP(16'h1B53A,4);
TASK_PP(16'h1B53B,4);
TASK_PP(16'h1B53C,4);
TASK_PP(16'h1B53D,4);
TASK_PP(16'h1B53E,4);
TASK_PP(16'h1B53F,4);
TASK_PP(16'h1B540,4);
TASK_PP(16'h1B541,4);
TASK_PP(16'h1B542,4);
TASK_PP(16'h1B543,4);
TASK_PP(16'h1B544,4);
TASK_PP(16'h1B545,4);
TASK_PP(16'h1B546,4);
TASK_PP(16'h1B547,4);
TASK_PP(16'h1B548,4);
TASK_PP(16'h1B549,4);
TASK_PP(16'h1B54A,4);
TASK_PP(16'h1B54B,4);
TASK_PP(16'h1B54C,4);
TASK_PP(16'h1B54D,4);
TASK_PP(16'h1B54E,4);
TASK_PP(16'h1B54F,4);
TASK_PP(16'h1B550,4);
TASK_PP(16'h1B551,4);
TASK_PP(16'h1B552,4);
TASK_PP(16'h1B553,4);
TASK_PP(16'h1B554,4);
TASK_PP(16'h1B555,4);
TASK_PP(16'h1B556,4);
TASK_PP(16'h1B557,4);
TASK_PP(16'h1B558,4);
TASK_PP(16'h1B559,4);
TASK_PP(16'h1B55A,4);
TASK_PP(16'h1B55B,4);
TASK_PP(16'h1B55C,4);
TASK_PP(16'h1B55D,4);
TASK_PP(16'h1B55E,4);
TASK_PP(16'h1B55F,4);
TASK_PP(16'h1B560,4);
TASK_PP(16'h1B561,4);
TASK_PP(16'h1B562,4);
TASK_PP(16'h1B563,4);
TASK_PP(16'h1B564,4);
TASK_PP(16'h1B565,4);
TASK_PP(16'h1B566,4);
TASK_PP(16'h1B567,4);
TASK_PP(16'h1B568,4);
TASK_PP(16'h1B569,4);
TASK_PP(16'h1B56A,4);
TASK_PP(16'h1B56B,4);
TASK_PP(16'h1B56C,4);
TASK_PP(16'h1B56D,4);
TASK_PP(16'h1B56E,4);
TASK_PP(16'h1B56F,4);
TASK_PP(16'h1B570,4);
TASK_PP(16'h1B571,4);
TASK_PP(16'h1B572,4);
TASK_PP(16'h1B573,4);
TASK_PP(16'h1B574,4);
TASK_PP(16'h1B575,4);
TASK_PP(16'h1B576,4);
TASK_PP(16'h1B577,4);
TASK_PP(16'h1B578,4);
TASK_PP(16'h1B579,4);
TASK_PP(16'h1B57A,4);
TASK_PP(16'h1B57B,4);
TASK_PP(16'h1B57C,4);
TASK_PP(16'h1B57D,4);
TASK_PP(16'h1B57E,4);
TASK_PP(16'h1B57F,4);
TASK_PP(16'h1B580,4);
TASK_PP(16'h1B581,4);
TASK_PP(16'h1B582,4);
TASK_PP(16'h1B583,4);
TASK_PP(16'h1B584,4);
TASK_PP(16'h1B585,4);
TASK_PP(16'h1B586,4);
TASK_PP(16'h1B587,4);
TASK_PP(16'h1B588,4);
TASK_PP(16'h1B589,4);
TASK_PP(16'h1B58A,4);
TASK_PP(16'h1B58B,4);
TASK_PP(16'h1B58C,4);
TASK_PP(16'h1B58D,4);
TASK_PP(16'h1B58E,4);
TASK_PP(16'h1B58F,4);
TASK_PP(16'h1B590,4);
TASK_PP(16'h1B591,4);
TASK_PP(16'h1B592,4);
TASK_PP(16'h1B593,4);
TASK_PP(16'h1B594,4);
TASK_PP(16'h1B595,4);
TASK_PP(16'h1B596,4);
TASK_PP(16'h1B597,4);
TASK_PP(16'h1B598,4);
TASK_PP(16'h1B599,4);
TASK_PP(16'h1B59A,4);
TASK_PP(16'h1B59B,4);
TASK_PP(16'h1B59C,4);
TASK_PP(16'h1B59D,4);
TASK_PP(16'h1B59E,4);
TASK_PP(16'h1B59F,4);
TASK_PP(16'h1B5A0,4);
TASK_PP(16'h1B5A1,4);
TASK_PP(16'h1B5A2,4);
TASK_PP(16'h1B5A3,4);
TASK_PP(16'h1B5A4,4);
TASK_PP(16'h1B5A5,4);
TASK_PP(16'h1B5A6,4);
TASK_PP(16'h1B5A7,4);
TASK_PP(16'h1B5A8,4);
TASK_PP(16'h1B5A9,4);
TASK_PP(16'h1B5AA,4);
TASK_PP(16'h1B5AB,4);
TASK_PP(16'h1B5AC,4);
TASK_PP(16'h1B5AD,4);
TASK_PP(16'h1B5AE,4);
TASK_PP(16'h1B5AF,4);
TASK_PP(16'h1B5B0,4);
TASK_PP(16'h1B5B1,4);
TASK_PP(16'h1B5B2,4);
TASK_PP(16'h1B5B3,4);
TASK_PP(16'h1B5B4,4);
TASK_PP(16'h1B5B5,4);
TASK_PP(16'h1B5B6,4);
TASK_PP(16'h1B5B7,4);
TASK_PP(16'h1B5B8,4);
TASK_PP(16'h1B5B9,4);
TASK_PP(16'h1B5BA,4);
TASK_PP(16'h1B5BB,4);
TASK_PP(16'h1B5BC,4);
TASK_PP(16'h1B5BD,4);
TASK_PP(16'h1B5BE,4);
TASK_PP(16'h1B5BF,4);
TASK_PP(16'h1B5C0,4);
TASK_PP(16'h1B5C1,4);
TASK_PP(16'h1B5C2,4);
TASK_PP(16'h1B5C3,4);
TASK_PP(16'h1B5C4,4);
TASK_PP(16'h1B5C5,4);
TASK_PP(16'h1B5C6,4);
TASK_PP(16'h1B5C7,4);
TASK_PP(16'h1B5C8,4);
TASK_PP(16'h1B5C9,4);
TASK_PP(16'h1B5CA,4);
TASK_PP(16'h1B5CB,4);
TASK_PP(16'h1B5CC,4);
TASK_PP(16'h1B5CD,4);
TASK_PP(16'h1B5CE,4);
TASK_PP(16'h1B5CF,4);
TASK_PP(16'h1B5D0,4);
TASK_PP(16'h1B5D1,4);
TASK_PP(16'h1B5D2,4);
TASK_PP(16'h1B5D3,4);
TASK_PP(16'h1B5D4,4);
TASK_PP(16'h1B5D5,4);
TASK_PP(16'h1B5D6,4);
TASK_PP(16'h1B5D7,4);
TASK_PP(16'h1B5D8,4);
TASK_PP(16'h1B5D9,4);
TASK_PP(16'h1B5DA,4);
TASK_PP(16'h1B5DB,4);
TASK_PP(16'h1B5DC,4);
TASK_PP(16'h1B5DD,4);
TASK_PP(16'h1B5DE,4);
TASK_PP(16'h1B5DF,4);
TASK_PP(16'h1B5E0,4);
TASK_PP(16'h1B5E1,4);
TASK_PP(16'h1B5E2,4);
TASK_PP(16'h1B5E3,4);
TASK_PP(16'h1B5E4,4);
TASK_PP(16'h1B5E5,4);
TASK_PP(16'h1B5E6,4);
TASK_PP(16'h1B5E7,4);
TASK_PP(16'h1B5E8,4);
TASK_PP(16'h1B5E9,4);
TASK_PP(16'h1B5EA,4);
TASK_PP(16'h1B5EB,4);
TASK_PP(16'h1B5EC,4);
TASK_PP(16'h1B5ED,4);
TASK_PP(16'h1B5EE,4);
TASK_PP(16'h1B5EF,4);
TASK_PP(16'h1B5F0,4);
TASK_PP(16'h1B5F1,4);
TASK_PP(16'h1B5F2,4);
TASK_PP(16'h1B5F3,4);
TASK_PP(16'h1B5F4,4);
TASK_PP(16'h1B5F5,4);
TASK_PP(16'h1B5F6,4);
TASK_PP(16'h1B5F7,4);
TASK_PP(16'h1B5F8,4);
TASK_PP(16'h1B5F9,4);
TASK_PP(16'h1B5FA,4);
TASK_PP(16'h1B5FB,4);
TASK_PP(16'h1B5FC,4);
TASK_PP(16'h1B5FD,4);
TASK_PP(16'h1B5FE,4);
TASK_PP(16'h1B5FF,4);
TASK_PP(16'h1B600,4);
TASK_PP(16'h1B601,4);
TASK_PP(16'h1B602,4);
TASK_PP(16'h1B603,4);
TASK_PP(16'h1B604,4);
TASK_PP(16'h1B605,4);
TASK_PP(16'h1B606,4);
TASK_PP(16'h1B607,4);
TASK_PP(16'h1B608,4);
TASK_PP(16'h1B609,4);
TASK_PP(16'h1B60A,4);
TASK_PP(16'h1B60B,4);
TASK_PP(16'h1B60C,4);
TASK_PP(16'h1B60D,4);
TASK_PP(16'h1B60E,4);
TASK_PP(16'h1B60F,4);
TASK_PP(16'h1B610,4);
TASK_PP(16'h1B611,4);
TASK_PP(16'h1B612,4);
TASK_PP(16'h1B613,4);
TASK_PP(16'h1B614,4);
TASK_PP(16'h1B615,4);
TASK_PP(16'h1B616,4);
TASK_PP(16'h1B617,4);
TASK_PP(16'h1B618,4);
TASK_PP(16'h1B619,4);
TASK_PP(16'h1B61A,4);
TASK_PP(16'h1B61B,4);
TASK_PP(16'h1B61C,4);
TASK_PP(16'h1B61D,4);
TASK_PP(16'h1B61E,4);
TASK_PP(16'h1B61F,4);
TASK_PP(16'h1B620,4);
TASK_PP(16'h1B621,4);
TASK_PP(16'h1B622,4);
TASK_PP(16'h1B623,4);
TASK_PP(16'h1B624,4);
TASK_PP(16'h1B625,4);
TASK_PP(16'h1B626,4);
TASK_PP(16'h1B627,4);
TASK_PP(16'h1B628,4);
TASK_PP(16'h1B629,4);
TASK_PP(16'h1B62A,4);
TASK_PP(16'h1B62B,4);
TASK_PP(16'h1B62C,4);
TASK_PP(16'h1B62D,4);
TASK_PP(16'h1B62E,4);
TASK_PP(16'h1B62F,4);
TASK_PP(16'h1B630,4);
TASK_PP(16'h1B631,4);
TASK_PP(16'h1B632,4);
TASK_PP(16'h1B633,4);
TASK_PP(16'h1B634,4);
TASK_PP(16'h1B635,4);
TASK_PP(16'h1B636,4);
TASK_PP(16'h1B637,4);
TASK_PP(16'h1B638,4);
TASK_PP(16'h1B639,4);
TASK_PP(16'h1B63A,4);
TASK_PP(16'h1B63B,4);
TASK_PP(16'h1B63C,4);
TASK_PP(16'h1B63D,4);
TASK_PP(16'h1B63E,4);
TASK_PP(16'h1B63F,4);
TASK_PP(16'h1B640,4);
TASK_PP(16'h1B641,4);
TASK_PP(16'h1B642,4);
TASK_PP(16'h1B643,4);
TASK_PP(16'h1B644,4);
TASK_PP(16'h1B645,4);
TASK_PP(16'h1B646,4);
TASK_PP(16'h1B647,4);
TASK_PP(16'h1B648,4);
TASK_PP(16'h1B649,4);
TASK_PP(16'h1B64A,4);
TASK_PP(16'h1B64B,4);
TASK_PP(16'h1B64C,4);
TASK_PP(16'h1B64D,4);
TASK_PP(16'h1B64E,4);
TASK_PP(16'h1B64F,4);
TASK_PP(16'h1B650,4);
TASK_PP(16'h1B651,4);
TASK_PP(16'h1B652,4);
TASK_PP(16'h1B653,4);
TASK_PP(16'h1B654,4);
TASK_PP(16'h1B655,4);
TASK_PP(16'h1B656,4);
TASK_PP(16'h1B657,4);
TASK_PP(16'h1B658,4);
TASK_PP(16'h1B659,4);
TASK_PP(16'h1B65A,4);
TASK_PP(16'h1B65B,4);
TASK_PP(16'h1B65C,4);
TASK_PP(16'h1B65D,4);
TASK_PP(16'h1B65E,4);
TASK_PP(16'h1B65F,4);
TASK_PP(16'h1B660,4);
TASK_PP(16'h1B661,4);
TASK_PP(16'h1B662,4);
TASK_PP(16'h1B663,4);
TASK_PP(16'h1B664,4);
TASK_PP(16'h1B665,4);
TASK_PP(16'h1B666,4);
TASK_PP(16'h1B667,4);
TASK_PP(16'h1B668,4);
TASK_PP(16'h1B669,4);
TASK_PP(16'h1B66A,4);
TASK_PP(16'h1B66B,4);
TASK_PP(16'h1B66C,4);
TASK_PP(16'h1B66D,4);
TASK_PP(16'h1B66E,4);
TASK_PP(16'h1B66F,4);
TASK_PP(16'h1B670,4);
TASK_PP(16'h1B671,4);
TASK_PP(16'h1B672,4);
TASK_PP(16'h1B673,4);
TASK_PP(16'h1B674,4);
TASK_PP(16'h1B675,4);
TASK_PP(16'h1B676,4);
TASK_PP(16'h1B677,4);
TASK_PP(16'h1B678,4);
TASK_PP(16'h1B679,4);
TASK_PP(16'h1B67A,4);
TASK_PP(16'h1B67B,4);
TASK_PP(16'h1B67C,4);
TASK_PP(16'h1B67D,4);
TASK_PP(16'h1B67E,4);
TASK_PP(16'h1B67F,4);
TASK_PP(16'h1B680,4);
TASK_PP(16'h1B681,4);
TASK_PP(16'h1B682,4);
TASK_PP(16'h1B683,4);
TASK_PP(16'h1B684,4);
TASK_PP(16'h1B685,4);
TASK_PP(16'h1B686,4);
TASK_PP(16'h1B687,4);
TASK_PP(16'h1B688,4);
TASK_PP(16'h1B689,4);
TASK_PP(16'h1B68A,4);
TASK_PP(16'h1B68B,4);
TASK_PP(16'h1B68C,4);
TASK_PP(16'h1B68D,4);
TASK_PP(16'h1B68E,4);
TASK_PP(16'h1B68F,4);
TASK_PP(16'h1B690,4);
TASK_PP(16'h1B691,4);
TASK_PP(16'h1B692,4);
TASK_PP(16'h1B693,4);
TASK_PP(16'h1B694,4);
TASK_PP(16'h1B695,4);
TASK_PP(16'h1B696,4);
TASK_PP(16'h1B697,4);
TASK_PP(16'h1B698,4);
TASK_PP(16'h1B699,4);
TASK_PP(16'h1B69A,4);
TASK_PP(16'h1B69B,4);
TASK_PP(16'h1B69C,4);
TASK_PP(16'h1B69D,4);
TASK_PP(16'h1B69E,4);
TASK_PP(16'h1B69F,4);
TASK_PP(16'h1B6A0,4);
TASK_PP(16'h1B6A1,4);
TASK_PP(16'h1B6A2,4);
TASK_PP(16'h1B6A3,4);
TASK_PP(16'h1B6A4,4);
TASK_PP(16'h1B6A5,4);
TASK_PP(16'h1B6A6,4);
TASK_PP(16'h1B6A7,4);
TASK_PP(16'h1B6A8,4);
TASK_PP(16'h1B6A9,4);
TASK_PP(16'h1B6AA,4);
TASK_PP(16'h1B6AB,4);
TASK_PP(16'h1B6AC,4);
TASK_PP(16'h1B6AD,4);
TASK_PP(16'h1B6AE,4);
TASK_PP(16'h1B6AF,4);
TASK_PP(16'h1B6B0,4);
TASK_PP(16'h1B6B1,4);
TASK_PP(16'h1B6B2,4);
TASK_PP(16'h1B6B3,4);
TASK_PP(16'h1B6B4,4);
TASK_PP(16'h1B6B5,4);
TASK_PP(16'h1B6B6,4);
TASK_PP(16'h1B6B7,4);
TASK_PP(16'h1B6B8,4);
TASK_PP(16'h1B6B9,4);
TASK_PP(16'h1B6BA,4);
TASK_PP(16'h1B6BB,4);
TASK_PP(16'h1B6BC,4);
TASK_PP(16'h1B6BD,4);
TASK_PP(16'h1B6BE,4);
TASK_PP(16'h1B6BF,4);
TASK_PP(16'h1B6C0,4);
TASK_PP(16'h1B6C1,4);
TASK_PP(16'h1B6C2,4);
TASK_PP(16'h1B6C3,4);
TASK_PP(16'h1B6C4,4);
TASK_PP(16'h1B6C5,4);
TASK_PP(16'h1B6C6,4);
TASK_PP(16'h1B6C7,4);
TASK_PP(16'h1B6C8,4);
TASK_PP(16'h1B6C9,4);
TASK_PP(16'h1B6CA,4);
TASK_PP(16'h1B6CB,4);
TASK_PP(16'h1B6CC,4);
TASK_PP(16'h1B6CD,4);
TASK_PP(16'h1B6CE,4);
TASK_PP(16'h1B6CF,4);
TASK_PP(16'h1B6D0,4);
TASK_PP(16'h1B6D1,4);
TASK_PP(16'h1B6D2,4);
TASK_PP(16'h1B6D3,4);
TASK_PP(16'h1B6D4,4);
TASK_PP(16'h1B6D5,4);
TASK_PP(16'h1B6D6,4);
TASK_PP(16'h1B6D7,4);
TASK_PP(16'h1B6D8,4);
TASK_PP(16'h1B6D9,4);
TASK_PP(16'h1B6DA,4);
TASK_PP(16'h1B6DB,4);
TASK_PP(16'h1B6DC,4);
TASK_PP(16'h1B6DD,4);
TASK_PP(16'h1B6DE,4);
TASK_PP(16'h1B6DF,4);
TASK_PP(16'h1B6E0,4);
TASK_PP(16'h1B6E1,4);
TASK_PP(16'h1B6E2,4);
TASK_PP(16'h1B6E3,4);
TASK_PP(16'h1B6E4,4);
TASK_PP(16'h1B6E5,4);
TASK_PP(16'h1B6E6,4);
TASK_PP(16'h1B6E7,4);
TASK_PP(16'h1B6E8,4);
TASK_PP(16'h1B6E9,4);
TASK_PP(16'h1B6EA,4);
TASK_PP(16'h1B6EB,4);
TASK_PP(16'h1B6EC,4);
TASK_PP(16'h1B6ED,4);
TASK_PP(16'h1B6EE,4);
TASK_PP(16'h1B6EF,4);
TASK_PP(16'h1B6F0,4);
TASK_PP(16'h1B6F1,4);
TASK_PP(16'h1B6F2,4);
TASK_PP(16'h1B6F3,4);
TASK_PP(16'h1B6F4,4);
TASK_PP(16'h1B6F5,4);
TASK_PP(16'h1B6F6,4);
TASK_PP(16'h1B6F7,4);
TASK_PP(16'h1B6F8,4);
TASK_PP(16'h1B6F9,4);
TASK_PP(16'h1B6FA,4);
TASK_PP(16'h1B6FB,4);
TASK_PP(16'h1B6FC,4);
TASK_PP(16'h1B6FD,4);
TASK_PP(16'h1B6FE,4);
TASK_PP(16'h1B6FF,4);
TASK_PP(16'h1B700,4);
TASK_PP(16'h1B701,4);
TASK_PP(16'h1B702,4);
TASK_PP(16'h1B703,4);
TASK_PP(16'h1B704,4);
TASK_PP(16'h1B705,4);
TASK_PP(16'h1B706,4);
TASK_PP(16'h1B707,4);
TASK_PP(16'h1B708,4);
TASK_PP(16'h1B709,4);
TASK_PP(16'h1B70A,4);
TASK_PP(16'h1B70B,4);
TASK_PP(16'h1B70C,4);
TASK_PP(16'h1B70D,4);
TASK_PP(16'h1B70E,4);
TASK_PP(16'h1B70F,4);
TASK_PP(16'h1B710,4);
TASK_PP(16'h1B711,4);
TASK_PP(16'h1B712,4);
TASK_PP(16'h1B713,4);
TASK_PP(16'h1B714,4);
TASK_PP(16'h1B715,4);
TASK_PP(16'h1B716,4);
TASK_PP(16'h1B717,4);
TASK_PP(16'h1B718,4);
TASK_PP(16'h1B719,4);
TASK_PP(16'h1B71A,4);
TASK_PP(16'h1B71B,4);
TASK_PP(16'h1B71C,4);
TASK_PP(16'h1B71D,4);
TASK_PP(16'h1B71E,4);
TASK_PP(16'h1B71F,4);
TASK_PP(16'h1B720,4);
TASK_PP(16'h1B721,4);
TASK_PP(16'h1B722,4);
TASK_PP(16'h1B723,4);
TASK_PP(16'h1B724,4);
TASK_PP(16'h1B725,4);
TASK_PP(16'h1B726,4);
TASK_PP(16'h1B727,4);
TASK_PP(16'h1B728,4);
TASK_PP(16'h1B729,4);
TASK_PP(16'h1B72A,4);
TASK_PP(16'h1B72B,4);
TASK_PP(16'h1B72C,4);
TASK_PP(16'h1B72D,4);
TASK_PP(16'h1B72E,4);
TASK_PP(16'h1B72F,4);
TASK_PP(16'h1B730,4);
TASK_PP(16'h1B731,4);
TASK_PP(16'h1B732,4);
TASK_PP(16'h1B733,4);
TASK_PP(16'h1B734,4);
TASK_PP(16'h1B735,4);
TASK_PP(16'h1B736,4);
TASK_PP(16'h1B737,4);
TASK_PP(16'h1B738,4);
TASK_PP(16'h1B739,4);
TASK_PP(16'h1B73A,4);
TASK_PP(16'h1B73B,4);
TASK_PP(16'h1B73C,4);
TASK_PP(16'h1B73D,4);
TASK_PP(16'h1B73E,4);
TASK_PP(16'h1B73F,4);
TASK_PP(16'h1B740,4);
TASK_PP(16'h1B741,4);
TASK_PP(16'h1B742,4);
TASK_PP(16'h1B743,4);
TASK_PP(16'h1B744,4);
TASK_PP(16'h1B745,4);
TASK_PP(16'h1B746,4);
TASK_PP(16'h1B747,4);
TASK_PP(16'h1B748,4);
TASK_PP(16'h1B749,4);
TASK_PP(16'h1B74A,4);
TASK_PP(16'h1B74B,4);
TASK_PP(16'h1B74C,4);
TASK_PP(16'h1B74D,4);
TASK_PP(16'h1B74E,4);
TASK_PP(16'h1B74F,4);
TASK_PP(16'h1B750,4);
TASK_PP(16'h1B751,4);
TASK_PP(16'h1B752,4);
TASK_PP(16'h1B753,4);
TASK_PP(16'h1B754,4);
TASK_PP(16'h1B755,4);
TASK_PP(16'h1B756,4);
TASK_PP(16'h1B757,4);
TASK_PP(16'h1B758,4);
TASK_PP(16'h1B759,4);
TASK_PP(16'h1B75A,4);
TASK_PP(16'h1B75B,4);
TASK_PP(16'h1B75C,4);
TASK_PP(16'h1B75D,4);
TASK_PP(16'h1B75E,4);
TASK_PP(16'h1B75F,4);
TASK_PP(16'h1B760,4);
TASK_PP(16'h1B761,4);
TASK_PP(16'h1B762,4);
TASK_PP(16'h1B763,4);
TASK_PP(16'h1B764,4);
TASK_PP(16'h1B765,4);
TASK_PP(16'h1B766,4);
TASK_PP(16'h1B767,4);
TASK_PP(16'h1B768,4);
TASK_PP(16'h1B769,4);
TASK_PP(16'h1B76A,4);
TASK_PP(16'h1B76B,4);
TASK_PP(16'h1B76C,4);
TASK_PP(16'h1B76D,4);
TASK_PP(16'h1B76E,4);
TASK_PP(16'h1B76F,4);
TASK_PP(16'h1B770,4);
TASK_PP(16'h1B771,4);
TASK_PP(16'h1B772,4);
TASK_PP(16'h1B773,4);
TASK_PP(16'h1B774,4);
TASK_PP(16'h1B775,4);
TASK_PP(16'h1B776,4);
TASK_PP(16'h1B777,4);
TASK_PP(16'h1B778,4);
TASK_PP(16'h1B779,4);
TASK_PP(16'h1B77A,4);
TASK_PP(16'h1B77B,4);
TASK_PP(16'h1B77C,4);
TASK_PP(16'h1B77D,4);
TASK_PP(16'h1B77E,4);
TASK_PP(16'h1B77F,4);
TASK_PP(16'h1B780,4);
TASK_PP(16'h1B781,4);
TASK_PP(16'h1B782,4);
TASK_PP(16'h1B783,4);
TASK_PP(16'h1B784,4);
TASK_PP(16'h1B785,4);
TASK_PP(16'h1B786,4);
TASK_PP(16'h1B787,4);
TASK_PP(16'h1B788,4);
TASK_PP(16'h1B789,4);
TASK_PP(16'h1B78A,4);
TASK_PP(16'h1B78B,4);
TASK_PP(16'h1B78C,4);
TASK_PP(16'h1B78D,4);
TASK_PP(16'h1B78E,4);
TASK_PP(16'h1B78F,4);
TASK_PP(16'h1B790,4);
TASK_PP(16'h1B791,4);
TASK_PP(16'h1B792,4);
TASK_PP(16'h1B793,4);
TASK_PP(16'h1B794,4);
TASK_PP(16'h1B795,4);
TASK_PP(16'h1B796,4);
TASK_PP(16'h1B797,4);
TASK_PP(16'h1B798,4);
TASK_PP(16'h1B799,4);
TASK_PP(16'h1B79A,4);
TASK_PP(16'h1B79B,4);
TASK_PP(16'h1B79C,4);
TASK_PP(16'h1B79D,4);
TASK_PP(16'h1B79E,4);
TASK_PP(16'h1B79F,4);
TASK_PP(16'h1B7A0,4);
TASK_PP(16'h1B7A1,4);
TASK_PP(16'h1B7A2,4);
TASK_PP(16'h1B7A3,4);
TASK_PP(16'h1B7A4,4);
TASK_PP(16'h1B7A5,4);
TASK_PP(16'h1B7A6,4);
TASK_PP(16'h1B7A7,4);
TASK_PP(16'h1B7A8,4);
TASK_PP(16'h1B7A9,4);
TASK_PP(16'h1B7AA,4);
TASK_PP(16'h1B7AB,4);
TASK_PP(16'h1B7AC,4);
TASK_PP(16'h1B7AD,4);
TASK_PP(16'h1B7AE,4);
TASK_PP(16'h1B7AF,4);
TASK_PP(16'h1B7B0,4);
TASK_PP(16'h1B7B1,4);
TASK_PP(16'h1B7B2,4);
TASK_PP(16'h1B7B3,4);
TASK_PP(16'h1B7B4,4);
TASK_PP(16'h1B7B5,4);
TASK_PP(16'h1B7B6,4);
TASK_PP(16'h1B7B7,4);
TASK_PP(16'h1B7B8,4);
TASK_PP(16'h1B7B9,4);
TASK_PP(16'h1B7BA,4);
TASK_PP(16'h1B7BB,4);
TASK_PP(16'h1B7BC,4);
TASK_PP(16'h1B7BD,4);
TASK_PP(16'h1B7BE,4);
TASK_PP(16'h1B7BF,4);
TASK_PP(16'h1B7C0,4);
TASK_PP(16'h1B7C1,4);
TASK_PP(16'h1B7C2,4);
TASK_PP(16'h1B7C3,4);
TASK_PP(16'h1B7C4,4);
TASK_PP(16'h1B7C5,4);
TASK_PP(16'h1B7C6,4);
TASK_PP(16'h1B7C7,4);
TASK_PP(16'h1B7C8,4);
TASK_PP(16'h1B7C9,4);
TASK_PP(16'h1B7CA,4);
TASK_PP(16'h1B7CB,4);
TASK_PP(16'h1B7CC,4);
TASK_PP(16'h1B7CD,4);
TASK_PP(16'h1B7CE,4);
TASK_PP(16'h1B7CF,4);
TASK_PP(16'h1B7D0,4);
TASK_PP(16'h1B7D1,4);
TASK_PP(16'h1B7D2,4);
TASK_PP(16'h1B7D3,4);
TASK_PP(16'h1B7D4,4);
TASK_PP(16'h1B7D5,4);
TASK_PP(16'h1B7D6,4);
TASK_PP(16'h1B7D7,4);
TASK_PP(16'h1B7D8,4);
TASK_PP(16'h1B7D9,4);
TASK_PP(16'h1B7DA,4);
TASK_PP(16'h1B7DB,4);
TASK_PP(16'h1B7DC,4);
TASK_PP(16'h1B7DD,4);
TASK_PP(16'h1B7DE,4);
TASK_PP(16'h1B7DF,4);
TASK_PP(16'h1B7E0,4);
TASK_PP(16'h1B7E1,4);
TASK_PP(16'h1B7E2,4);
TASK_PP(16'h1B7E3,4);
TASK_PP(16'h1B7E4,4);
TASK_PP(16'h1B7E5,4);
TASK_PP(16'h1B7E6,4);
TASK_PP(16'h1B7E7,4);
TASK_PP(16'h1B7E8,4);
TASK_PP(16'h1B7E9,4);
TASK_PP(16'h1B7EA,4);
TASK_PP(16'h1B7EB,4);
TASK_PP(16'h1B7EC,4);
TASK_PP(16'h1B7ED,4);
TASK_PP(16'h1B7EE,4);
TASK_PP(16'h1B7EF,4);
TASK_PP(16'h1B7F0,4);
TASK_PP(16'h1B7F1,4);
TASK_PP(16'h1B7F2,4);
TASK_PP(16'h1B7F3,4);
TASK_PP(16'h1B7F4,4);
TASK_PP(16'h1B7F5,4);
TASK_PP(16'h1B7F6,4);
TASK_PP(16'h1B7F7,4);
TASK_PP(16'h1B7F8,4);
TASK_PP(16'h1B7F9,4);
TASK_PP(16'h1B7FA,4);
TASK_PP(16'h1B7FB,4);
TASK_PP(16'h1B7FC,4);
TASK_PP(16'h1B7FD,4);
TASK_PP(16'h1B7FE,4);
TASK_PP(16'h1B7FF,4);
TASK_PP(16'h1B800,4);
TASK_PP(16'h1B801,4);
TASK_PP(16'h1B802,4);
TASK_PP(16'h1B803,4);
TASK_PP(16'h1B804,4);
TASK_PP(16'h1B805,4);
TASK_PP(16'h1B806,4);
TASK_PP(16'h1B807,4);
TASK_PP(16'h1B808,4);
TASK_PP(16'h1B809,4);
TASK_PP(16'h1B80A,4);
TASK_PP(16'h1B80B,4);
TASK_PP(16'h1B80C,4);
TASK_PP(16'h1B80D,4);
TASK_PP(16'h1B80E,4);
TASK_PP(16'h1B80F,4);
TASK_PP(16'h1B810,4);
TASK_PP(16'h1B811,4);
TASK_PP(16'h1B812,4);
TASK_PP(16'h1B813,4);
TASK_PP(16'h1B814,4);
TASK_PP(16'h1B815,4);
TASK_PP(16'h1B816,4);
TASK_PP(16'h1B817,4);
TASK_PP(16'h1B818,4);
TASK_PP(16'h1B819,4);
TASK_PP(16'h1B81A,4);
TASK_PP(16'h1B81B,4);
TASK_PP(16'h1B81C,4);
TASK_PP(16'h1B81D,4);
TASK_PP(16'h1B81E,4);
TASK_PP(16'h1B81F,4);
TASK_PP(16'h1B820,4);
TASK_PP(16'h1B821,4);
TASK_PP(16'h1B822,4);
TASK_PP(16'h1B823,4);
TASK_PP(16'h1B824,4);
TASK_PP(16'h1B825,4);
TASK_PP(16'h1B826,4);
TASK_PP(16'h1B827,4);
TASK_PP(16'h1B828,4);
TASK_PP(16'h1B829,4);
TASK_PP(16'h1B82A,4);
TASK_PP(16'h1B82B,4);
TASK_PP(16'h1B82C,4);
TASK_PP(16'h1B82D,4);
TASK_PP(16'h1B82E,4);
TASK_PP(16'h1B82F,4);
TASK_PP(16'h1B830,4);
TASK_PP(16'h1B831,4);
TASK_PP(16'h1B832,4);
TASK_PP(16'h1B833,4);
TASK_PP(16'h1B834,4);
TASK_PP(16'h1B835,4);
TASK_PP(16'h1B836,4);
TASK_PP(16'h1B837,4);
TASK_PP(16'h1B838,4);
TASK_PP(16'h1B839,4);
TASK_PP(16'h1B83A,4);
TASK_PP(16'h1B83B,4);
TASK_PP(16'h1B83C,4);
TASK_PP(16'h1B83D,4);
TASK_PP(16'h1B83E,4);
TASK_PP(16'h1B83F,4);
TASK_PP(16'h1B840,4);
TASK_PP(16'h1B841,4);
TASK_PP(16'h1B842,4);
TASK_PP(16'h1B843,4);
TASK_PP(16'h1B844,4);
TASK_PP(16'h1B845,4);
TASK_PP(16'h1B846,4);
TASK_PP(16'h1B847,4);
TASK_PP(16'h1B848,4);
TASK_PP(16'h1B849,4);
TASK_PP(16'h1B84A,4);
TASK_PP(16'h1B84B,4);
TASK_PP(16'h1B84C,4);
TASK_PP(16'h1B84D,4);
TASK_PP(16'h1B84E,4);
TASK_PP(16'h1B84F,4);
TASK_PP(16'h1B850,4);
TASK_PP(16'h1B851,4);
TASK_PP(16'h1B852,4);
TASK_PP(16'h1B853,4);
TASK_PP(16'h1B854,4);
TASK_PP(16'h1B855,4);
TASK_PP(16'h1B856,4);
TASK_PP(16'h1B857,4);
TASK_PP(16'h1B858,4);
TASK_PP(16'h1B859,4);
TASK_PP(16'h1B85A,4);
TASK_PP(16'h1B85B,4);
TASK_PP(16'h1B85C,4);
TASK_PP(16'h1B85D,4);
TASK_PP(16'h1B85E,4);
TASK_PP(16'h1B85F,4);
TASK_PP(16'h1B860,4);
TASK_PP(16'h1B861,4);
TASK_PP(16'h1B862,4);
TASK_PP(16'h1B863,4);
TASK_PP(16'h1B864,4);
TASK_PP(16'h1B865,4);
TASK_PP(16'h1B866,4);
TASK_PP(16'h1B867,4);
TASK_PP(16'h1B868,4);
TASK_PP(16'h1B869,4);
TASK_PP(16'h1B86A,4);
TASK_PP(16'h1B86B,4);
TASK_PP(16'h1B86C,4);
TASK_PP(16'h1B86D,4);
TASK_PP(16'h1B86E,4);
TASK_PP(16'h1B86F,4);
TASK_PP(16'h1B870,4);
TASK_PP(16'h1B871,4);
TASK_PP(16'h1B872,4);
TASK_PP(16'h1B873,4);
TASK_PP(16'h1B874,4);
TASK_PP(16'h1B875,4);
TASK_PP(16'h1B876,4);
TASK_PP(16'h1B877,4);
TASK_PP(16'h1B878,4);
TASK_PP(16'h1B879,4);
TASK_PP(16'h1B87A,4);
TASK_PP(16'h1B87B,4);
TASK_PP(16'h1B87C,4);
TASK_PP(16'h1B87D,4);
TASK_PP(16'h1B87E,4);
TASK_PP(16'h1B87F,4);
TASK_PP(16'h1B880,4);
TASK_PP(16'h1B881,4);
TASK_PP(16'h1B882,4);
TASK_PP(16'h1B883,4);
TASK_PP(16'h1B884,4);
TASK_PP(16'h1B885,4);
TASK_PP(16'h1B886,4);
TASK_PP(16'h1B887,4);
TASK_PP(16'h1B888,4);
TASK_PP(16'h1B889,4);
TASK_PP(16'h1B88A,4);
TASK_PP(16'h1B88B,4);
TASK_PP(16'h1B88C,4);
TASK_PP(16'h1B88D,4);
TASK_PP(16'h1B88E,4);
TASK_PP(16'h1B88F,4);
TASK_PP(16'h1B890,4);
TASK_PP(16'h1B891,4);
TASK_PP(16'h1B892,4);
TASK_PP(16'h1B893,4);
TASK_PP(16'h1B894,4);
TASK_PP(16'h1B895,4);
TASK_PP(16'h1B896,4);
TASK_PP(16'h1B897,4);
TASK_PP(16'h1B898,4);
TASK_PP(16'h1B899,4);
TASK_PP(16'h1B89A,4);
TASK_PP(16'h1B89B,4);
TASK_PP(16'h1B89C,4);
TASK_PP(16'h1B89D,4);
TASK_PP(16'h1B89E,4);
TASK_PP(16'h1B89F,4);
TASK_PP(16'h1B8A0,4);
TASK_PP(16'h1B8A1,4);
TASK_PP(16'h1B8A2,4);
TASK_PP(16'h1B8A3,4);
TASK_PP(16'h1B8A4,4);
TASK_PP(16'h1B8A5,4);
TASK_PP(16'h1B8A6,4);
TASK_PP(16'h1B8A7,4);
TASK_PP(16'h1B8A8,4);
TASK_PP(16'h1B8A9,4);
TASK_PP(16'h1B8AA,4);
TASK_PP(16'h1B8AB,4);
TASK_PP(16'h1B8AC,4);
TASK_PP(16'h1B8AD,4);
TASK_PP(16'h1B8AE,4);
TASK_PP(16'h1B8AF,4);
TASK_PP(16'h1B8B0,4);
TASK_PP(16'h1B8B1,4);
TASK_PP(16'h1B8B2,4);
TASK_PP(16'h1B8B3,4);
TASK_PP(16'h1B8B4,4);
TASK_PP(16'h1B8B5,4);
TASK_PP(16'h1B8B6,4);
TASK_PP(16'h1B8B7,4);
TASK_PP(16'h1B8B8,4);
TASK_PP(16'h1B8B9,4);
TASK_PP(16'h1B8BA,4);
TASK_PP(16'h1B8BB,4);
TASK_PP(16'h1B8BC,4);
TASK_PP(16'h1B8BD,4);
TASK_PP(16'h1B8BE,4);
TASK_PP(16'h1B8BF,4);
TASK_PP(16'h1B8C0,4);
TASK_PP(16'h1B8C1,4);
TASK_PP(16'h1B8C2,4);
TASK_PP(16'h1B8C3,4);
TASK_PP(16'h1B8C4,4);
TASK_PP(16'h1B8C5,4);
TASK_PP(16'h1B8C6,4);
TASK_PP(16'h1B8C7,4);
TASK_PP(16'h1B8C8,4);
TASK_PP(16'h1B8C9,4);
TASK_PP(16'h1B8CA,4);
TASK_PP(16'h1B8CB,4);
TASK_PP(16'h1B8CC,4);
TASK_PP(16'h1B8CD,4);
TASK_PP(16'h1B8CE,4);
TASK_PP(16'h1B8CF,4);
TASK_PP(16'h1B8D0,4);
TASK_PP(16'h1B8D1,4);
TASK_PP(16'h1B8D2,4);
TASK_PP(16'h1B8D3,4);
TASK_PP(16'h1B8D4,4);
TASK_PP(16'h1B8D5,4);
TASK_PP(16'h1B8D6,4);
TASK_PP(16'h1B8D7,4);
TASK_PP(16'h1B8D8,4);
TASK_PP(16'h1B8D9,4);
TASK_PP(16'h1B8DA,4);
TASK_PP(16'h1B8DB,4);
TASK_PP(16'h1B8DC,4);
TASK_PP(16'h1B8DD,4);
TASK_PP(16'h1B8DE,4);
TASK_PP(16'h1B8DF,4);
TASK_PP(16'h1B8E0,4);
TASK_PP(16'h1B8E1,4);
TASK_PP(16'h1B8E2,4);
TASK_PP(16'h1B8E3,4);
TASK_PP(16'h1B8E4,4);
TASK_PP(16'h1B8E5,4);
TASK_PP(16'h1B8E6,4);
TASK_PP(16'h1B8E7,4);
TASK_PP(16'h1B8E8,4);
TASK_PP(16'h1B8E9,4);
TASK_PP(16'h1B8EA,4);
TASK_PP(16'h1B8EB,4);
TASK_PP(16'h1B8EC,4);
TASK_PP(16'h1B8ED,4);
TASK_PP(16'h1B8EE,4);
TASK_PP(16'h1B8EF,4);
TASK_PP(16'h1B8F0,4);
TASK_PP(16'h1B8F1,4);
TASK_PP(16'h1B8F2,4);
TASK_PP(16'h1B8F3,4);
TASK_PP(16'h1B8F4,4);
TASK_PP(16'h1B8F5,4);
TASK_PP(16'h1B8F6,4);
TASK_PP(16'h1B8F7,4);
TASK_PP(16'h1B8F8,4);
TASK_PP(16'h1B8F9,4);
TASK_PP(16'h1B8FA,4);
TASK_PP(16'h1B8FB,4);
TASK_PP(16'h1B8FC,4);
TASK_PP(16'h1B8FD,4);
TASK_PP(16'h1B8FE,4);
TASK_PP(16'h1B8FF,4);
TASK_PP(16'h1B900,4);
TASK_PP(16'h1B901,4);
TASK_PP(16'h1B902,4);
TASK_PP(16'h1B903,4);
TASK_PP(16'h1B904,4);
TASK_PP(16'h1B905,4);
TASK_PP(16'h1B906,4);
TASK_PP(16'h1B907,4);
TASK_PP(16'h1B908,4);
TASK_PP(16'h1B909,4);
TASK_PP(16'h1B90A,4);
TASK_PP(16'h1B90B,4);
TASK_PP(16'h1B90C,4);
TASK_PP(16'h1B90D,4);
TASK_PP(16'h1B90E,4);
TASK_PP(16'h1B90F,4);
TASK_PP(16'h1B910,4);
TASK_PP(16'h1B911,4);
TASK_PP(16'h1B912,4);
TASK_PP(16'h1B913,4);
TASK_PP(16'h1B914,4);
TASK_PP(16'h1B915,4);
TASK_PP(16'h1B916,4);
TASK_PP(16'h1B917,4);
TASK_PP(16'h1B918,4);
TASK_PP(16'h1B919,4);
TASK_PP(16'h1B91A,4);
TASK_PP(16'h1B91B,4);
TASK_PP(16'h1B91C,4);
TASK_PP(16'h1B91D,4);
TASK_PP(16'h1B91E,4);
TASK_PP(16'h1B91F,4);
TASK_PP(16'h1B920,4);
TASK_PP(16'h1B921,4);
TASK_PP(16'h1B922,4);
TASK_PP(16'h1B923,4);
TASK_PP(16'h1B924,4);
TASK_PP(16'h1B925,4);
TASK_PP(16'h1B926,4);
TASK_PP(16'h1B927,4);
TASK_PP(16'h1B928,4);
TASK_PP(16'h1B929,4);
TASK_PP(16'h1B92A,4);
TASK_PP(16'h1B92B,4);
TASK_PP(16'h1B92C,4);
TASK_PP(16'h1B92D,4);
TASK_PP(16'h1B92E,4);
TASK_PP(16'h1B92F,4);
TASK_PP(16'h1B930,4);
TASK_PP(16'h1B931,4);
TASK_PP(16'h1B932,4);
TASK_PP(16'h1B933,4);
TASK_PP(16'h1B934,4);
TASK_PP(16'h1B935,4);
TASK_PP(16'h1B936,4);
TASK_PP(16'h1B937,4);
TASK_PP(16'h1B938,4);
TASK_PP(16'h1B939,4);
TASK_PP(16'h1B93A,4);
TASK_PP(16'h1B93B,4);
TASK_PP(16'h1B93C,4);
TASK_PP(16'h1B93D,4);
TASK_PP(16'h1B93E,4);
TASK_PP(16'h1B93F,4);
TASK_PP(16'h1B940,4);
TASK_PP(16'h1B941,4);
TASK_PP(16'h1B942,4);
TASK_PP(16'h1B943,4);
TASK_PP(16'h1B944,4);
TASK_PP(16'h1B945,4);
TASK_PP(16'h1B946,4);
TASK_PP(16'h1B947,4);
TASK_PP(16'h1B948,4);
TASK_PP(16'h1B949,4);
TASK_PP(16'h1B94A,4);
TASK_PP(16'h1B94B,4);
TASK_PP(16'h1B94C,4);
TASK_PP(16'h1B94D,4);
TASK_PP(16'h1B94E,4);
TASK_PP(16'h1B94F,4);
TASK_PP(16'h1B950,4);
TASK_PP(16'h1B951,4);
TASK_PP(16'h1B952,4);
TASK_PP(16'h1B953,4);
TASK_PP(16'h1B954,4);
TASK_PP(16'h1B955,4);
TASK_PP(16'h1B956,4);
TASK_PP(16'h1B957,4);
TASK_PP(16'h1B958,4);
TASK_PP(16'h1B959,4);
TASK_PP(16'h1B95A,4);
TASK_PP(16'h1B95B,4);
TASK_PP(16'h1B95C,4);
TASK_PP(16'h1B95D,4);
TASK_PP(16'h1B95E,4);
TASK_PP(16'h1B95F,4);
TASK_PP(16'h1B960,4);
TASK_PP(16'h1B961,4);
TASK_PP(16'h1B962,4);
TASK_PP(16'h1B963,4);
TASK_PP(16'h1B964,4);
TASK_PP(16'h1B965,4);
TASK_PP(16'h1B966,4);
TASK_PP(16'h1B967,4);
TASK_PP(16'h1B968,4);
TASK_PP(16'h1B969,4);
TASK_PP(16'h1B96A,4);
TASK_PP(16'h1B96B,4);
TASK_PP(16'h1B96C,4);
TASK_PP(16'h1B96D,4);
TASK_PP(16'h1B96E,4);
TASK_PP(16'h1B96F,4);
TASK_PP(16'h1B970,4);
TASK_PP(16'h1B971,4);
TASK_PP(16'h1B972,4);
TASK_PP(16'h1B973,4);
TASK_PP(16'h1B974,4);
TASK_PP(16'h1B975,4);
TASK_PP(16'h1B976,4);
TASK_PP(16'h1B977,4);
TASK_PP(16'h1B978,4);
TASK_PP(16'h1B979,4);
TASK_PP(16'h1B97A,4);
TASK_PP(16'h1B97B,4);
TASK_PP(16'h1B97C,4);
TASK_PP(16'h1B97D,4);
TASK_PP(16'h1B97E,4);
TASK_PP(16'h1B97F,4);
TASK_PP(16'h1B980,4);
TASK_PP(16'h1B981,4);
TASK_PP(16'h1B982,4);
TASK_PP(16'h1B983,4);
TASK_PP(16'h1B984,4);
TASK_PP(16'h1B985,4);
TASK_PP(16'h1B986,4);
TASK_PP(16'h1B987,4);
TASK_PP(16'h1B988,4);
TASK_PP(16'h1B989,4);
TASK_PP(16'h1B98A,4);
TASK_PP(16'h1B98B,4);
TASK_PP(16'h1B98C,4);
TASK_PP(16'h1B98D,4);
TASK_PP(16'h1B98E,4);
TASK_PP(16'h1B98F,4);
TASK_PP(16'h1B990,4);
TASK_PP(16'h1B991,4);
TASK_PP(16'h1B992,4);
TASK_PP(16'h1B993,4);
TASK_PP(16'h1B994,4);
TASK_PP(16'h1B995,4);
TASK_PP(16'h1B996,4);
TASK_PP(16'h1B997,4);
TASK_PP(16'h1B998,4);
TASK_PP(16'h1B999,4);
TASK_PP(16'h1B99A,4);
TASK_PP(16'h1B99B,4);
TASK_PP(16'h1B99C,4);
TASK_PP(16'h1B99D,4);
TASK_PP(16'h1B99E,4);
TASK_PP(16'h1B99F,4);
TASK_PP(16'h1B9A0,4);
TASK_PP(16'h1B9A1,4);
TASK_PP(16'h1B9A2,4);
TASK_PP(16'h1B9A3,4);
TASK_PP(16'h1B9A4,4);
TASK_PP(16'h1B9A5,4);
TASK_PP(16'h1B9A6,4);
TASK_PP(16'h1B9A7,4);
TASK_PP(16'h1B9A8,4);
TASK_PP(16'h1B9A9,4);
TASK_PP(16'h1B9AA,4);
TASK_PP(16'h1B9AB,4);
TASK_PP(16'h1B9AC,4);
TASK_PP(16'h1B9AD,4);
TASK_PP(16'h1B9AE,4);
TASK_PP(16'h1B9AF,4);
TASK_PP(16'h1B9B0,4);
TASK_PP(16'h1B9B1,4);
TASK_PP(16'h1B9B2,4);
TASK_PP(16'h1B9B3,4);
TASK_PP(16'h1B9B4,4);
TASK_PP(16'h1B9B5,4);
TASK_PP(16'h1B9B6,4);
TASK_PP(16'h1B9B7,4);
TASK_PP(16'h1B9B8,4);
TASK_PP(16'h1B9B9,4);
TASK_PP(16'h1B9BA,4);
TASK_PP(16'h1B9BB,4);
TASK_PP(16'h1B9BC,4);
TASK_PP(16'h1B9BD,4);
TASK_PP(16'h1B9BE,4);
TASK_PP(16'h1B9BF,4);
TASK_PP(16'h1B9C0,4);
TASK_PP(16'h1B9C1,4);
TASK_PP(16'h1B9C2,4);
TASK_PP(16'h1B9C3,4);
TASK_PP(16'h1B9C4,4);
TASK_PP(16'h1B9C5,4);
TASK_PP(16'h1B9C6,4);
TASK_PP(16'h1B9C7,4);
TASK_PP(16'h1B9C8,4);
TASK_PP(16'h1B9C9,4);
TASK_PP(16'h1B9CA,4);
TASK_PP(16'h1B9CB,4);
TASK_PP(16'h1B9CC,4);
TASK_PP(16'h1B9CD,4);
TASK_PP(16'h1B9CE,4);
TASK_PP(16'h1B9CF,4);
TASK_PP(16'h1B9D0,4);
TASK_PP(16'h1B9D1,4);
TASK_PP(16'h1B9D2,4);
TASK_PP(16'h1B9D3,4);
TASK_PP(16'h1B9D4,4);
TASK_PP(16'h1B9D5,4);
TASK_PP(16'h1B9D6,4);
TASK_PP(16'h1B9D7,4);
TASK_PP(16'h1B9D8,4);
TASK_PP(16'h1B9D9,4);
TASK_PP(16'h1B9DA,4);
TASK_PP(16'h1B9DB,4);
TASK_PP(16'h1B9DC,4);
TASK_PP(16'h1B9DD,4);
TASK_PP(16'h1B9DE,4);
TASK_PP(16'h1B9DF,4);
TASK_PP(16'h1B9E0,4);
TASK_PP(16'h1B9E1,4);
TASK_PP(16'h1B9E2,4);
TASK_PP(16'h1B9E3,4);
TASK_PP(16'h1B9E4,4);
TASK_PP(16'h1B9E5,4);
TASK_PP(16'h1B9E6,4);
TASK_PP(16'h1B9E7,4);
TASK_PP(16'h1B9E8,4);
TASK_PP(16'h1B9E9,4);
TASK_PP(16'h1B9EA,4);
TASK_PP(16'h1B9EB,4);
TASK_PP(16'h1B9EC,4);
TASK_PP(16'h1B9ED,4);
TASK_PP(16'h1B9EE,4);
TASK_PP(16'h1B9EF,4);
TASK_PP(16'h1B9F0,4);
TASK_PP(16'h1B9F1,4);
TASK_PP(16'h1B9F2,4);
TASK_PP(16'h1B9F3,4);
TASK_PP(16'h1B9F4,4);
TASK_PP(16'h1B9F5,4);
TASK_PP(16'h1B9F6,4);
TASK_PP(16'h1B9F7,4);
TASK_PP(16'h1B9F8,4);
TASK_PP(16'h1B9F9,4);
TASK_PP(16'h1B9FA,4);
TASK_PP(16'h1B9FB,4);
TASK_PP(16'h1B9FC,4);
TASK_PP(16'h1B9FD,4);
TASK_PP(16'h1B9FE,4);
TASK_PP(16'h1B9FF,4);
TASK_PP(16'h1BA00,4);
TASK_PP(16'h1BA01,4);
TASK_PP(16'h1BA02,4);
TASK_PP(16'h1BA03,4);
TASK_PP(16'h1BA04,4);
TASK_PP(16'h1BA05,4);
TASK_PP(16'h1BA06,4);
TASK_PP(16'h1BA07,4);
TASK_PP(16'h1BA08,4);
TASK_PP(16'h1BA09,4);
TASK_PP(16'h1BA0A,4);
TASK_PP(16'h1BA0B,4);
TASK_PP(16'h1BA0C,4);
TASK_PP(16'h1BA0D,4);
TASK_PP(16'h1BA0E,4);
TASK_PP(16'h1BA0F,4);
TASK_PP(16'h1BA10,4);
TASK_PP(16'h1BA11,4);
TASK_PP(16'h1BA12,4);
TASK_PP(16'h1BA13,4);
TASK_PP(16'h1BA14,4);
TASK_PP(16'h1BA15,4);
TASK_PP(16'h1BA16,4);
TASK_PP(16'h1BA17,4);
TASK_PP(16'h1BA18,4);
TASK_PP(16'h1BA19,4);
TASK_PP(16'h1BA1A,4);
TASK_PP(16'h1BA1B,4);
TASK_PP(16'h1BA1C,4);
TASK_PP(16'h1BA1D,4);
TASK_PP(16'h1BA1E,4);
TASK_PP(16'h1BA1F,4);
TASK_PP(16'h1BA20,4);
TASK_PP(16'h1BA21,4);
TASK_PP(16'h1BA22,4);
TASK_PP(16'h1BA23,4);
TASK_PP(16'h1BA24,4);
TASK_PP(16'h1BA25,4);
TASK_PP(16'h1BA26,4);
TASK_PP(16'h1BA27,4);
TASK_PP(16'h1BA28,4);
TASK_PP(16'h1BA29,4);
TASK_PP(16'h1BA2A,4);
TASK_PP(16'h1BA2B,4);
TASK_PP(16'h1BA2C,4);
TASK_PP(16'h1BA2D,4);
TASK_PP(16'h1BA2E,4);
TASK_PP(16'h1BA2F,4);
TASK_PP(16'h1BA30,4);
TASK_PP(16'h1BA31,4);
TASK_PP(16'h1BA32,4);
TASK_PP(16'h1BA33,4);
TASK_PP(16'h1BA34,4);
TASK_PP(16'h1BA35,4);
TASK_PP(16'h1BA36,4);
TASK_PP(16'h1BA37,4);
TASK_PP(16'h1BA38,4);
TASK_PP(16'h1BA39,4);
TASK_PP(16'h1BA3A,4);
TASK_PP(16'h1BA3B,4);
TASK_PP(16'h1BA3C,4);
TASK_PP(16'h1BA3D,4);
TASK_PP(16'h1BA3E,4);
TASK_PP(16'h1BA3F,4);
TASK_PP(16'h1BA40,4);
TASK_PP(16'h1BA41,4);
TASK_PP(16'h1BA42,4);
TASK_PP(16'h1BA43,4);
TASK_PP(16'h1BA44,4);
TASK_PP(16'h1BA45,4);
TASK_PP(16'h1BA46,4);
TASK_PP(16'h1BA47,4);
TASK_PP(16'h1BA48,4);
TASK_PP(16'h1BA49,4);
TASK_PP(16'h1BA4A,4);
TASK_PP(16'h1BA4B,4);
TASK_PP(16'h1BA4C,4);
TASK_PP(16'h1BA4D,4);
TASK_PP(16'h1BA4E,4);
TASK_PP(16'h1BA4F,4);
TASK_PP(16'h1BA50,4);
TASK_PP(16'h1BA51,4);
TASK_PP(16'h1BA52,4);
TASK_PP(16'h1BA53,4);
TASK_PP(16'h1BA54,4);
TASK_PP(16'h1BA55,4);
TASK_PP(16'h1BA56,4);
TASK_PP(16'h1BA57,4);
TASK_PP(16'h1BA58,4);
TASK_PP(16'h1BA59,4);
TASK_PP(16'h1BA5A,4);
TASK_PP(16'h1BA5B,4);
TASK_PP(16'h1BA5C,4);
TASK_PP(16'h1BA5D,4);
TASK_PP(16'h1BA5E,4);
TASK_PP(16'h1BA5F,4);
TASK_PP(16'h1BA60,4);
TASK_PP(16'h1BA61,4);
TASK_PP(16'h1BA62,4);
TASK_PP(16'h1BA63,4);
TASK_PP(16'h1BA64,4);
TASK_PP(16'h1BA65,4);
TASK_PP(16'h1BA66,4);
TASK_PP(16'h1BA67,4);
TASK_PP(16'h1BA68,4);
TASK_PP(16'h1BA69,4);
TASK_PP(16'h1BA6A,4);
TASK_PP(16'h1BA6B,4);
TASK_PP(16'h1BA6C,4);
TASK_PP(16'h1BA6D,4);
TASK_PP(16'h1BA6E,4);
TASK_PP(16'h1BA6F,4);
TASK_PP(16'h1BA70,4);
TASK_PP(16'h1BA71,4);
TASK_PP(16'h1BA72,4);
TASK_PP(16'h1BA73,4);
TASK_PP(16'h1BA74,4);
TASK_PP(16'h1BA75,4);
TASK_PP(16'h1BA76,4);
TASK_PP(16'h1BA77,4);
TASK_PP(16'h1BA78,4);
TASK_PP(16'h1BA79,4);
TASK_PP(16'h1BA7A,4);
TASK_PP(16'h1BA7B,4);
TASK_PP(16'h1BA7C,4);
TASK_PP(16'h1BA7D,4);
TASK_PP(16'h1BA7E,4);
TASK_PP(16'h1BA7F,4);
TASK_PP(16'h1BA80,4);
TASK_PP(16'h1BA81,4);
TASK_PP(16'h1BA82,4);
TASK_PP(16'h1BA83,4);
TASK_PP(16'h1BA84,4);
TASK_PP(16'h1BA85,4);
TASK_PP(16'h1BA86,4);
TASK_PP(16'h1BA87,4);
TASK_PP(16'h1BA88,4);
TASK_PP(16'h1BA89,4);
TASK_PP(16'h1BA8A,4);
TASK_PP(16'h1BA8B,4);
TASK_PP(16'h1BA8C,4);
TASK_PP(16'h1BA8D,4);
TASK_PP(16'h1BA8E,4);
TASK_PP(16'h1BA8F,4);
TASK_PP(16'h1BA90,4);
TASK_PP(16'h1BA91,4);
TASK_PP(16'h1BA92,4);
TASK_PP(16'h1BA93,4);
TASK_PP(16'h1BA94,4);
TASK_PP(16'h1BA95,4);
TASK_PP(16'h1BA96,4);
TASK_PP(16'h1BA97,4);
TASK_PP(16'h1BA98,4);
TASK_PP(16'h1BA99,4);
TASK_PP(16'h1BA9A,4);
TASK_PP(16'h1BA9B,4);
TASK_PP(16'h1BA9C,4);
TASK_PP(16'h1BA9D,4);
TASK_PP(16'h1BA9E,4);
TASK_PP(16'h1BA9F,4);
TASK_PP(16'h1BAA0,4);
TASK_PP(16'h1BAA1,4);
TASK_PP(16'h1BAA2,4);
TASK_PP(16'h1BAA3,4);
TASK_PP(16'h1BAA4,4);
TASK_PP(16'h1BAA5,4);
TASK_PP(16'h1BAA6,4);
TASK_PP(16'h1BAA7,4);
TASK_PP(16'h1BAA8,4);
TASK_PP(16'h1BAA9,4);
TASK_PP(16'h1BAAA,4);
TASK_PP(16'h1BAAB,4);
TASK_PP(16'h1BAAC,4);
TASK_PP(16'h1BAAD,4);
TASK_PP(16'h1BAAE,4);
TASK_PP(16'h1BAAF,4);
TASK_PP(16'h1BAB0,4);
TASK_PP(16'h1BAB1,4);
TASK_PP(16'h1BAB2,4);
TASK_PP(16'h1BAB3,4);
TASK_PP(16'h1BAB4,4);
TASK_PP(16'h1BAB5,4);
TASK_PP(16'h1BAB6,4);
TASK_PP(16'h1BAB7,4);
TASK_PP(16'h1BAB8,4);
TASK_PP(16'h1BAB9,4);
TASK_PP(16'h1BABA,4);
TASK_PP(16'h1BABB,4);
TASK_PP(16'h1BABC,4);
TASK_PP(16'h1BABD,4);
TASK_PP(16'h1BABE,4);
TASK_PP(16'h1BABF,4);
TASK_PP(16'h1BAC0,4);
TASK_PP(16'h1BAC1,4);
TASK_PP(16'h1BAC2,4);
TASK_PP(16'h1BAC3,4);
TASK_PP(16'h1BAC4,4);
TASK_PP(16'h1BAC5,4);
TASK_PP(16'h1BAC6,4);
TASK_PP(16'h1BAC7,4);
TASK_PP(16'h1BAC8,4);
TASK_PP(16'h1BAC9,4);
TASK_PP(16'h1BACA,4);
TASK_PP(16'h1BACB,4);
TASK_PP(16'h1BACC,4);
TASK_PP(16'h1BACD,4);
TASK_PP(16'h1BACE,4);
TASK_PP(16'h1BACF,4);
TASK_PP(16'h1BAD0,4);
TASK_PP(16'h1BAD1,4);
TASK_PP(16'h1BAD2,4);
TASK_PP(16'h1BAD3,4);
TASK_PP(16'h1BAD4,4);
TASK_PP(16'h1BAD5,4);
TASK_PP(16'h1BAD6,4);
TASK_PP(16'h1BAD7,4);
TASK_PP(16'h1BAD8,4);
TASK_PP(16'h1BAD9,4);
TASK_PP(16'h1BADA,4);
TASK_PP(16'h1BADB,4);
TASK_PP(16'h1BADC,4);
TASK_PP(16'h1BADD,4);
TASK_PP(16'h1BADE,4);
TASK_PP(16'h1BADF,4);
TASK_PP(16'h1BAE0,4);
TASK_PP(16'h1BAE1,4);
TASK_PP(16'h1BAE2,4);
TASK_PP(16'h1BAE3,4);
TASK_PP(16'h1BAE4,4);
TASK_PP(16'h1BAE5,4);
TASK_PP(16'h1BAE6,4);
TASK_PP(16'h1BAE7,4);
TASK_PP(16'h1BAE8,4);
TASK_PP(16'h1BAE9,4);
TASK_PP(16'h1BAEA,4);
TASK_PP(16'h1BAEB,4);
TASK_PP(16'h1BAEC,4);
TASK_PP(16'h1BAED,4);
TASK_PP(16'h1BAEE,4);
TASK_PP(16'h1BAEF,4);
TASK_PP(16'h1BAF0,4);
TASK_PP(16'h1BAF1,4);
TASK_PP(16'h1BAF2,4);
TASK_PP(16'h1BAF3,4);
TASK_PP(16'h1BAF4,4);
TASK_PP(16'h1BAF5,4);
TASK_PP(16'h1BAF6,4);
TASK_PP(16'h1BAF7,4);
TASK_PP(16'h1BAF8,4);
TASK_PP(16'h1BAF9,4);
TASK_PP(16'h1BAFA,4);
TASK_PP(16'h1BAFB,4);
TASK_PP(16'h1BAFC,4);
TASK_PP(16'h1BAFD,4);
TASK_PP(16'h1BAFE,4);
TASK_PP(16'h1BAFF,4);
TASK_PP(16'h1BB00,4);
TASK_PP(16'h1BB01,4);
TASK_PP(16'h1BB02,4);
TASK_PP(16'h1BB03,4);
TASK_PP(16'h1BB04,4);
TASK_PP(16'h1BB05,4);
TASK_PP(16'h1BB06,4);
TASK_PP(16'h1BB07,4);
TASK_PP(16'h1BB08,4);
TASK_PP(16'h1BB09,4);
TASK_PP(16'h1BB0A,4);
TASK_PP(16'h1BB0B,4);
TASK_PP(16'h1BB0C,4);
TASK_PP(16'h1BB0D,4);
TASK_PP(16'h1BB0E,4);
TASK_PP(16'h1BB0F,4);
TASK_PP(16'h1BB10,4);
TASK_PP(16'h1BB11,4);
TASK_PP(16'h1BB12,4);
TASK_PP(16'h1BB13,4);
TASK_PP(16'h1BB14,4);
TASK_PP(16'h1BB15,4);
TASK_PP(16'h1BB16,4);
TASK_PP(16'h1BB17,4);
TASK_PP(16'h1BB18,4);
TASK_PP(16'h1BB19,4);
TASK_PP(16'h1BB1A,4);
TASK_PP(16'h1BB1B,4);
TASK_PP(16'h1BB1C,4);
TASK_PP(16'h1BB1D,4);
TASK_PP(16'h1BB1E,4);
TASK_PP(16'h1BB1F,4);
TASK_PP(16'h1BB20,4);
TASK_PP(16'h1BB21,4);
TASK_PP(16'h1BB22,4);
TASK_PP(16'h1BB23,4);
TASK_PP(16'h1BB24,4);
TASK_PP(16'h1BB25,4);
TASK_PP(16'h1BB26,4);
TASK_PP(16'h1BB27,4);
TASK_PP(16'h1BB28,4);
TASK_PP(16'h1BB29,4);
TASK_PP(16'h1BB2A,4);
TASK_PP(16'h1BB2B,4);
TASK_PP(16'h1BB2C,4);
TASK_PP(16'h1BB2D,4);
TASK_PP(16'h1BB2E,4);
TASK_PP(16'h1BB2F,4);
TASK_PP(16'h1BB30,4);
TASK_PP(16'h1BB31,4);
TASK_PP(16'h1BB32,4);
TASK_PP(16'h1BB33,4);
TASK_PP(16'h1BB34,4);
TASK_PP(16'h1BB35,4);
TASK_PP(16'h1BB36,4);
TASK_PP(16'h1BB37,4);
TASK_PP(16'h1BB38,4);
TASK_PP(16'h1BB39,4);
TASK_PP(16'h1BB3A,4);
TASK_PP(16'h1BB3B,4);
TASK_PP(16'h1BB3C,4);
TASK_PP(16'h1BB3D,4);
TASK_PP(16'h1BB3E,4);
TASK_PP(16'h1BB3F,4);
TASK_PP(16'h1BB40,4);
TASK_PP(16'h1BB41,4);
TASK_PP(16'h1BB42,4);
TASK_PP(16'h1BB43,4);
TASK_PP(16'h1BB44,4);
TASK_PP(16'h1BB45,4);
TASK_PP(16'h1BB46,4);
TASK_PP(16'h1BB47,4);
TASK_PP(16'h1BB48,4);
TASK_PP(16'h1BB49,4);
TASK_PP(16'h1BB4A,4);
TASK_PP(16'h1BB4B,4);
TASK_PP(16'h1BB4C,4);
TASK_PP(16'h1BB4D,4);
TASK_PP(16'h1BB4E,4);
TASK_PP(16'h1BB4F,4);
TASK_PP(16'h1BB50,4);
TASK_PP(16'h1BB51,4);
TASK_PP(16'h1BB52,4);
TASK_PP(16'h1BB53,4);
TASK_PP(16'h1BB54,4);
TASK_PP(16'h1BB55,4);
TASK_PP(16'h1BB56,4);
TASK_PP(16'h1BB57,4);
TASK_PP(16'h1BB58,4);
TASK_PP(16'h1BB59,4);
TASK_PP(16'h1BB5A,4);
TASK_PP(16'h1BB5B,4);
TASK_PP(16'h1BB5C,4);
TASK_PP(16'h1BB5D,4);
TASK_PP(16'h1BB5E,4);
TASK_PP(16'h1BB5F,4);
TASK_PP(16'h1BB60,4);
TASK_PP(16'h1BB61,4);
TASK_PP(16'h1BB62,4);
TASK_PP(16'h1BB63,4);
TASK_PP(16'h1BB64,4);
TASK_PP(16'h1BB65,4);
TASK_PP(16'h1BB66,4);
TASK_PP(16'h1BB67,4);
TASK_PP(16'h1BB68,4);
TASK_PP(16'h1BB69,4);
TASK_PP(16'h1BB6A,4);
TASK_PP(16'h1BB6B,4);
TASK_PP(16'h1BB6C,4);
TASK_PP(16'h1BB6D,4);
TASK_PP(16'h1BB6E,4);
TASK_PP(16'h1BB6F,4);
TASK_PP(16'h1BB70,4);
TASK_PP(16'h1BB71,4);
TASK_PP(16'h1BB72,4);
TASK_PP(16'h1BB73,4);
TASK_PP(16'h1BB74,4);
TASK_PP(16'h1BB75,4);
TASK_PP(16'h1BB76,4);
TASK_PP(16'h1BB77,4);
TASK_PP(16'h1BB78,4);
TASK_PP(16'h1BB79,4);
TASK_PP(16'h1BB7A,4);
TASK_PP(16'h1BB7B,4);
TASK_PP(16'h1BB7C,4);
TASK_PP(16'h1BB7D,4);
TASK_PP(16'h1BB7E,4);
TASK_PP(16'h1BB7F,4);
TASK_PP(16'h1BB80,4);
TASK_PP(16'h1BB81,4);
TASK_PP(16'h1BB82,4);
TASK_PP(16'h1BB83,4);
TASK_PP(16'h1BB84,4);
TASK_PP(16'h1BB85,4);
TASK_PP(16'h1BB86,4);
TASK_PP(16'h1BB87,4);
TASK_PP(16'h1BB88,4);
TASK_PP(16'h1BB89,4);
TASK_PP(16'h1BB8A,4);
TASK_PP(16'h1BB8B,4);
TASK_PP(16'h1BB8C,4);
TASK_PP(16'h1BB8D,4);
TASK_PP(16'h1BB8E,4);
TASK_PP(16'h1BB8F,4);
TASK_PP(16'h1BB90,4);
TASK_PP(16'h1BB91,4);
TASK_PP(16'h1BB92,4);
TASK_PP(16'h1BB93,4);
TASK_PP(16'h1BB94,4);
TASK_PP(16'h1BB95,4);
TASK_PP(16'h1BB96,4);
TASK_PP(16'h1BB97,4);
TASK_PP(16'h1BB98,4);
TASK_PP(16'h1BB99,4);
TASK_PP(16'h1BB9A,4);
TASK_PP(16'h1BB9B,4);
TASK_PP(16'h1BB9C,4);
TASK_PP(16'h1BB9D,4);
TASK_PP(16'h1BB9E,4);
TASK_PP(16'h1BB9F,4);
TASK_PP(16'h1BBA0,4);
TASK_PP(16'h1BBA1,4);
TASK_PP(16'h1BBA2,4);
TASK_PP(16'h1BBA3,4);
TASK_PP(16'h1BBA4,4);
TASK_PP(16'h1BBA5,4);
TASK_PP(16'h1BBA6,4);
TASK_PP(16'h1BBA7,4);
TASK_PP(16'h1BBA8,4);
TASK_PP(16'h1BBA9,4);
TASK_PP(16'h1BBAA,4);
TASK_PP(16'h1BBAB,4);
TASK_PP(16'h1BBAC,4);
TASK_PP(16'h1BBAD,4);
TASK_PP(16'h1BBAE,4);
TASK_PP(16'h1BBAF,4);
TASK_PP(16'h1BBB0,4);
TASK_PP(16'h1BBB1,4);
TASK_PP(16'h1BBB2,4);
TASK_PP(16'h1BBB3,4);
TASK_PP(16'h1BBB4,4);
TASK_PP(16'h1BBB5,4);
TASK_PP(16'h1BBB6,4);
TASK_PP(16'h1BBB7,4);
TASK_PP(16'h1BBB8,4);
TASK_PP(16'h1BBB9,4);
TASK_PP(16'h1BBBA,4);
TASK_PP(16'h1BBBB,4);
TASK_PP(16'h1BBBC,4);
TASK_PP(16'h1BBBD,4);
TASK_PP(16'h1BBBE,4);
TASK_PP(16'h1BBBF,4);
TASK_PP(16'h1BBC0,4);
TASK_PP(16'h1BBC1,4);
TASK_PP(16'h1BBC2,4);
TASK_PP(16'h1BBC3,4);
TASK_PP(16'h1BBC4,4);
TASK_PP(16'h1BBC5,4);
TASK_PP(16'h1BBC6,4);
TASK_PP(16'h1BBC7,4);
TASK_PP(16'h1BBC8,4);
TASK_PP(16'h1BBC9,4);
TASK_PP(16'h1BBCA,4);
TASK_PP(16'h1BBCB,4);
TASK_PP(16'h1BBCC,4);
TASK_PP(16'h1BBCD,4);
TASK_PP(16'h1BBCE,4);
TASK_PP(16'h1BBCF,4);
TASK_PP(16'h1BBD0,4);
TASK_PP(16'h1BBD1,4);
TASK_PP(16'h1BBD2,4);
TASK_PP(16'h1BBD3,4);
TASK_PP(16'h1BBD4,4);
TASK_PP(16'h1BBD5,4);
TASK_PP(16'h1BBD6,4);
TASK_PP(16'h1BBD7,4);
TASK_PP(16'h1BBD8,4);
TASK_PP(16'h1BBD9,4);
TASK_PP(16'h1BBDA,4);
TASK_PP(16'h1BBDB,4);
TASK_PP(16'h1BBDC,4);
TASK_PP(16'h1BBDD,4);
TASK_PP(16'h1BBDE,4);
TASK_PP(16'h1BBDF,4);
TASK_PP(16'h1BBE0,4);
TASK_PP(16'h1BBE1,4);
TASK_PP(16'h1BBE2,4);
TASK_PP(16'h1BBE3,4);
TASK_PP(16'h1BBE4,4);
TASK_PP(16'h1BBE5,4);
TASK_PP(16'h1BBE6,4);
TASK_PP(16'h1BBE7,4);
TASK_PP(16'h1BBE8,4);
TASK_PP(16'h1BBE9,4);
TASK_PP(16'h1BBEA,4);
TASK_PP(16'h1BBEB,4);
TASK_PP(16'h1BBEC,4);
TASK_PP(16'h1BBED,4);
TASK_PP(16'h1BBEE,4);
TASK_PP(16'h1BBEF,4);
TASK_PP(16'h1BBF0,4);
TASK_PP(16'h1BBF1,4);
TASK_PP(16'h1BBF2,4);
TASK_PP(16'h1BBF3,4);
TASK_PP(16'h1BBF4,4);
TASK_PP(16'h1BBF5,4);
TASK_PP(16'h1BBF6,4);
TASK_PP(16'h1BBF7,4);
TASK_PP(16'h1BBF8,4);
TASK_PP(16'h1BBF9,4);
TASK_PP(16'h1BBFA,4);
TASK_PP(16'h1BBFB,4);
TASK_PP(16'h1BBFC,4);
TASK_PP(16'h1BBFD,4);
TASK_PP(16'h1BBFE,4);
TASK_PP(16'h1BBFF,4);
TASK_PP(16'h1BC00,4);
TASK_PP(16'h1BC01,4);
TASK_PP(16'h1BC02,4);
TASK_PP(16'h1BC03,4);
TASK_PP(16'h1BC04,4);
TASK_PP(16'h1BC05,4);
TASK_PP(16'h1BC06,4);
TASK_PP(16'h1BC07,4);
TASK_PP(16'h1BC08,4);
TASK_PP(16'h1BC09,4);
TASK_PP(16'h1BC0A,4);
TASK_PP(16'h1BC0B,4);
TASK_PP(16'h1BC0C,4);
TASK_PP(16'h1BC0D,4);
TASK_PP(16'h1BC0E,4);
TASK_PP(16'h1BC0F,4);
TASK_PP(16'h1BC10,4);
TASK_PP(16'h1BC11,4);
TASK_PP(16'h1BC12,4);
TASK_PP(16'h1BC13,4);
TASK_PP(16'h1BC14,4);
TASK_PP(16'h1BC15,4);
TASK_PP(16'h1BC16,4);
TASK_PP(16'h1BC17,4);
TASK_PP(16'h1BC18,4);
TASK_PP(16'h1BC19,4);
TASK_PP(16'h1BC1A,4);
TASK_PP(16'h1BC1B,4);
TASK_PP(16'h1BC1C,4);
TASK_PP(16'h1BC1D,4);
TASK_PP(16'h1BC1E,4);
TASK_PP(16'h1BC1F,4);
TASK_PP(16'h1BC20,4);
TASK_PP(16'h1BC21,4);
TASK_PP(16'h1BC22,4);
TASK_PP(16'h1BC23,4);
TASK_PP(16'h1BC24,4);
TASK_PP(16'h1BC25,4);
TASK_PP(16'h1BC26,4);
TASK_PP(16'h1BC27,4);
TASK_PP(16'h1BC28,4);
TASK_PP(16'h1BC29,4);
TASK_PP(16'h1BC2A,4);
TASK_PP(16'h1BC2B,4);
TASK_PP(16'h1BC2C,4);
TASK_PP(16'h1BC2D,4);
TASK_PP(16'h1BC2E,4);
TASK_PP(16'h1BC2F,4);
TASK_PP(16'h1BC30,4);
TASK_PP(16'h1BC31,4);
TASK_PP(16'h1BC32,4);
TASK_PP(16'h1BC33,4);
TASK_PP(16'h1BC34,4);
TASK_PP(16'h1BC35,4);
TASK_PP(16'h1BC36,4);
TASK_PP(16'h1BC37,4);
TASK_PP(16'h1BC38,4);
TASK_PP(16'h1BC39,4);
TASK_PP(16'h1BC3A,4);
TASK_PP(16'h1BC3B,4);
TASK_PP(16'h1BC3C,4);
TASK_PP(16'h1BC3D,4);
TASK_PP(16'h1BC3E,4);
TASK_PP(16'h1BC3F,4);
TASK_PP(16'h1BC40,4);
TASK_PP(16'h1BC41,4);
TASK_PP(16'h1BC42,4);
TASK_PP(16'h1BC43,4);
TASK_PP(16'h1BC44,4);
TASK_PP(16'h1BC45,4);
TASK_PP(16'h1BC46,4);
TASK_PP(16'h1BC47,4);
TASK_PP(16'h1BC48,4);
TASK_PP(16'h1BC49,4);
TASK_PP(16'h1BC4A,4);
TASK_PP(16'h1BC4B,4);
TASK_PP(16'h1BC4C,4);
TASK_PP(16'h1BC4D,4);
TASK_PP(16'h1BC4E,4);
TASK_PP(16'h1BC4F,4);
TASK_PP(16'h1BC50,4);
TASK_PP(16'h1BC51,4);
TASK_PP(16'h1BC52,4);
TASK_PP(16'h1BC53,4);
TASK_PP(16'h1BC54,4);
TASK_PP(16'h1BC55,4);
TASK_PP(16'h1BC56,4);
TASK_PP(16'h1BC57,4);
TASK_PP(16'h1BC58,4);
TASK_PP(16'h1BC59,4);
TASK_PP(16'h1BC5A,4);
TASK_PP(16'h1BC5B,4);
TASK_PP(16'h1BC5C,4);
TASK_PP(16'h1BC5D,4);
TASK_PP(16'h1BC5E,4);
TASK_PP(16'h1BC5F,4);
TASK_PP(16'h1BC60,4);
TASK_PP(16'h1BC61,4);
TASK_PP(16'h1BC62,4);
TASK_PP(16'h1BC63,4);
TASK_PP(16'h1BC64,4);
TASK_PP(16'h1BC65,4);
TASK_PP(16'h1BC66,4);
TASK_PP(16'h1BC67,4);
TASK_PP(16'h1BC68,4);
TASK_PP(16'h1BC69,4);
TASK_PP(16'h1BC6A,4);
TASK_PP(16'h1BC6B,4);
TASK_PP(16'h1BC6C,4);
TASK_PP(16'h1BC6D,4);
TASK_PP(16'h1BC6E,4);
TASK_PP(16'h1BC6F,4);
TASK_PP(16'h1BC70,4);
TASK_PP(16'h1BC71,4);
TASK_PP(16'h1BC72,4);
TASK_PP(16'h1BC73,4);
TASK_PP(16'h1BC74,4);
TASK_PP(16'h1BC75,4);
TASK_PP(16'h1BC76,4);
TASK_PP(16'h1BC77,4);
TASK_PP(16'h1BC78,4);
TASK_PP(16'h1BC79,4);
TASK_PP(16'h1BC7A,4);
TASK_PP(16'h1BC7B,4);
TASK_PP(16'h1BC7C,4);
TASK_PP(16'h1BC7D,4);
TASK_PP(16'h1BC7E,4);
TASK_PP(16'h1BC7F,4);
TASK_PP(16'h1BC80,4);
TASK_PP(16'h1BC81,4);
TASK_PP(16'h1BC82,4);
TASK_PP(16'h1BC83,4);
TASK_PP(16'h1BC84,4);
TASK_PP(16'h1BC85,4);
TASK_PP(16'h1BC86,4);
TASK_PP(16'h1BC87,4);
TASK_PP(16'h1BC88,4);
TASK_PP(16'h1BC89,4);
TASK_PP(16'h1BC8A,4);
TASK_PP(16'h1BC8B,4);
TASK_PP(16'h1BC8C,4);
TASK_PP(16'h1BC8D,4);
TASK_PP(16'h1BC8E,4);
TASK_PP(16'h1BC8F,4);
TASK_PP(16'h1BC90,4);
TASK_PP(16'h1BC91,4);
TASK_PP(16'h1BC92,4);
TASK_PP(16'h1BC93,4);
TASK_PP(16'h1BC94,4);
TASK_PP(16'h1BC95,4);
TASK_PP(16'h1BC96,4);
TASK_PP(16'h1BC97,4);
TASK_PP(16'h1BC98,4);
TASK_PP(16'h1BC99,4);
TASK_PP(16'h1BC9A,4);
TASK_PP(16'h1BC9B,4);
TASK_PP(16'h1BC9C,4);
TASK_PP(16'h1BC9D,4);
TASK_PP(16'h1BC9E,4);
TASK_PP(16'h1BC9F,4);
TASK_PP(16'h1BCA0,4);
TASK_PP(16'h1BCA1,4);
TASK_PP(16'h1BCA2,4);
TASK_PP(16'h1BCA3,4);
TASK_PP(16'h1BCA4,4);
TASK_PP(16'h1BCA5,4);
TASK_PP(16'h1BCA6,4);
TASK_PP(16'h1BCA7,4);
TASK_PP(16'h1BCA8,4);
TASK_PP(16'h1BCA9,4);
TASK_PP(16'h1BCAA,4);
TASK_PP(16'h1BCAB,4);
TASK_PP(16'h1BCAC,4);
TASK_PP(16'h1BCAD,4);
TASK_PP(16'h1BCAE,4);
TASK_PP(16'h1BCAF,4);
TASK_PP(16'h1BCB0,4);
TASK_PP(16'h1BCB1,4);
TASK_PP(16'h1BCB2,4);
TASK_PP(16'h1BCB3,4);
TASK_PP(16'h1BCB4,4);
TASK_PP(16'h1BCB5,4);
TASK_PP(16'h1BCB6,4);
TASK_PP(16'h1BCB7,4);
TASK_PP(16'h1BCB8,4);
TASK_PP(16'h1BCB9,4);
TASK_PP(16'h1BCBA,4);
TASK_PP(16'h1BCBB,4);
TASK_PP(16'h1BCBC,4);
TASK_PP(16'h1BCBD,4);
TASK_PP(16'h1BCBE,4);
TASK_PP(16'h1BCBF,4);
TASK_PP(16'h1BCC0,4);
TASK_PP(16'h1BCC1,4);
TASK_PP(16'h1BCC2,4);
TASK_PP(16'h1BCC3,4);
TASK_PP(16'h1BCC4,4);
TASK_PP(16'h1BCC5,4);
TASK_PP(16'h1BCC6,4);
TASK_PP(16'h1BCC7,4);
TASK_PP(16'h1BCC8,4);
TASK_PP(16'h1BCC9,4);
TASK_PP(16'h1BCCA,4);
TASK_PP(16'h1BCCB,4);
TASK_PP(16'h1BCCC,4);
TASK_PP(16'h1BCCD,4);
TASK_PP(16'h1BCCE,4);
TASK_PP(16'h1BCCF,4);
TASK_PP(16'h1BCD0,4);
TASK_PP(16'h1BCD1,4);
TASK_PP(16'h1BCD2,4);
TASK_PP(16'h1BCD3,4);
TASK_PP(16'h1BCD4,4);
TASK_PP(16'h1BCD5,4);
TASK_PP(16'h1BCD6,4);
TASK_PP(16'h1BCD7,4);
TASK_PP(16'h1BCD8,4);
TASK_PP(16'h1BCD9,4);
TASK_PP(16'h1BCDA,4);
TASK_PP(16'h1BCDB,4);
TASK_PP(16'h1BCDC,4);
TASK_PP(16'h1BCDD,4);
TASK_PP(16'h1BCDE,4);
TASK_PP(16'h1BCDF,4);
TASK_PP(16'h1BCE0,4);
TASK_PP(16'h1BCE1,4);
TASK_PP(16'h1BCE2,4);
TASK_PP(16'h1BCE3,4);
TASK_PP(16'h1BCE4,4);
TASK_PP(16'h1BCE5,4);
TASK_PP(16'h1BCE6,4);
TASK_PP(16'h1BCE7,4);
TASK_PP(16'h1BCE8,4);
TASK_PP(16'h1BCE9,4);
TASK_PP(16'h1BCEA,4);
TASK_PP(16'h1BCEB,4);
TASK_PP(16'h1BCEC,4);
TASK_PP(16'h1BCED,4);
TASK_PP(16'h1BCEE,4);
TASK_PP(16'h1BCEF,4);
TASK_PP(16'h1BCF0,4);
TASK_PP(16'h1BCF1,4);
TASK_PP(16'h1BCF2,4);
TASK_PP(16'h1BCF3,4);
TASK_PP(16'h1BCF4,4);
TASK_PP(16'h1BCF5,4);
TASK_PP(16'h1BCF6,4);
TASK_PP(16'h1BCF7,4);
TASK_PP(16'h1BCF8,4);
TASK_PP(16'h1BCF9,4);
TASK_PP(16'h1BCFA,4);
TASK_PP(16'h1BCFB,4);
TASK_PP(16'h1BCFC,4);
TASK_PP(16'h1BCFD,4);
TASK_PP(16'h1BCFE,4);
TASK_PP(16'h1BCFF,4);
TASK_PP(16'h1BD00,4);
TASK_PP(16'h1BD01,4);
TASK_PP(16'h1BD02,4);
TASK_PP(16'h1BD03,4);
TASK_PP(16'h1BD04,4);
TASK_PP(16'h1BD05,4);
TASK_PP(16'h1BD06,4);
TASK_PP(16'h1BD07,4);
TASK_PP(16'h1BD08,4);
TASK_PP(16'h1BD09,4);
TASK_PP(16'h1BD0A,4);
TASK_PP(16'h1BD0B,4);
TASK_PP(16'h1BD0C,4);
TASK_PP(16'h1BD0D,4);
TASK_PP(16'h1BD0E,4);
TASK_PP(16'h1BD0F,4);
TASK_PP(16'h1BD10,4);
TASK_PP(16'h1BD11,4);
TASK_PP(16'h1BD12,4);
TASK_PP(16'h1BD13,4);
TASK_PP(16'h1BD14,4);
TASK_PP(16'h1BD15,4);
TASK_PP(16'h1BD16,4);
TASK_PP(16'h1BD17,4);
TASK_PP(16'h1BD18,4);
TASK_PP(16'h1BD19,4);
TASK_PP(16'h1BD1A,4);
TASK_PP(16'h1BD1B,4);
TASK_PP(16'h1BD1C,4);
TASK_PP(16'h1BD1D,4);
TASK_PP(16'h1BD1E,4);
TASK_PP(16'h1BD1F,4);
TASK_PP(16'h1BD20,4);
TASK_PP(16'h1BD21,4);
TASK_PP(16'h1BD22,4);
TASK_PP(16'h1BD23,4);
TASK_PP(16'h1BD24,4);
TASK_PP(16'h1BD25,4);
TASK_PP(16'h1BD26,4);
TASK_PP(16'h1BD27,4);
TASK_PP(16'h1BD28,4);
TASK_PP(16'h1BD29,4);
TASK_PP(16'h1BD2A,4);
TASK_PP(16'h1BD2B,4);
TASK_PP(16'h1BD2C,4);
TASK_PP(16'h1BD2D,4);
TASK_PP(16'h1BD2E,4);
TASK_PP(16'h1BD2F,4);
TASK_PP(16'h1BD30,4);
TASK_PP(16'h1BD31,4);
TASK_PP(16'h1BD32,4);
TASK_PP(16'h1BD33,4);
TASK_PP(16'h1BD34,4);
TASK_PP(16'h1BD35,4);
TASK_PP(16'h1BD36,4);
TASK_PP(16'h1BD37,4);
TASK_PP(16'h1BD38,4);
TASK_PP(16'h1BD39,4);
TASK_PP(16'h1BD3A,4);
TASK_PP(16'h1BD3B,4);
TASK_PP(16'h1BD3C,4);
TASK_PP(16'h1BD3D,4);
TASK_PP(16'h1BD3E,4);
TASK_PP(16'h1BD3F,4);
TASK_PP(16'h1BD40,4);
TASK_PP(16'h1BD41,4);
TASK_PP(16'h1BD42,4);
TASK_PP(16'h1BD43,4);
TASK_PP(16'h1BD44,4);
TASK_PP(16'h1BD45,4);
TASK_PP(16'h1BD46,4);
TASK_PP(16'h1BD47,4);
TASK_PP(16'h1BD48,4);
TASK_PP(16'h1BD49,4);
TASK_PP(16'h1BD4A,4);
TASK_PP(16'h1BD4B,4);
TASK_PP(16'h1BD4C,4);
TASK_PP(16'h1BD4D,4);
TASK_PP(16'h1BD4E,4);
TASK_PP(16'h1BD4F,4);
TASK_PP(16'h1BD50,4);
TASK_PP(16'h1BD51,4);
TASK_PP(16'h1BD52,4);
TASK_PP(16'h1BD53,4);
TASK_PP(16'h1BD54,4);
TASK_PP(16'h1BD55,4);
TASK_PP(16'h1BD56,4);
TASK_PP(16'h1BD57,4);
TASK_PP(16'h1BD58,4);
TASK_PP(16'h1BD59,4);
TASK_PP(16'h1BD5A,4);
TASK_PP(16'h1BD5B,4);
TASK_PP(16'h1BD5C,4);
TASK_PP(16'h1BD5D,4);
TASK_PP(16'h1BD5E,4);
TASK_PP(16'h1BD5F,4);
TASK_PP(16'h1BD60,4);
TASK_PP(16'h1BD61,4);
TASK_PP(16'h1BD62,4);
TASK_PP(16'h1BD63,4);
TASK_PP(16'h1BD64,4);
TASK_PP(16'h1BD65,4);
TASK_PP(16'h1BD66,4);
TASK_PP(16'h1BD67,4);
TASK_PP(16'h1BD68,4);
TASK_PP(16'h1BD69,4);
TASK_PP(16'h1BD6A,4);
TASK_PP(16'h1BD6B,4);
TASK_PP(16'h1BD6C,4);
TASK_PP(16'h1BD6D,4);
TASK_PP(16'h1BD6E,4);
TASK_PP(16'h1BD6F,4);
TASK_PP(16'h1BD70,4);
TASK_PP(16'h1BD71,4);
TASK_PP(16'h1BD72,4);
TASK_PP(16'h1BD73,4);
TASK_PP(16'h1BD74,4);
TASK_PP(16'h1BD75,4);
TASK_PP(16'h1BD76,4);
TASK_PP(16'h1BD77,4);
TASK_PP(16'h1BD78,4);
TASK_PP(16'h1BD79,4);
TASK_PP(16'h1BD7A,4);
TASK_PP(16'h1BD7B,4);
TASK_PP(16'h1BD7C,4);
TASK_PP(16'h1BD7D,4);
TASK_PP(16'h1BD7E,4);
TASK_PP(16'h1BD7F,4);
TASK_PP(16'h1BD80,4);
TASK_PP(16'h1BD81,4);
TASK_PP(16'h1BD82,4);
TASK_PP(16'h1BD83,4);
TASK_PP(16'h1BD84,4);
TASK_PP(16'h1BD85,4);
TASK_PP(16'h1BD86,4);
TASK_PP(16'h1BD87,4);
TASK_PP(16'h1BD88,4);
TASK_PP(16'h1BD89,4);
TASK_PP(16'h1BD8A,4);
TASK_PP(16'h1BD8B,4);
TASK_PP(16'h1BD8C,4);
TASK_PP(16'h1BD8D,4);
TASK_PP(16'h1BD8E,4);
TASK_PP(16'h1BD8F,4);
TASK_PP(16'h1BD90,4);
TASK_PP(16'h1BD91,4);
TASK_PP(16'h1BD92,4);
TASK_PP(16'h1BD93,4);
TASK_PP(16'h1BD94,4);
TASK_PP(16'h1BD95,4);
TASK_PP(16'h1BD96,4);
TASK_PP(16'h1BD97,4);
TASK_PP(16'h1BD98,4);
TASK_PP(16'h1BD99,4);
TASK_PP(16'h1BD9A,4);
TASK_PP(16'h1BD9B,4);
TASK_PP(16'h1BD9C,4);
TASK_PP(16'h1BD9D,4);
TASK_PP(16'h1BD9E,4);
TASK_PP(16'h1BD9F,4);
TASK_PP(16'h1BDA0,4);
TASK_PP(16'h1BDA1,4);
TASK_PP(16'h1BDA2,4);
TASK_PP(16'h1BDA3,4);
TASK_PP(16'h1BDA4,4);
TASK_PP(16'h1BDA5,4);
TASK_PP(16'h1BDA6,4);
TASK_PP(16'h1BDA7,4);
TASK_PP(16'h1BDA8,4);
TASK_PP(16'h1BDA9,4);
TASK_PP(16'h1BDAA,4);
TASK_PP(16'h1BDAB,4);
TASK_PP(16'h1BDAC,4);
TASK_PP(16'h1BDAD,4);
TASK_PP(16'h1BDAE,4);
TASK_PP(16'h1BDAF,4);
TASK_PP(16'h1BDB0,4);
TASK_PP(16'h1BDB1,4);
TASK_PP(16'h1BDB2,4);
TASK_PP(16'h1BDB3,4);
TASK_PP(16'h1BDB4,4);
TASK_PP(16'h1BDB5,4);
TASK_PP(16'h1BDB6,4);
TASK_PP(16'h1BDB7,4);
TASK_PP(16'h1BDB8,4);
TASK_PP(16'h1BDB9,4);
TASK_PP(16'h1BDBA,4);
TASK_PP(16'h1BDBB,4);
TASK_PP(16'h1BDBC,4);
TASK_PP(16'h1BDBD,4);
TASK_PP(16'h1BDBE,4);
TASK_PP(16'h1BDBF,4);
TASK_PP(16'h1BDC0,4);
TASK_PP(16'h1BDC1,4);
TASK_PP(16'h1BDC2,4);
TASK_PP(16'h1BDC3,4);
TASK_PP(16'h1BDC4,4);
TASK_PP(16'h1BDC5,4);
TASK_PP(16'h1BDC6,4);
TASK_PP(16'h1BDC7,4);
TASK_PP(16'h1BDC8,4);
TASK_PP(16'h1BDC9,4);
TASK_PP(16'h1BDCA,4);
TASK_PP(16'h1BDCB,4);
TASK_PP(16'h1BDCC,4);
TASK_PP(16'h1BDCD,4);
TASK_PP(16'h1BDCE,4);
TASK_PP(16'h1BDCF,4);
TASK_PP(16'h1BDD0,4);
TASK_PP(16'h1BDD1,4);
TASK_PP(16'h1BDD2,4);
TASK_PP(16'h1BDD3,4);
TASK_PP(16'h1BDD4,4);
TASK_PP(16'h1BDD5,4);
TASK_PP(16'h1BDD6,4);
TASK_PP(16'h1BDD7,4);
TASK_PP(16'h1BDD8,4);
TASK_PP(16'h1BDD9,4);
TASK_PP(16'h1BDDA,4);
TASK_PP(16'h1BDDB,4);
TASK_PP(16'h1BDDC,4);
TASK_PP(16'h1BDDD,4);
TASK_PP(16'h1BDDE,4);
TASK_PP(16'h1BDDF,4);
TASK_PP(16'h1BDE0,4);
TASK_PP(16'h1BDE1,4);
TASK_PP(16'h1BDE2,4);
TASK_PP(16'h1BDE3,4);
TASK_PP(16'h1BDE4,4);
TASK_PP(16'h1BDE5,4);
TASK_PP(16'h1BDE6,4);
TASK_PP(16'h1BDE7,4);
TASK_PP(16'h1BDE8,4);
TASK_PP(16'h1BDE9,4);
TASK_PP(16'h1BDEA,4);
TASK_PP(16'h1BDEB,4);
TASK_PP(16'h1BDEC,4);
TASK_PP(16'h1BDED,4);
TASK_PP(16'h1BDEE,4);
TASK_PP(16'h1BDEF,4);
TASK_PP(16'h1BDF0,4);
TASK_PP(16'h1BDF1,4);
TASK_PP(16'h1BDF2,4);
TASK_PP(16'h1BDF3,4);
TASK_PP(16'h1BDF4,4);
TASK_PP(16'h1BDF5,4);
TASK_PP(16'h1BDF6,4);
TASK_PP(16'h1BDF7,4);
TASK_PP(16'h1BDF8,4);
TASK_PP(16'h1BDF9,4);
TASK_PP(16'h1BDFA,4);
TASK_PP(16'h1BDFB,4);
TASK_PP(16'h1BDFC,4);
TASK_PP(16'h1BDFD,4);
TASK_PP(16'h1BDFE,4);
TASK_PP(16'h1BDFF,4);
TASK_PP(16'h1BE00,4);
TASK_PP(16'h1BE01,4);
TASK_PP(16'h1BE02,4);
TASK_PP(16'h1BE03,4);
TASK_PP(16'h1BE04,4);
TASK_PP(16'h1BE05,4);
TASK_PP(16'h1BE06,4);
TASK_PP(16'h1BE07,4);
TASK_PP(16'h1BE08,4);
TASK_PP(16'h1BE09,4);
TASK_PP(16'h1BE0A,4);
TASK_PP(16'h1BE0B,4);
TASK_PP(16'h1BE0C,4);
TASK_PP(16'h1BE0D,4);
TASK_PP(16'h1BE0E,4);
TASK_PP(16'h1BE0F,4);
TASK_PP(16'h1BE10,4);
TASK_PP(16'h1BE11,4);
TASK_PP(16'h1BE12,4);
TASK_PP(16'h1BE13,4);
TASK_PP(16'h1BE14,4);
TASK_PP(16'h1BE15,4);
TASK_PP(16'h1BE16,4);
TASK_PP(16'h1BE17,4);
TASK_PP(16'h1BE18,4);
TASK_PP(16'h1BE19,4);
TASK_PP(16'h1BE1A,4);
TASK_PP(16'h1BE1B,4);
TASK_PP(16'h1BE1C,4);
TASK_PP(16'h1BE1D,4);
TASK_PP(16'h1BE1E,4);
TASK_PP(16'h1BE1F,4);
TASK_PP(16'h1BE20,4);
TASK_PP(16'h1BE21,4);
TASK_PP(16'h1BE22,4);
TASK_PP(16'h1BE23,4);
TASK_PP(16'h1BE24,4);
TASK_PP(16'h1BE25,4);
TASK_PP(16'h1BE26,4);
TASK_PP(16'h1BE27,4);
TASK_PP(16'h1BE28,4);
TASK_PP(16'h1BE29,4);
TASK_PP(16'h1BE2A,4);
TASK_PP(16'h1BE2B,4);
TASK_PP(16'h1BE2C,4);
TASK_PP(16'h1BE2D,4);
TASK_PP(16'h1BE2E,4);
TASK_PP(16'h1BE2F,4);
TASK_PP(16'h1BE30,4);
TASK_PP(16'h1BE31,4);
TASK_PP(16'h1BE32,4);
TASK_PP(16'h1BE33,4);
TASK_PP(16'h1BE34,4);
TASK_PP(16'h1BE35,4);
TASK_PP(16'h1BE36,4);
TASK_PP(16'h1BE37,4);
TASK_PP(16'h1BE38,4);
TASK_PP(16'h1BE39,4);
TASK_PP(16'h1BE3A,4);
TASK_PP(16'h1BE3B,4);
TASK_PP(16'h1BE3C,4);
TASK_PP(16'h1BE3D,4);
TASK_PP(16'h1BE3E,4);
TASK_PP(16'h1BE3F,4);
TASK_PP(16'h1BE40,4);
TASK_PP(16'h1BE41,4);
TASK_PP(16'h1BE42,4);
TASK_PP(16'h1BE43,4);
TASK_PP(16'h1BE44,4);
TASK_PP(16'h1BE45,4);
TASK_PP(16'h1BE46,4);
TASK_PP(16'h1BE47,4);
TASK_PP(16'h1BE48,4);
TASK_PP(16'h1BE49,4);
TASK_PP(16'h1BE4A,4);
TASK_PP(16'h1BE4B,4);
TASK_PP(16'h1BE4C,4);
TASK_PP(16'h1BE4D,4);
TASK_PP(16'h1BE4E,4);
TASK_PP(16'h1BE4F,4);
TASK_PP(16'h1BE50,4);
TASK_PP(16'h1BE51,4);
TASK_PP(16'h1BE52,4);
TASK_PP(16'h1BE53,4);
TASK_PP(16'h1BE54,4);
TASK_PP(16'h1BE55,4);
TASK_PP(16'h1BE56,4);
TASK_PP(16'h1BE57,4);
TASK_PP(16'h1BE58,4);
TASK_PP(16'h1BE59,4);
TASK_PP(16'h1BE5A,4);
TASK_PP(16'h1BE5B,4);
TASK_PP(16'h1BE5C,4);
TASK_PP(16'h1BE5D,4);
TASK_PP(16'h1BE5E,4);
TASK_PP(16'h1BE5F,4);
TASK_PP(16'h1BE60,4);
TASK_PP(16'h1BE61,4);
TASK_PP(16'h1BE62,4);
TASK_PP(16'h1BE63,4);
TASK_PP(16'h1BE64,4);
TASK_PP(16'h1BE65,4);
TASK_PP(16'h1BE66,4);
TASK_PP(16'h1BE67,4);
TASK_PP(16'h1BE68,4);
TASK_PP(16'h1BE69,4);
TASK_PP(16'h1BE6A,4);
TASK_PP(16'h1BE6B,4);
TASK_PP(16'h1BE6C,4);
TASK_PP(16'h1BE6D,4);
TASK_PP(16'h1BE6E,4);
TASK_PP(16'h1BE6F,4);
TASK_PP(16'h1BE70,4);
TASK_PP(16'h1BE71,4);
TASK_PP(16'h1BE72,4);
TASK_PP(16'h1BE73,4);
TASK_PP(16'h1BE74,4);
TASK_PP(16'h1BE75,4);
TASK_PP(16'h1BE76,4);
TASK_PP(16'h1BE77,4);
TASK_PP(16'h1BE78,4);
TASK_PP(16'h1BE79,4);
TASK_PP(16'h1BE7A,4);
TASK_PP(16'h1BE7B,4);
TASK_PP(16'h1BE7C,4);
TASK_PP(16'h1BE7D,4);
TASK_PP(16'h1BE7E,4);
TASK_PP(16'h1BE7F,4);
TASK_PP(16'h1BE80,4);
TASK_PP(16'h1BE81,4);
TASK_PP(16'h1BE82,4);
TASK_PP(16'h1BE83,4);
TASK_PP(16'h1BE84,4);
TASK_PP(16'h1BE85,4);
TASK_PP(16'h1BE86,4);
TASK_PP(16'h1BE87,4);
TASK_PP(16'h1BE88,4);
TASK_PP(16'h1BE89,4);
TASK_PP(16'h1BE8A,4);
TASK_PP(16'h1BE8B,4);
TASK_PP(16'h1BE8C,4);
TASK_PP(16'h1BE8D,4);
TASK_PP(16'h1BE8E,4);
TASK_PP(16'h1BE8F,4);
TASK_PP(16'h1BE90,4);
TASK_PP(16'h1BE91,4);
TASK_PP(16'h1BE92,4);
TASK_PP(16'h1BE93,4);
TASK_PP(16'h1BE94,4);
TASK_PP(16'h1BE95,4);
TASK_PP(16'h1BE96,4);
TASK_PP(16'h1BE97,4);
TASK_PP(16'h1BE98,4);
TASK_PP(16'h1BE99,4);
TASK_PP(16'h1BE9A,4);
TASK_PP(16'h1BE9B,4);
TASK_PP(16'h1BE9C,4);
TASK_PP(16'h1BE9D,4);
TASK_PP(16'h1BE9E,4);
TASK_PP(16'h1BE9F,4);
TASK_PP(16'h1BEA0,4);
TASK_PP(16'h1BEA1,4);
TASK_PP(16'h1BEA2,4);
TASK_PP(16'h1BEA3,4);
TASK_PP(16'h1BEA4,4);
TASK_PP(16'h1BEA5,4);
TASK_PP(16'h1BEA6,4);
TASK_PP(16'h1BEA7,4);
TASK_PP(16'h1BEA8,4);
TASK_PP(16'h1BEA9,4);
TASK_PP(16'h1BEAA,4);
TASK_PP(16'h1BEAB,4);
TASK_PP(16'h1BEAC,4);
TASK_PP(16'h1BEAD,4);
TASK_PP(16'h1BEAE,4);
TASK_PP(16'h1BEAF,4);
TASK_PP(16'h1BEB0,4);
TASK_PP(16'h1BEB1,4);
TASK_PP(16'h1BEB2,4);
TASK_PP(16'h1BEB3,4);
TASK_PP(16'h1BEB4,4);
TASK_PP(16'h1BEB5,4);
TASK_PP(16'h1BEB6,4);
TASK_PP(16'h1BEB7,4);
TASK_PP(16'h1BEB8,4);
TASK_PP(16'h1BEB9,4);
TASK_PP(16'h1BEBA,4);
TASK_PP(16'h1BEBB,4);
TASK_PP(16'h1BEBC,4);
TASK_PP(16'h1BEBD,4);
TASK_PP(16'h1BEBE,4);
TASK_PP(16'h1BEBF,4);
TASK_PP(16'h1BEC0,4);
TASK_PP(16'h1BEC1,4);
TASK_PP(16'h1BEC2,4);
TASK_PP(16'h1BEC3,4);
TASK_PP(16'h1BEC4,4);
TASK_PP(16'h1BEC5,4);
TASK_PP(16'h1BEC6,4);
TASK_PP(16'h1BEC7,4);
TASK_PP(16'h1BEC8,4);
TASK_PP(16'h1BEC9,4);
TASK_PP(16'h1BECA,4);
TASK_PP(16'h1BECB,4);
TASK_PP(16'h1BECC,4);
TASK_PP(16'h1BECD,4);
TASK_PP(16'h1BECE,4);
TASK_PP(16'h1BECF,4);
TASK_PP(16'h1BED0,4);
TASK_PP(16'h1BED1,4);
TASK_PP(16'h1BED2,4);
TASK_PP(16'h1BED3,4);
TASK_PP(16'h1BED4,4);
TASK_PP(16'h1BED5,4);
TASK_PP(16'h1BED6,4);
TASK_PP(16'h1BED7,4);
TASK_PP(16'h1BED8,4);
TASK_PP(16'h1BED9,4);
TASK_PP(16'h1BEDA,4);
TASK_PP(16'h1BEDB,4);
TASK_PP(16'h1BEDC,4);
TASK_PP(16'h1BEDD,4);
TASK_PP(16'h1BEDE,4);
TASK_PP(16'h1BEDF,4);
TASK_PP(16'h1BEE0,4);
TASK_PP(16'h1BEE1,4);
TASK_PP(16'h1BEE2,4);
TASK_PP(16'h1BEE3,4);
TASK_PP(16'h1BEE4,4);
TASK_PP(16'h1BEE5,4);
TASK_PP(16'h1BEE6,4);
TASK_PP(16'h1BEE7,4);
TASK_PP(16'h1BEE8,4);
TASK_PP(16'h1BEE9,4);
TASK_PP(16'h1BEEA,4);
TASK_PP(16'h1BEEB,4);
TASK_PP(16'h1BEEC,4);
TASK_PP(16'h1BEED,4);
TASK_PP(16'h1BEEE,4);
TASK_PP(16'h1BEEF,4);
TASK_PP(16'h1BEF0,4);
TASK_PP(16'h1BEF1,4);
TASK_PP(16'h1BEF2,4);
TASK_PP(16'h1BEF3,4);
TASK_PP(16'h1BEF4,4);
TASK_PP(16'h1BEF5,4);
TASK_PP(16'h1BEF6,4);
TASK_PP(16'h1BEF7,4);
TASK_PP(16'h1BEF8,4);
TASK_PP(16'h1BEF9,4);
TASK_PP(16'h1BEFA,4);
TASK_PP(16'h1BEFB,4);
TASK_PP(16'h1BEFC,4);
TASK_PP(16'h1BEFD,4);
TASK_PP(16'h1BEFE,4);
TASK_PP(16'h1BEFF,4);
TASK_PP(16'h1BF00,4);
TASK_PP(16'h1BF01,4);
TASK_PP(16'h1BF02,4);
TASK_PP(16'h1BF03,4);
TASK_PP(16'h1BF04,4);
TASK_PP(16'h1BF05,4);
TASK_PP(16'h1BF06,4);
TASK_PP(16'h1BF07,4);
TASK_PP(16'h1BF08,4);
TASK_PP(16'h1BF09,4);
TASK_PP(16'h1BF0A,4);
TASK_PP(16'h1BF0B,4);
TASK_PP(16'h1BF0C,4);
TASK_PP(16'h1BF0D,4);
TASK_PP(16'h1BF0E,4);
TASK_PP(16'h1BF0F,4);
TASK_PP(16'h1BF10,4);
TASK_PP(16'h1BF11,4);
TASK_PP(16'h1BF12,4);
TASK_PP(16'h1BF13,4);
TASK_PP(16'h1BF14,4);
TASK_PP(16'h1BF15,4);
TASK_PP(16'h1BF16,4);
TASK_PP(16'h1BF17,4);
TASK_PP(16'h1BF18,4);
TASK_PP(16'h1BF19,4);
TASK_PP(16'h1BF1A,4);
TASK_PP(16'h1BF1B,4);
TASK_PP(16'h1BF1C,4);
TASK_PP(16'h1BF1D,4);
TASK_PP(16'h1BF1E,4);
TASK_PP(16'h1BF1F,4);
TASK_PP(16'h1BF20,4);
TASK_PP(16'h1BF21,4);
TASK_PP(16'h1BF22,4);
TASK_PP(16'h1BF23,4);
TASK_PP(16'h1BF24,4);
TASK_PP(16'h1BF25,4);
TASK_PP(16'h1BF26,4);
TASK_PP(16'h1BF27,4);
TASK_PP(16'h1BF28,4);
TASK_PP(16'h1BF29,4);
TASK_PP(16'h1BF2A,4);
TASK_PP(16'h1BF2B,4);
TASK_PP(16'h1BF2C,4);
TASK_PP(16'h1BF2D,4);
TASK_PP(16'h1BF2E,4);
TASK_PP(16'h1BF2F,4);
TASK_PP(16'h1BF30,4);
TASK_PP(16'h1BF31,4);
TASK_PP(16'h1BF32,4);
TASK_PP(16'h1BF33,4);
TASK_PP(16'h1BF34,4);
TASK_PP(16'h1BF35,4);
TASK_PP(16'h1BF36,4);
TASK_PP(16'h1BF37,4);
TASK_PP(16'h1BF38,4);
TASK_PP(16'h1BF39,4);
TASK_PP(16'h1BF3A,4);
TASK_PP(16'h1BF3B,4);
TASK_PP(16'h1BF3C,4);
TASK_PP(16'h1BF3D,4);
TASK_PP(16'h1BF3E,4);
TASK_PP(16'h1BF3F,4);
TASK_PP(16'h1BF40,4);
TASK_PP(16'h1BF41,4);
TASK_PP(16'h1BF42,4);
TASK_PP(16'h1BF43,4);
TASK_PP(16'h1BF44,4);
TASK_PP(16'h1BF45,4);
TASK_PP(16'h1BF46,4);
TASK_PP(16'h1BF47,4);
TASK_PP(16'h1BF48,4);
TASK_PP(16'h1BF49,4);
TASK_PP(16'h1BF4A,4);
TASK_PP(16'h1BF4B,4);
TASK_PP(16'h1BF4C,4);
TASK_PP(16'h1BF4D,4);
TASK_PP(16'h1BF4E,4);
TASK_PP(16'h1BF4F,4);
TASK_PP(16'h1BF50,4);
TASK_PP(16'h1BF51,4);
TASK_PP(16'h1BF52,4);
TASK_PP(16'h1BF53,4);
TASK_PP(16'h1BF54,4);
TASK_PP(16'h1BF55,4);
TASK_PP(16'h1BF56,4);
TASK_PP(16'h1BF57,4);
TASK_PP(16'h1BF58,4);
TASK_PP(16'h1BF59,4);
TASK_PP(16'h1BF5A,4);
TASK_PP(16'h1BF5B,4);
TASK_PP(16'h1BF5C,4);
TASK_PP(16'h1BF5D,4);
TASK_PP(16'h1BF5E,4);
TASK_PP(16'h1BF5F,4);
TASK_PP(16'h1BF60,4);
TASK_PP(16'h1BF61,4);
TASK_PP(16'h1BF62,4);
TASK_PP(16'h1BF63,4);
TASK_PP(16'h1BF64,4);
TASK_PP(16'h1BF65,4);
TASK_PP(16'h1BF66,4);
TASK_PP(16'h1BF67,4);
TASK_PP(16'h1BF68,4);
TASK_PP(16'h1BF69,4);
TASK_PP(16'h1BF6A,4);
TASK_PP(16'h1BF6B,4);
TASK_PP(16'h1BF6C,4);
TASK_PP(16'h1BF6D,4);
TASK_PP(16'h1BF6E,4);
TASK_PP(16'h1BF6F,4);
TASK_PP(16'h1BF70,4);
TASK_PP(16'h1BF71,4);
TASK_PP(16'h1BF72,4);
TASK_PP(16'h1BF73,4);
TASK_PP(16'h1BF74,4);
TASK_PP(16'h1BF75,4);
TASK_PP(16'h1BF76,4);
TASK_PP(16'h1BF77,4);
TASK_PP(16'h1BF78,4);
TASK_PP(16'h1BF79,4);
TASK_PP(16'h1BF7A,4);
TASK_PP(16'h1BF7B,4);
TASK_PP(16'h1BF7C,4);
TASK_PP(16'h1BF7D,4);
TASK_PP(16'h1BF7E,4);
TASK_PP(16'h1BF7F,4);
TASK_PP(16'h1BF80,4);
TASK_PP(16'h1BF81,4);
TASK_PP(16'h1BF82,4);
TASK_PP(16'h1BF83,4);
TASK_PP(16'h1BF84,4);
TASK_PP(16'h1BF85,4);
TASK_PP(16'h1BF86,4);
TASK_PP(16'h1BF87,4);
TASK_PP(16'h1BF88,4);
TASK_PP(16'h1BF89,4);
TASK_PP(16'h1BF8A,4);
TASK_PP(16'h1BF8B,4);
TASK_PP(16'h1BF8C,4);
TASK_PP(16'h1BF8D,4);
TASK_PP(16'h1BF8E,4);
TASK_PP(16'h1BF8F,4);
TASK_PP(16'h1BF90,4);
TASK_PP(16'h1BF91,4);
TASK_PP(16'h1BF92,4);
TASK_PP(16'h1BF93,4);
TASK_PP(16'h1BF94,4);
TASK_PP(16'h1BF95,4);
TASK_PP(16'h1BF96,4);
TASK_PP(16'h1BF97,4);
TASK_PP(16'h1BF98,4);
TASK_PP(16'h1BF99,4);
TASK_PP(16'h1BF9A,4);
TASK_PP(16'h1BF9B,4);
TASK_PP(16'h1BF9C,4);
TASK_PP(16'h1BF9D,4);
TASK_PP(16'h1BF9E,4);
TASK_PP(16'h1BF9F,4);
TASK_PP(16'h1BFA0,4);
TASK_PP(16'h1BFA1,4);
TASK_PP(16'h1BFA2,4);
TASK_PP(16'h1BFA3,4);
TASK_PP(16'h1BFA4,4);
TASK_PP(16'h1BFA5,4);
TASK_PP(16'h1BFA6,4);
TASK_PP(16'h1BFA7,4);
TASK_PP(16'h1BFA8,4);
TASK_PP(16'h1BFA9,4);
TASK_PP(16'h1BFAA,4);
TASK_PP(16'h1BFAB,4);
TASK_PP(16'h1BFAC,4);
TASK_PP(16'h1BFAD,4);
TASK_PP(16'h1BFAE,4);
TASK_PP(16'h1BFAF,4);
TASK_PP(16'h1BFB0,4);
TASK_PP(16'h1BFB1,4);
TASK_PP(16'h1BFB2,4);
TASK_PP(16'h1BFB3,4);
TASK_PP(16'h1BFB4,4);
TASK_PP(16'h1BFB5,4);
TASK_PP(16'h1BFB6,4);
TASK_PP(16'h1BFB7,4);
TASK_PP(16'h1BFB8,4);
TASK_PP(16'h1BFB9,4);
TASK_PP(16'h1BFBA,4);
TASK_PP(16'h1BFBB,4);
TASK_PP(16'h1BFBC,4);
TASK_PP(16'h1BFBD,4);
TASK_PP(16'h1BFBE,4);
TASK_PP(16'h1BFBF,4);
TASK_PP(16'h1BFC0,4);
TASK_PP(16'h1BFC1,4);
TASK_PP(16'h1BFC2,4);
TASK_PP(16'h1BFC3,4);
TASK_PP(16'h1BFC4,4);
TASK_PP(16'h1BFC5,4);
TASK_PP(16'h1BFC6,4);
TASK_PP(16'h1BFC7,4);
TASK_PP(16'h1BFC8,4);
TASK_PP(16'h1BFC9,4);
TASK_PP(16'h1BFCA,4);
TASK_PP(16'h1BFCB,4);
TASK_PP(16'h1BFCC,4);
TASK_PP(16'h1BFCD,4);
TASK_PP(16'h1BFCE,4);
TASK_PP(16'h1BFCF,4);
TASK_PP(16'h1BFD0,4);
TASK_PP(16'h1BFD1,4);
TASK_PP(16'h1BFD2,4);
TASK_PP(16'h1BFD3,4);
TASK_PP(16'h1BFD4,4);
TASK_PP(16'h1BFD5,4);
TASK_PP(16'h1BFD6,4);
TASK_PP(16'h1BFD7,4);
TASK_PP(16'h1BFD8,4);
TASK_PP(16'h1BFD9,4);
TASK_PP(16'h1BFDA,4);
TASK_PP(16'h1BFDB,4);
TASK_PP(16'h1BFDC,4);
TASK_PP(16'h1BFDD,4);
TASK_PP(16'h1BFDE,4);
TASK_PP(16'h1BFDF,4);
TASK_PP(16'h1BFE0,4);
TASK_PP(16'h1BFE1,4);
TASK_PP(16'h1BFE2,4);
TASK_PP(16'h1BFE3,4);
TASK_PP(16'h1BFE4,4);
TASK_PP(16'h1BFE5,4);
TASK_PP(16'h1BFE6,4);
TASK_PP(16'h1BFE7,4);
TASK_PP(16'h1BFE8,4);
TASK_PP(16'h1BFE9,4);
TASK_PP(16'h1BFEA,4);
TASK_PP(16'h1BFEB,4);
TASK_PP(16'h1BFEC,4);
TASK_PP(16'h1BFED,4);
TASK_PP(16'h1BFEE,4);
TASK_PP(16'h1BFEF,4);
TASK_PP(16'h1BFF0,4);
TASK_PP(16'h1BFF1,4);
TASK_PP(16'h1BFF2,4);
TASK_PP(16'h1BFF3,4);
TASK_PP(16'h1BFF4,4);
TASK_PP(16'h1BFF5,4);
TASK_PP(16'h1BFF6,4);
TASK_PP(16'h1BFF7,4);
TASK_PP(16'h1BFF8,4);
TASK_PP(16'h1BFF9,4);
TASK_PP(16'h1BFFA,4);
TASK_PP(16'h1BFFB,4);
TASK_PP(16'h1BFFC,4);
TASK_PP(16'h1BFFD,4);
TASK_PP(16'h1BFFE,4);
TASK_PP(16'h1BFFF,4);
TASK_PP(16'h1C000,4);
TASK_PP(16'h1C001,4);
TASK_PP(16'h1C002,4);
TASK_PP(16'h1C003,4);
TASK_PP(16'h1C004,4);
TASK_PP(16'h1C005,4);
TASK_PP(16'h1C006,4);
TASK_PP(16'h1C007,4);
TASK_PP(16'h1C008,4);
TASK_PP(16'h1C009,4);
TASK_PP(16'h1C00A,4);
TASK_PP(16'h1C00B,4);
TASK_PP(16'h1C00C,4);
TASK_PP(16'h1C00D,4);
TASK_PP(16'h1C00E,4);
TASK_PP(16'h1C00F,4);
TASK_PP(16'h1C010,4);
TASK_PP(16'h1C011,4);
TASK_PP(16'h1C012,4);
TASK_PP(16'h1C013,4);
TASK_PP(16'h1C014,4);
TASK_PP(16'h1C015,4);
TASK_PP(16'h1C016,4);
TASK_PP(16'h1C017,4);
TASK_PP(16'h1C018,4);
TASK_PP(16'h1C019,4);
TASK_PP(16'h1C01A,4);
TASK_PP(16'h1C01B,4);
TASK_PP(16'h1C01C,4);
TASK_PP(16'h1C01D,4);
TASK_PP(16'h1C01E,4);
TASK_PP(16'h1C01F,4);
TASK_PP(16'h1C020,4);
TASK_PP(16'h1C021,4);
TASK_PP(16'h1C022,4);
TASK_PP(16'h1C023,4);
TASK_PP(16'h1C024,4);
TASK_PP(16'h1C025,4);
TASK_PP(16'h1C026,4);
TASK_PP(16'h1C027,4);
TASK_PP(16'h1C028,4);
TASK_PP(16'h1C029,4);
TASK_PP(16'h1C02A,4);
TASK_PP(16'h1C02B,4);
TASK_PP(16'h1C02C,4);
TASK_PP(16'h1C02D,4);
TASK_PP(16'h1C02E,4);
TASK_PP(16'h1C02F,4);
TASK_PP(16'h1C030,4);
TASK_PP(16'h1C031,4);
TASK_PP(16'h1C032,4);
TASK_PP(16'h1C033,4);
TASK_PP(16'h1C034,4);
TASK_PP(16'h1C035,4);
TASK_PP(16'h1C036,4);
TASK_PP(16'h1C037,4);
TASK_PP(16'h1C038,4);
TASK_PP(16'h1C039,4);
TASK_PP(16'h1C03A,4);
TASK_PP(16'h1C03B,4);
TASK_PP(16'h1C03C,4);
TASK_PP(16'h1C03D,4);
TASK_PP(16'h1C03E,4);
TASK_PP(16'h1C03F,4);
TASK_PP(16'h1C040,4);
TASK_PP(16'h1C041,4);
TASK_PP(16'h1C042,4);
TASK_PP(16'h1C043,4);
TASK_PP(16'h1C044,4);
TASK_PP(16'h1C045,4);
TASK_PP(16'h1C046,4);
TASK_PP(16'h1C047,4);
TASK_PP(16'h1C048,4);
TASK_PP(16'h1C049,4);
TASK_PP(16'h1C04A,4);
TASK_PP(16'h1C04B,4);
TASK_PP(16'h1C04C,4);
TASK_PP(16'h1C04D,4);
TASK_PP(16'h1C04E,4);
TASK_PP(16'h1C04F,4);
TASK_PP(16'h1C050,4);
TASK_PP(16'h1C051,4);
TASK_PP(16'h1C052,4);
TASK_PP(16'h1C053,4);
TASK_PP(16'h1C054,4);
TASK_PP(16'h1C055,4);
TASK_PP(16'h1C056,4);
TASK_PP(16'h1C057,4);
TASK_PP(16'h1C058,4);
TASK_PP(16'h1C059,4);
TASK_PP(16'h1C05A,4);
TASK_PP(16'h1C05B,4);
TASK_PP(16'h1C05C,4);
TASK_PP(16'h1C05D,4);
TASK_PP(16'h1C05E,4);
TASK_PP(16'h1C05F,4);
TASK_PP(16'h1C060,4);
TASK_PP(16'h1C061,4);
TASK_PP(16'h1C062,4);
TASK_PP(16'h1C063,4);
TASK_PP(16'h1C064,4);
TASK_PP(16'h1C065,4);
TASK_PP(16'h1C066,4);
TASK_PP(16'h1C067,4);
TASK_PP(16'h1C068,4);
TASK_PP(16'h1C069,4);
TASK_PP(16'h1C06A,4);
TASK_PP(16'h1C06B,4);
TASK_PP(16'h1C06C,4);
TASK_PP(16'h1C06D,4);
TASK_PP(16'h1C06E,4);
TASK_PP(16'h1C06F,4);
TASK_PP(16'h1C070,4);
TASK_PP(16'h1C071,4);
TASK_PP(16'h1C072,4);
TASK_PP(16'h1C073,4);
TASK_PP(16'h1C074,4);
TASK_PP(16'h1C075,4);
TASK_PP(16'h1C076,4);
TASK_PP(16'h1C077,4);
TASK_PP(16'h1C078,4);
TASK_PP(16'h1C079,4);
TASK_PP(16'h1C07A,4);
TASK_PP(16'h1C07B,4);
TASK_PP(16'h1C07C,4);
TASK_PP(16'h1C07D,4);
TASK_PP(16'h1C07E,4);
TASK_PP(16'h1C07F,4);
TASK_PP(16'h1C080,4);
TASK_PP(16'h1C081,4);
TASK_PP(16'h1C082,4);
TASK_PP(16'h1C083,4);
TASK_PP(16'h1C084,4);
TASK_PP(16'h1C085,4);
TASK_PP(16'h1C086,4);
TASK_PP(16'h1C087,4);
TASK_PP(16'h1C088,4);
TASK_PP(16'h1C089,4);
TASK_PP(16'h1C08A,4);
TASK_PP(16'h1C08B,4);
TASK_PP(16'h1C08C,4);
TASK_PP(16'h1C08D,4);
TASK_PP(16'h1C08E,4);
TASK_PP(16'h1C08F,4);
TASK_PP(16'h1C090,4);
TASK_PP(16'h1C091,4);
TASK_PP(16'h1C092,4);
TASK_PP(16'h1C093,4);
TASK_PP(16'h1C094,4);
TASK_PP(16'h1C095,4);
TASK_PP(16'h1C096,4);
TASK_PP(16'h1C097,4);
TASK_PP(16'h1C098,4);
TASK_PP(16'h1C099,4);
TASK_PP(16'h1C09A,4);
TASK_PP(16'h1C09B,4);
TASK_PP(16'h1C09C,4);
TASK_PP(16'h1C09D,4);
TASK_PP(16'h1C09E,4);
TASK_PP(16'h1C09F,4);
TASK_PP(16'h1C0A0,4);
TASK_PP(16'h1C0A1,4);
TASK_PP(16'h1C0A2,4);
TASK_PP(16'h1C0A3,4);
TASK_PP(16'h1C0A4,4);
TASK_PP(16'h1C0A5,4);
TASK_PP(16'h1C0A6,4);
TASK_PP(16'h1C0A7,4);
TASK_PP(16'h1C0A8,4);
TASK_PP(16'h1C0A9,4);
TASK_PP(16'h1C0AA,4);
TASK_PP(16'h1C0AB,4);
TASK_PP(16'h1C0AC,4);
TASK_PP(16'h1C0AD,4);
TASK_PP(16'h1C0AE,4);
TASK_PP(16'h1C0AF,4);
TASK_PP(16'h1C0B0,4);
TASK_PP(16'h1C0B1,4);
TASK_PP(16'h1C0B2,4);
TASK_PP(16'h1C0B3,4);
TASK_PP(16'h1C0B4,4);
TASK_PP(16'h1C0B5,4);
TASK_PP(16'h1C0B6,4);
TASK_PP(16'h1C0B7,4);
TASK_PP(16'h1C0B8,4);
TASK_PP(16'h1C0B9,4);
TASK_PP(16'h1C0BA,4);
TASK_PP(16'h1C0BB,4);
TASK_PP(16'h1C0BC,4);
TASK_PP(16'h1C0BD,4);
TASK_PP(16'h1C0BE,4);
TASK_PP(16'h1C0BF,4);
TASK_PP(16'h1C0C0,4);
TASK_PP(16'h1C0C1,4);
TASK_PP(16'h1C0C2,4);
TASK_PP(16'h1C0C3,4);
TASK_PP(16'h1C0C4,4);
TASK_PP(16'h1C0C5,4);
TASK_PP(16'h1C0C6,4);
TASK_PP(16'h1C0C7,4);
TASK_PP(16'h1C0C8,4);
TASK_PP(16'h1C0C9,4);
TASK_PP(16'h1C0CA,4);
TASK_PP(16'h1C0CB,4);
TASK_PP(16'h1C0CC,4);
TASK_PP(16'h1C0CD,4);
TASK_PP(16'h1C0CE,4);
TASK_PP(16'h1C0CF,4);
TASK_PP(16'h1C0D0,4);
TASK_PP(16'h1C0D1,4);
TASK_PP(16'h1C0D2,4);
TASK_PP(16'h1C0D3,4);
TASK_PP(16'h1C0D4,4);
TASK_PP(16'h1C0D5,4);
TASK_PP(16'h1C0D6,4);
TASK_PP(16'h1C0D7,4);
TASK_PP(16'h1C0D8,4);
TASK_PP(16'h1C0D9,4);
TASK_PP(16'h1C0DA,4);
TASK_PP(16'h1C0DB,4);
TASK_PP(16'h1C0DC,4);
TASK_PP(16'h1C0DD,4);
TASK_PP(16'h1C0DE,4);
TASK_PP(16'h1C0DF,4);
TASK_PP(16'h1C0E0,4);
TASK_PP(16'h1C0E1,4);
TASK_PP(16'h1C0E2,4);
TASK_PP(16'h1C0E3,4);
TASK_PP(16'h1C0E4,4);
TASK_PP(16'h1C0E5,4);
TASK_PP(16'h1C0E6,4);
TASK_PP(16'h1C0E7,4);
TASK_PP(16'h1C0E8,4);
TASK_PP(16'h1C0E9,4);
TASK_PP(16'h1C0EA,4);
TASK_PP(16'h1C0EB,4);
TASK_PP(16'h1C0EC,4);
TASK_PP(16'h1C0ED,4);
TASK_PP(16'h1C0EE,4);
TASK_PP(16'h1C0EF,4);
TASK_PP(16'h1C0F0,4);
TASK_PP(16'h1C0F1,4);
TASK_PP(16'h1C0F2,4);
TASK_PP(16'h1C0F3,4);
TASK_PP(16'h1C0F4,4);
TASK_PP(16'h1C0F5,4);
TASK_PP(16'h1C0F6,4);
TASK_PP(16'h1C0F7,4);
TASK_PP(16'h1C0F8,4);
TASK_PP(16'h1C0F9,4);
TASK_PP(16'h1C0FA,4);
TASK_PP(16'h1C0FB,4);
TASK_PP(16'h1C0FC,4);
TASK_PP(16'h1C0FD,4);
TASK_PP(16'h1C0FE,4);
TASK_PP(16'h1C0FF,4);
TASK_PP(16'h1C100,4);
TASK_PP(16'h1C101,4);
TASK_PP(16'h1C102,4);
TASK_PP(16'h1C103,4);
TASK_PP(16'h1C104,4);
TASK_PP(16'h1C105,4);
TASK_PP(16'h1C106,4);
TASK_PP(16'h1C107,4);
TASK_PP(16'h1C108,4);
TASK_PP(16'h1C109,4);
TASK_PP(16'h1C10A,4);
TASK_PP(16'h1C10B,4);
TASK_PP(16'h1C10C,4);
TASK_PP(16'h1C10D,4);
TASK_PP(16'h1C10E,4);
TASK_PP(16'h1C10F,4);
TASK_PP(16'h1C110,4);
TASK_PP(16'h1C111,4);
TASK_PP(16'h1C112,4);
TASK_PP(16'h1C113,4);
TASK_PP(16'h1C114,4);
TASK_PP(16'h1C115,4);
TASK_PP(16'h1C116,4);
TASK_PP(16'h1C117,4);
TASK_PP(16'h1C118,4);
TASK_PP(16'h1C119,4);
TASK_PP(16'h1C11A,4);
TASK_PP(16'h1C11B,4);
TASK_PP(16'h1C11C,4);
TASK_PP(16'h1C11D,4);
TASK_PP(16'h1C11E,4);
TASK_PP(16'h1C11F,4);
TASK_PP(16'h1C120,4);
TASK_PP(16'h1C121,4);
TASK_PP(16'h1C122,4);
TASK_PP(16'h1C123,4);
TASK_PP(16'h1C124,4);
TASK_PP(16'h1C125,4);
TASK_PP(16'h1C126,4);
TASK_PP(16'h1C127,4);
TASK_PP(16'h1C128,4);
TASK_PP(16'h1C129,4);
TASK_PP(16'h1C12A,4);
TASK_PP(16'h1C12B,4);
TASK_PP(16'h1C12C,4);
TASK_PP(16'h1C12D,4);
TASK_PP(16'h1C12E,4);
TASK_PP(16'h1C12F,4);
TASK_PP(16'h1C130,4);
TASK_PP(16'h1C131,4);
TASK_PP(16'h1C132,4);
TASK_PP(16'h1C133,4);
TASK_PP(16'h1C134,4);
TASK_PP(16'h1C135,4);
TASK_PP(16'h1C136,4);
TASK_PP(16'h1C137,4);
TASK_PP(16'h1C138,4);
TASK_PP(16'h1C139,4);
TASK_PP(16'h1C13A,4);
TASK_PP(16'h1C13B,4);
TASK_PP(16'h1C13C,4);
TASK_PP(16'h1C13D,4);
TASK_PP(16'h1C13E,4);
TASK_PP(16'h1C13F,4);
TASK_PP(16'h1C140,4);
TASK_PP(16'h1C141,4);
TASK_PP(16'h1C142,4);
TASK_PP(16'h1C143,4);
TASK_PP(16'h1C144,4);
TASK_PP(16'h1C145,4);
TASK_PP(16'h1C146,4);
TASK_PP(16'h1C147,4);
TASK_PP(16'h1C148,4);
TASK_PP(16'h1C149,4);
TASK_PP(16'h1C14A,4);
TASK_PP(16'h1C14B,4);
TASK_PP(16'h1C14C,4);
TASK_PP(16'h1C14D,4);
TASK_PP(16'h1C14E,4);
TASK_PP(16'h1C14F,4);
TASK_PP(16'h1C150,4);
TASK_PP(16'h1C151,4);
TASK_PP(16'h1C152,4);
TASK_PP(16'h1C153,4);
TASK_PP(16'h1C154,4);
TASK_PP(16'h1C155,4);
TASK_PP(16'h1C156,4);
TASK_PP(16'h1C157,4);
TASK_PP(16'h1C158,4);
TASK_PP(16'h1C159,4);
TASK_PP(16'h1C15A,4);
TASK_PP(16'h1C15B,4);
TASK_PP(16'h1C15C,4);
TASK_PP(16'h1C15D,4);
TASK_PP(16'h1C15E,4);
TASK_PP(16'h1C15F,4);
TASK_PP(16'h1C160,4);
TASK_PP(16'h1C161,4);
TASK_PP(16'h1C162,4);
TASK_PP(16'h1C163,4);
TASK_PP(16'h1C164,4);
TASK_PP(16'h1C165,4);
TASK_PP(16'h1C166,4);
TASK_PP(16'h1C167,4);
TASK_PP(16'h1C168,4);
TASK_PP(16'h1C169,4);
TASK_PP(16'h1C16A,4);
TASK_PP(16'h1C16B,4);
TASK_PP(16'h1C16C,4);
TASK_PP(16'h1C16D,4);
TASK_PP(16'h1C16E,4);
TASK_PP(16'h1C16F,4);
TASK_PP(16'h1C170,4);
TASK_PP(16'h1C171,4);
TASK_PP(16'h1C172,4);
TASK_PP(16'h1C173,4);
TASK_PP(16'h1C174,4);
TASK_PP(16'h1C175,4);
TASK_PP(16'h1C176,4);
TASK_PP(16'h1C177,4);
TASK_PP(16'h1C178,4);
TASK_PP(16'h1C179,4);
TASK_PP(16'h1C17A,4);
TASK_PP(16'h1C17B,4);
TASK_PP(16'h1C17C,4);
TASK_PP(16'h1C17D,4);
TASK_PP(16'h1C17E,4);
TASK_PP(16'h1C17F,4);
TASK_PP(16'h1C180,4);
TASK_PP(16'h1C181,4);
TASK_PP(16'h1C182,4);
TASK_PP(16'h1C183,4);
TASK_PP(16'h1C184,4);
TASK_PP(16'h1C185,4);
TASK_PP(16'h1C186,4);
TASK_PP(16'h1C187,4);
TASK_PP(16'h1C188,4);
TASK_PP(16'h1C189,4);
TASK_PP(16'h1C18A,4);
TASK_PP(16'h1C18B,4);
TASK_PP(16'h1C18C,4);
TASK_PP(16'h1C18D,4);
TASK_PP(16'h1C18E,4);
TASK_PP(16'h1C18F,4);
TASK_PP(16'h1C190,4);
TASK_PP(16'h1C191,4);
TASK_PP(16'h1C192,4);
TASK_PP(16'h1C193,4);
TASK_PP(16'h1C194,4);
TASK_PP(16'h1C195,4);
TASK_PP(16'h1C196,4);
TASK_PP(16'h1C197,4);
TASK_PP(16'h1C198,4);
TASK_PP(16'h1C199,4);
TASK_PP(16'h1C19A,4);
TASK_PP(16'h1C19B,4);
TASK_PP(16'h1C19C,4);
TASK_PP(16'h1C19D,4);
TASK_PP(16'h1C19E,4);
TASK_PP(16'h1C19F,4);
TASK_PP(16'h1C1A0,4);
TASK_PP(16'h1C1A1,4);
TASK_PP(16'h1C1A2,4);
TASK_PP(16'h1C1A3,4);
TASK_PP(16'h1C1A4,4);
TASK_PP(16'h1C1A5,4);
TASK_PP(16'h1C1A6,4);
TASK_PP(16'h1C1A7,4);
TASK_PP(16'h1C1A8,4);
TASK_PP(16'h1C1A9,4);
TASK_PP(16'h1C1AA,4);
TASK_PP(16'h1C1AB,4);
TASK_PP(16'h1C1AC,4);
TASK_PP(16'h1C1AD,4);
TASK_PP(16'h1C1AE,4);
TASK_PP(16'h1C1AF,4);
TASK_PP(16'h1C1B0,4);
TASK_PP(16'h1C1B1,4);
TASK_PP(16'h1C1B2,4);
TASK_PP(16'h1C1B3,4);
TASK_PP(16'h1C1B4,4);
TASK_PP(16'h1C1B5,4);
TASK_PP(16'h1C1B6,4);
TASK_PP(16'h1C1B7,4);
TASK_PP(16'h1C1B8,4);
TASK_PP(16'h1C1B9,4);
TASK_PP(16'h1C1BA,4);
TASK_PP(16'h1C1BB,4);
TASK_PP(16'h1C1BC,4);
TASK_PP(16'h1C1BD,4);
TASK_PP(16'h1C1BE,4);
TASK_PP(16'h1C1BF,4);
TASK_PP(16'h1C1C0,4);
TASK_PP(16'h1C1C1,4);
TASK_PP(16'h1C1C2,4);
TASK_PP(16'h1C1C3,4);
TASK_PP(16'h1C1C4,4);
TASK_PP(16'h1C1C5,4);
TASK_PP(16'h1C1C6,4);
TASK_PP(16'h1C1C7,4);
TASK_PP(16'h1C1C8,4);
TASK_PP(16'h1C1C9,4);
TASK_PP(16'h1C1CA,4);
TASK_PP(16'h1C1CB,4);
TASK_PP(16'h1C1CC,4);
TASK_PP(16'h1C1CD,4);
TASK_PP(16'h1C1CE,4);
TASK_PP(16'h1C1CF,4);
TASK_PP(16'h1C1D0,4);
TASK_PP(16'h1C1D1,4);
TASK_PP(16'h1C1D2,4);
TASK_PP(16'h1C1D3,4);
TASK_PP(16'h1C1D4,4);
TASK_PP(16'h1C1D5,4);
TASK_PP(16'h1C1D6,4);
TASK_PP(16'h1C1D7,4);
TASK_PP(16'h1C1D8,4);
TASK_PP(16'h1C1D9,4);
TASK_PP(16'h1C1DA,4);
TASK_PP(16'h1C1DB,4);
TASK_PP(16'h1C1DC,4);
TASK_PP(16'h1C1DD,4);
TASK_PP(16'h1C1DE,4);
TASK_PP(16'h1C1DF,4);
TASK_PP(16'h1C1E0,4);
TASK_PP(16'h1C1E1,4);
TASK_PP(16'h1C1E2,4);
TASK_PP(16'h1C1E3,4);
TASK_PP(16'h1C1E4,4);
TASK_PP(16'h1C1E5,4);
TASK_PP(16'h1C1E6,4);
TASK_PP(16'h1C1E7,4);
TASK_PP(16'h1C1E8,4);
TASK_PP(16'h1C1E9,4);
TASK_PP(16'h1C1EA,4);
TASK_PP(16'h1C1EB,4);
TASK_PP(16'h1C1EC,4);
TASK_PP(16'h1C1ED,4);
TASK_PP(16'h1C1EE,4);
TASK_PP(16'h1C1EF,4);
TASK_PP(16'h1C1F0,4);
TASK_PP(16'h1C1F1,4);
TASK_PP(16'h1C1F2,4);
TASK_PP(16'h1C1F3,4);
TASK_PP(16'h1C1F4,4);
TASK_PP(16'h1C1F5,4);
TASK_PP(16'h1C1F6,4);
TASK_PP(16'h1C1F7,4);
TASK_PP(16'h1C1F8,4);
TASK_PP(16'h1C1F9,4);
TASK_PP(16'h1C1FA,4);
TASK_PP(16'h1C1FB,4);
TASK_PP(16'h1C1FC,4);
TASK_PP(16'h1C1FD,4);
TASK_PP(16'h1C1FE,4);
TASK_PP(16'h1C1FF,4);
TASK_PP(16'h1C200,4);
TASK_PP(16'h1C201,4);
TASK_PP(16'h1C202,4);
TASK_PP(16'h1C203,4);
TASK_PP(16'h1C204,4);
TASK_PP(16'h1C205,4);
TASK_PP(16'h1C206,4);
TASK_PP(16'h1C207,4);
TASK_PP(16'h1C208,4);
TASK_PP(16'h1C209,4);
TASK_PP(16'h1C20A,4);
TASK_PP(16'h1C20B,4);
TASK_PP(16'h1C20C,4);
TASK_PP(16'h1C20D,4);
TASK_PP(16'h1C20E,4);
TASK_PP(16'h1C20F,4);
TASK_PP(16'h1C210,4);
TASK_PP(16'h1C211,4);
TASK_PP(16'h1C212,4);
TASK_PP(16'h1C213,4);
TASK_PP(16'h1C214,4);
TASK_PP(16'h1C215,4);
TASK_PP(16'h1C216,4);
TASK_PP(16'h1C217,4);
TASK_PP(16'h1C218,4);
TASK_PP(16'h1C219,4);
TASK_PP(16'h1C21A,4);
TASK_PP(16'h1C21B,4);
TASK_PP(16'h1C21C,4);
TASK_PP(16'h1C21D,4);
TASK_PP(16'h1C21E,4);
TASK_PP(16'h1C21F,4);
TASK_PP(16'h1C220,4);
TASK_PP(16'h1C221,4);
TASK_PP(16'h1C222,4);
TASK_PP(16'h1C223,4);
TASK_PP(16'h1C224,4);
TASK_PP(16'h1C225,4);
TASK_PP(16'h1C226,4);
TASK_PP(16'h1C227,4);
TASK_PP(16'h1C228,4);
TASK_PP(16'h1C229,4);
TASK_PP(16'h1C22A,4);
TASK_PP(16'h1C22B,4);
TASK_PP(16'h1C22C,4);
TASK_PP(16'h1C22D,4);
TASK_PP(16'h1C22E,4);
TASK_PP(16'h1C22F,4);
TASK_PP(16'h1C230,4);
TASK_PP(16'h1C231,4);
TASK_PP(16'h1C232,4);
TASK_PP(16'h1C233,4);
TASK_PP(16'h1C234,4);
TASK_PP(16'h1C235,4);
TASK_PP(16'h1C236,4);
TASK_PP(16'h1C237,4);
TASK_PP(16'h1C238,4);
TASK_PP(16'h1C239,4);
TASK_PP(16'h1C23A,4);
TASK_PP(16'h1C23B,4);
TASK_PP(16'h1C23C,4);
TASK_PP(16'h1C23D,4);
TASK_PP(16'h1C23E,4);
TASK_PP(16'h1C23F,4);
TASK_PP(16'h1C240,4);
TASK_PP(16'h1C241,4);
TASK_PP(16'h1C242,4);
TASK_PP(16'h1C243,4);
TASK_PP(16'h1C244,4);
TASK_PP(16'h1C245,4);
TASK_PP(16'h1C246,4);
TASK_PP(16'h1C247,4);
TASK_PP(16'h1C248,4);
TASK_PP(16'h1C249,4);
TASK_PP(16'h1C24A,4);
TASK_PP(16'h1C24B,4);
TASK_PP(16'h1C24C,4);
TASK_PP(16'h1C24D,4);
TASK_PP(16'h1C24E,4);
TASK_PP(16'h1C24F,4);
TASK_PP(16'h1C250,4);
TASK_PP(16'h1C251,4);
TASK_PP(16'h1C252,4);
TASK_PP(16'h1C253,4);
TASK_PP(16'h1C254,4);
TASK_PP(16'h1C255,4);
TASK_PP(16'h1C256,4);
TASK_PP(16'h1C257,4);
TASK_PP(16'h1C258,4);
TASK_PP(16'h1C259,4);
TASK_PP(16'h1C25A,4);
TASK_PP(16'h1C25B,4);
TASK_PP(16'h1C25C,4);
TASK_PP(16'h1C25D,4);
TASK_PP(16'h1C25E,4);
TASK_PP(16'h1C25F,4);
TASK_PP(16'h1C260,4);
TASK_PP(16'h1C261,4);
TASK_PP(16'h1C262,4);
TASK_PP(16'h1C263,4);
TASK_PP(16'h1C264,4);
TASK_PP(16'h1C265,4);
TASK_PP(16'h1C266,4);
TASK_PP(16'h1C267,4);
TASK_PP(16'h1C268,4);
TASK_PP(16'h1C269,4);
TASK_PP(16'h1C26A,4);
TASK_PP(16'h1C26B,4);
TASK_PP(16'h1C26C,4);
TASK_PP(16'h1C26D,4);
TASK_PP(16'h1C26E,4);
TASK_PP(16'h1C26F,4);
TASK_PP(16'h1C270,4);
TASK_PP(16'h1C271,4);
TASK_PP(16'h1C272,4);
TASK_PP(16'h1C273,4);
TASK_PP(16'h1C274,4);
TASK_PP(16'h1C275,4);
TASK_PP(16'h1C276,4);
TASK_PP(16'h1C277,4);
TASK_PP(16'h1C278,4);
TASK_PP(16'h1C279,4);
TASK_PP(16'h1C27A,4);
TASK_PP(16'h1C27B,4);
TASK_PP(16'h1C27C,4);
TASK_PP(16'h1C27D,4);
TASK_PP(16'h1C27E,4);
TASK_PP(16'h1C27F,4);
TASK_PP(16'h1C280,4);
TASK_PP(16'h1C281,4);
TASK_PP(16'h1C282,4);
TASK_PP(16'h1C283,4);
TASK_PP(16'h1C284,4);
TASK_PP(16'h1C285,4);
TASK_PP(16'h1C286,4);
TASK_PP(16'h1C287,4);
TASK_PP(16'h1C288,4);
TASK_PP(16'h1C289,4);
TASK_PP(16'h1C28A,4);
TASK_PP(16'h1C28B,4);
TASK_PP(16'h1C28C,4);
TASK_PP(16'h1C28D,4);
TASK_PP(16'h1C28E,4);
TASK_PP(16'h1C28F,4);
TASK_PP(16'h1C290,4);
TASK_PP(16'h1C291,4);
TASK_PP(16'h1C292,4);
TASK_PP(16'h1C293,4);
TASK_PP(16'h1C294,4);
TASK_PP(16'h1C295,4);
TASK_PP(16'h1C296,4);
TASK_PP(16'h1C297,4);
TASK_PP(16'h1C298,4);
TASK_PP(16'h1C299,4);
TASK_PP(16'h1C29A,4);
TASK_PP(16'h1C29B,4);
TASK_PP(16'h1C29C,4);
TASK_PP(16'h1C29D,4);
TASK_PP(16'h1C29E,4);
TASK_PP(16'h1C29F,4);
TASK_PP(16'h1C2A0,4);
TASK_PP(16'h1C2A1,4);
TASK_PP(16'h1C2A2,4);
TASK_PP(16'h1C2A3,4);
TASK_PP(16'h1C2A4,4);
TASK_PP(16'h1C2A5,4);
TASK_PP(16'h1C2A6,4);
TASK_PP(16'h1C2A7,4);
TASK_PP(16'h1C2A8,4);
TASK_PP(16'h1C2A9,4);
TASK_PP(16'h1C2AA,4);
TASK_PP(16'h1C2AB,4);
TASK_PP(16'h1C2AC,4);
TASK_PP(16'h1C2AD,4);
TASK_PP(16'h1C2AE,4);
TASK_PP(16'h1C2AF,4);
TASK_PP(16'h1C2B0,4);
TASK_PP(16'h1C2B1,4);
TASK_PP(16'h1C2B2,4);
TASK_PP(16'h1C2B3,4);
TASK_PP(16'h1C2B4,4);
TASK_PP(16'h1C2B5,4);
TASK_PP(16'h1C2B6,4);
TASK_PP(16'h1C2B7,4);
TASK_PP(16'h1C2B8,4);
TASK_PP(16'h1C2B9,4);
TASK_PP(16'h1C2BA,4);
TASK_PP(16'h1C2BB,4);
TASK_PP(16'h1C2BC,4);
TASK_PP(16'h1C2BD,4);
TASK_PP(16'h1C2BE,4);
TASK_PP(16'h1C2BF,4);
TASK_PP(16'h1C2C0,4);
TASK_PP(16'h1C2C1,4);
TASK_PP(16'h1C2C2,4);
TASK_PP(16'h1C2C3,4);
TASK_PP(16'h1C2C4,4);
TASK_PP(16'h1C2C5,4);
TASK_PP(16'h1C2C6,4);
TASK_PP(16'h1C2C7,4);
TASK_PP(16'h1C2C8,4);
TASK_PP(16'h1C2C9,4);
TASK_PP(16'h1C2CA,4);
TASK_PP(16'h1C2CB,4);
TASK_PP(16'h1C2CC,4);
TASK_PP(16'h1C2CD,4);
TASK_PP(16'h1C2CE,4);
TASK_PP(16'h1C2CF,4);
TASK_PP(16'h1C2D0,4);
TASK_PP(16'h1C2D1,4);
TASK_PP(16'h1C2D2,4);
TASK_PP(16'h1C2D3,4);
TASK_PP(16'h1C2D4,4);
TASK_PP(16'h1C2D5,4);
TASK_PP(16'h1C2D6,4);
TASK_PP(16'h1C2D7,4);
TASK_PP(16'h1C2D8,4);
TASK_PP(16'h1C2D9,4);
TASK_PP(16'h1C2DA,4);
TASK_PP(16'h1C2DB,4);
TASK_PP(16'h1C2DC,4);
TASK_PP(16'h1C2DD,4);
TASK_PP(16'h1C2DE,4);
TASK_PP(16'h1C2DF,4);
TASK_PP(16'h1C2E0,4);
TASK_PP(16'h1C2E1,4);
TASK_PP(16'h1C2E2,4);
TASK_PP(16'h1C2E3,4);
TASK_PP(16'h1C2E4,4);
TASK_PP(16'h1C2E5,4);
TASK_PP(16'h1C2E6,4);
TASK_PP(16'h1C2E7,4);
TASK_PP(16'h1C2E8,4);
TASK_PP(16'h1C2E9,4);
TASK_PP(16'h1C2EA,4);
TASK_PP(16'h1C2EB,4);
TASK_PP(16'h1C2EC,4);
TASK_PP(16'h1C2ED,4);
TASK_PP(16'h1C2EE,4);
TASK_PP(16'h1C2EF,4);
TASK_PP(16'h1C2F0,4);
TASK_PP(16'h1C2F1,4);
TASK_PP(16'h1C2F2,4);
TASK_PP(16'h1C2F3,4);
TASK_PP(16'h1C2F4,4);
TASK_PP(16'h1C2F5,4);
TASK_PP(16'h1C2F6,4);
TASK_PP(16'h1C2F7,4);
TASK_PP(16'h1C2F8,4);
TASK_PP(16'h1C2F9,4);
TASK_PP(16'h1C2FA,4);
TASK_PP(16'h1C2FB,4);
TASK_PP(16'h1C2FC,4);
TASK_PP(16'h1C2FD,4);
TASK_PP(16'h1C2FE,4);
TASK_PP(16'h1C2FF,4);
TASK_PP(16'h1C300,4);
TASK_PP(16'h1C301,4);
TASK_PP(16'h1C302,4);
TASK_PP(16'h1C303,4);
TASK_PP(16'h1C304,4);
TASK_PP(16'h1C305,4);
TASK_PP(16'h1C306,4);
TASK_PP(16'h1C307,4);
TASK_PP(16'h1C308,4);
TASK_PP(16'h1C309,4);
TASK_PP(16'h1C30A,4);
TASK_PP(16'h1C30B,4);
TASK_PP(16'h1C30C,4);
TASK_PP(16'h1C30D,4);
TASK_PP(16'h1C30E,4);
TASK_PP(16'h1C30F,4);
TASK_PP(16'h1C310,4);
TASK_PP(16'h1C311,4);
TASK_PP(16'h1C312,4);
TASK_PP(16'h1C313,4);
TASK_PP(16'h1C314,4);
TASK_PP(16'h1C315,4);
TASK_PP(16'h1C316,4);
TASK_PP(16'h1C317,4);
TASK_PP(16'h1C318,4);
TASK_PP(16'h1C319,4);
TASK_PP(16'h1C31A,4);
TASK_PP(16'h1C31B,4);
TASK_PP(16'h1C31C,4);
TASK_PP(16'h1C31D,4);
TASK_PP(16'h1C31E,4);
TASK_PP(16'h1C31F,4);
TASK_PP(16'h1C320,4);
TASK_PP(16'h1C321,4);
TASK_PP(16'h1C322,4);
TASK_PP(16'h1C323,4);
TASK_PP(16'h1C324,4);
TASK_PP(16'h1C325,4);
TASK_PP(16'h1C326,4);
TASK_PP(16'h1C327,4);
TASK_PP(16'h1C328,4);
TASK_PP(16'h1C329,4);
TASK_PP(16'h1C32A,4);
TASK_PP(16'h1C32B,4);
TASK_PP(16'h1C32C,4);
TASK_PP(16'h1C32D,4);
TASK_PP(16'h1C32E,4);
TASK_PP(16'h1C32F,4);
TASK_PP(16'h1C330,4);
TASK_PP(16'h1C331,4);
TASK_PP(16'h1C332,4);
TASK_PP(16'h1C333,4);
TASK_PP(16'h1C334,4);
TASK_PP(16'h1C335,4);
TASK_PP(16'h1C336,4);
TASK_PP(16'h1C337,4);
TASK_PP(16'h1C338,4);
TASK_PP(16'h1C339,4);
TASK_PP(16'h1C33A,4);
TASK_PP(16'h1C33B,4);
TASK_PP(16'h1C33C,4);
TASK_PP(16'h1C33D,4);
TASK_PP(16'h1C33E,4);
TASK_PP(16'h1C33F,4);
TASK_PP(16'h1C340,4);
TASK_PP(16'h1C341,4);
TASK_PP(16'h1C342,4);
TASK_PP(16'h1C343,4);
TASK_PP(16'h1C344,4);
TASK_PP(16'h1C345,4);
TASK_PP(16'h1C346,4);
TASK_PP(16'h1C347,4);
TASK_PP(16'h1C348,4);
TASK_PP(16'h1C349,4);
TASK_PP(16'h1C34A,4);
TASK_PP(16'h1C34B,4);
TASK_PP(16'h1C34C,4);
TASK_PP(16'h1C34D,4);
TASK_PP(16'h1C34E,4);
TASK_PP(16'h1C34F,4);
TASK_PP(16'h1C350,4);
TASK_PP(16'h1C351,4);
TASK_PP(16'h1C352,4);
TASK_PP(16'h1C353,4);
TASK_PP(16'h1C354,4);
TASK_PP(16'h1C355,4);
TASK_PP(16'h1C356,4);
TASK_PP(16'h1C357,4);
TASK_PP(16'h1C358,4);
TASK_PP(16'h1C359,4);
TASK_PP(16'h1C35A,4);
TASK_PP(16'h1C35B,4);
TASK_PP(16'h1C35C,4);
TASK_PP(16'h1C35D,4);
TASK_PP(16'h1C35E,4);
TASK_PP(16'h1C35F,4);
TASK_PP(16'h1C360,4);
TASK_PP(16'h1C361,4);
TASK_PP(16'h1C362,4);
TASK_PP(16'h1C363,4);
TASK_PP(16'h1C364,4);
TASK_PP(16'h1C365,4);
TASK_PP(16'h1C366,4);
TASK_PP(16'h1C367,4);
TASK_PP(16'h1C368,4);
TASK_PP(16'h1C369,4);
TASK_PP(16'h1C36A,4);
TASK_PP(16'h1C36B,4);
TASK_PP(16'h1C36C,4);
TASK_PP(16'h1C36D,4);
TASK_PP(16'h1C36E,4);
TASK_PP(16'h1C36F,4);
TASK_PP(16'h1C370,4);
TASK_PP(16'h1C371,4);
TASK_PP(16'h1C372,4);
TASK_PP(16'h1C373,4);
TASK_PP(16'h1C374,4);
TASK_PP(16'h1C375,4);
TASK_PP(16'h1C376,4);
TASK_PP(16'h1C377,4);
TASK_PP(16'h1C378,4);
TASK_PP(16'h1C379,4);
TASK_PP(16'h1C37A,4);
TASK_PP(16'h1C37B,4);
TASK_PP(16'h1C37C,4);
TASK_PP(16'h1C37D,4);
TASK_PP(16'h1C37E,4);
TASK_PP(16'h1C37F,4);
TASK_PP(16'h1C380,4);
TASK_PP(16'h1C381,4);
TASK_PP(16'h1C382,4);
TASK_PP(16'h1C383,4);
TASK_PP(16'h1C384,4);
TASK_PP(16'h1C385,4);
TASK_PP(16'h1C386,4);
TASK_PP(16'h1C387,4);
TASK_PP(16'h1C388,4);
TASK_PP(16'h1C389,4);
TASK_PP(16'h1C38A,4);
TASK_PP(16'h1C38B,4);
TASK_PP(16'h1C38C,4);
TASK_PP(16'h1C38D,4);
TASK_PP(16'h1C38E,4);
TASK_PP(16'h1C38F,4);
TASK_PP(16'h1C390,4);
TASK_PP(16'h1C391,4);
TASK_PP(16'h1C392,4);
TASK_PP(16'h1C393,4);
TASK_PP(16'h1C394,4);
TASK_PP(16'h1C395,4);
TASK_PP(16'h1C396,4);
TASK_PP(16'h1C397,4);
TASK_PP(16'h1C398,4);
TASK_PP(16'h1C399,4);
TASK_PP(16'h1C39A,4);
TASK_PP(16'h1C39B,4);
TASK_PP(16'h1C39C,4);
TASK_PP(16'h1C39D,4);
TASK_PP(16'h1C39E,4);
TASK_PP(16'h1C39F,4);
TASK_PP(16'h1C3A0,4);
TASK_PP(16'h1C3A1,4);
TASK_PP(16'h1C3A2,4);
TASK_PP(16'h1C3A3,4);
TASK_PP(16'h1C3A4,4);
TASK_PP(16'h1C3A5,4);
TASK_PP(16'h1C3A6,4);
TASK_PP(16'h1C3A7,4);
TASK_PP(16'h1C3A8,4);
TASK_PP(16'h1C3A9,4);
TASK_PP(16'h1C3AA,4);
TASK_PP(16'h1C3AB,4);
TASK_PP(16'h1C3AC,4);
TASK_PP(16'h1C3AD,4);
TASK_PP(16'h1C3AE,4);
TASK_PP(16'h1C3AF,4);
TASK_PP(16'h1C3B0,4);
TASK_PP(16'h1C3B1,4);
TASK_PP(16'h1C3B2,4);
TASK_PP(16'h1C3B3,4);
TASK_PP(16'h1C3B4,4);
TASK_PP(16'h1C3B5,4);
TASK_PP(16'h1C3B6,4);
TASK_PP(16'h1C3B7,4);
TASK_PP(16'h1C3B8,4);
TASK_PP(16'h1C3B9,4);
TASK_PP(16'h1C3BA,4);
TASK_PP(16'h1C3BB,4);
TASK_PP(16'h1C3BC,4);
TASK_PP(16'h1C3BD,4);
TASK_PP(16'h1C3BE,4);
TASK_PP(16'h1C3BF,4);
TASK_PP(16'h1C3C0,4);
TASK_PP(16'h1C3C1,4);
TASK_PP(16'h1C3C2,4);
TASK_PP(16'h1C3C3,4);
TASK_PP(16'h1C3C4,4);
TASK_PP(16'h1C3C5,4);
TASK_PP(16'h1C3C6,4);
TASK_PP(16'h1C3C7,4);
TASK_PP(16'h1C3C8,4);
TASK_PP(16'h1C3C9,4);
TASK_PP(16'h1C3CA,4);
TASK_PP(16'h1C3CB,4);
TASK_PP(16'h1C3CC,4);
TASK_PP(16'h1C3CD,4);
TASK_PP(16'h1C3CE,4);
TASK_PP(16'h1C3CF,4);
TASK_PP(16'h1C3D0,4);
TASK_PP(16'h1C3D1,4);
TASK_PP(16'h1C3D2,4);
TASK_PP(16'h1C3D3,4);
TASK_PP(16'h1C3D4,4);
TASK_PP(16'h1C3D5,4);
TASK_PP(16'h1C3D6,4);
TASK_PP(16'h1C3D7,4);
TASK_PP(16'h1C3D8,4);
TASK_PP(16'h1C3D9,4);
TASK_PP(16'h1C3DA,4);
TASK_PP(16'h1C3DB,4);
TASK_PP(16'h1C3DC,4);
TASK_PP(16'h1C3DD,4);
TASK_PP(16'h1C3DE,4);
TASK_PP(16'h1C3DF,4);
TASK_PP(16'h1C3E0,4);
TASK_PP(16'h1C3E1,4);
TASK_PP(16'h1C3E2,4);
TASK_PP(16'h1C3E3,4);
TASK_PP(16'h1C3E4,4);
TASK_PP(16'h1C3E5,4);
TASK_PP(16'h1C3E6,4);
TASK_PP(16'h1C3E7,4);
TASK_PP(16'h1C3E8,4);
TASK_PP(16'h1C3E9,4);
TASK_PP(16'h1C3EA,4);
TASK_PP(16'h1C3EB,4);
TASK_PP(16'h1C3EC,4);
TASK_PP(16'h1C3ED,4);
TASK_PP(16'h1C3EE,4);
TASK_PP(16'h1C3EF,4);
TASK_PP(16'h1C3F0,4);
TASK_PP(16'h1C3F1,4);
TASK_PP(16'h1C3F2,4);
TASK_PP(16'h1C3F3,4);
TASK_PP(16'h1C3F4,4);
TASK_PP(16'h1C3F5,4);
TASK_PP(16'h1C3F6,4);
TASK_PP(16'h1C3F7,4);
TASK_PP(16'h1C3F8,4);
TASK_PP(16'h1C3F9,4);
TASK_PP(16'h1C3FA,4);
TASK_PP(16'h1C3FB,4);
TASK_PP(16'h1C3FC,4);
TASK_PP(16'h1C3FD,4);
TASK_PP(16'h1C3FE,4);
TASK_PP(16'h1C3FF,4);
TASK_PP(16'h1C400,4);
TASK_PP(16'h1C401,4);
TASK_PP(16'h1C402,4);
TASK_PP(16'h1C403,4);
TASK_PP(16'h1C404,4);
TASK_PP(16'h1C405,4);
TASK_PP(16'h1C406,4);
TASK_PP(16'h1C407,4);
TASK_PP(16'h1C408,4);
TASK_PP(16'h1C409,4);
TASK_PP(16'h1C40A,4);
TASK_PP(16'h1C40B,4);
TASK_PP(16'h1C40C,4);
TASK_PP(16'h1C40D,4);
TASK_PP(16'h1C40E,4);
TASK_PP(16'h1C40F,4);
TASK_PP(16'h1C410,4);
TASK_PP(16'h1C411,4);
TASK_PP(16'h1C412,4);
TASK_PP(16'h1C413,4);
TASK_PP(16'h1C414,4);
TASK_PP(16'h1C415,4);
TASK_PP(16'h1C416,4);
TASK_PP(16'h1C417,4);
TASK_PP(16'h1C418,4);
TASK_PP(16'h1C419,4);
TASK_PP(16'h1C41A,4);
TASK_PP(16'h1C41B,4);
TASK_PP(16'h1C41C,4);
TASK_PP(16'h1C41D,4);
TASK_PP(16'h1C41E,4);
TASK_PP(16'h1C41F,4);
TASK_PP(16'h1C420,4);
TASK_PP(16'h1C421,4);
TASK_PP(16'h1C422,4);
TASK_PP(16'h1C423,4);
TASK_PP(16'h1C424,4);
TASK_PP(16'h1C425,4);
TASK_PP(16'h1C426,4);
TASK_PP(16'h1C427,4);
TASK_PP(16'h1C428,4);
TASK_PP(16'h1C429,4);
TASK_PP(16'h1C42A,4);
TASK_PP(16'h1C42B,4);
TASK_PP(16'h1C42C,4);
TASK_PP(16'h1C42D,4);
TASK_PP(16'h1C42E,4);
TASK_PP(16'h1C42F,4);
TASK_PP(16'h1C430,4);
TASK_PP(16'h1C431,4);
TASK_PP(16'h1C432,4);
TASK_PP(16'h1C433,4);
TASK_PP(16'h1C434,4);
TASK_PP(16'h1C435,4);
TASK_PP(16'h1C436,4);
TASK_PP(16'h1C437,4);
TASK_PP(16'h1C438,4);
TASK_PP(16'h1C439,4);
TASK_PP(16'h1C43A,4);
TASK_PP(16'h1C43B,4);
TASK_PP(16'h1C43C,4);
TASK_PP(16'h1C43D,4);
TASK_PP(16'h1C43E,4);
TASK_PP(16'h1C43F,4);
TASK_PP(16'h1C440,4);
TASK_PP(16'h1C441,4);
TASK_PP(16'h1C442,4);
TASK_PP(16'h1C443,4);
TASK_PP(16'h1C444,4);
TASK_PP(16'h1C445,4);
TASK_PP(16'h1C446,4);
TASK_PP(16'h1C447,4);
TASK_PP(16'h1C448,4);
TASK_PP(16'h1C449,4);
TASK_PP(16'h1C44A,4);
TASK_PP(16'h1C44B,4);
TASK_PP(16'h1C44C,4);
TASK_PP(16'h1C44D,4);
TASK_PP(16'h1C44E,4);
TASK_PP(16'h1C44F,4);
TASK_PP(16'h1C450,4);
TASK_PP(16'h1C451,4);
TASK_PP(16'h1C452,4);
TASK_PP(16'h1C453,4);
TASK_PP(16'h1C454,4);
TASK_PP(16'h1C455,4);
TASK_PP(16'h1C456,4);
TASK_PP(16'h1C457,4);
TASK_PP(16'h1C458,4);
TASK_PP(16'h1C459,4);
TASK_PP(16'h1C45A,4);
TASK_PP(16'h1C45B,4);
TASK_PP(16'h1C45C,4);
TASK_PP(16'h1C45D,4);
TASK_PP(16'h1C45E,4);
TASK_PP(16'h1C45F,4);
TASK_PP(16'h1C460,4);
TASK_PP(16'h1C461,4);
TASK_PP(16'h1C462,4);
TASK_PP(16'h1C463,4);
TASK_PP(16'h1C464,4);
TASK_PP(16'h1C465,4);
TASK_PP(16'h1C466,4);
TASK_PP(16'h1C467,4);
TASK_PP(16'h1C468,4);
TASK_PP(16'h1C469,4);
TASK_PP(16'h1C46A,4);
TASK_PP(16'h1C46B,4);
TASK_PP(16'h1C46C,4);
TASK_PP(16'h1C46D,4);
TASK_PP(16'h1C46E,4);
TASK_PP(16'h1C46F,4);
TASK_PP(16'h1C470,4);
TASK_PP(16'h1C471,4);
TASK_PP(16'h1C472,4);
TASK_PP(16'h1C473,4);
TASK_PP(16'h1C474,4);
TASK_PP(16'h1C475,4);
TASK_PP(16'h1C476,4);
TASK_PP(16'h1C477,4);
TASK_PP(16'h1C478,4);
TASK_PP(16'h1C479,4);
TASK_PP(16'h1C47A,4);
TASK_PP(16'h1C47B,4);
TASK_PP(16'h1C47C,4);
TASK_PP(16'h1C47D,4);
TASK_PP(16'h1C47E,4);
TASK_PP(16'h1C47F,4);
TASK_PP(16'h1C480,4);
TASK_PP(16'h1C481,4);
TASK_PP(16'h1C482,4);
TASK_PP(16'h1C483,4);
TASK_PP(16'h1C484,4);
TASK_PP(16'h1C485,4);
TASK_PP(16'h1C486,4);
TASK_PP(16'h1C487,4);
TASK_PP(16'h1C488,4);
TASK_PP(16'h1C489,4);
TASK_PP(16'h1C48A,4);
TASK_PP(16'h1C48B,4);
TASK_PP(16'h1C48C,4);
TASK_PP(16'h1C48D,4);
TASK_PP(16'h1C48E,4);
TASK_PP(16'h1C48F,4);
TASK_PP(16'h1C490,4);
TASK_PP(16'h1C491,4);
TASK_PP(16'h1C492,4);
TASK_PP(16'h1C493,4);
TASK_PP(16'h1C494,4);
TASK_PP(16'h1C495,4);
TASK_PP(16'h1C496,4);
TASK_PP(16'h1C497,4);
TASK_PP(16'h1C498,4);
TASK_PP(16'h1C499,4);
TASK_PP(16'h1C49A,4);
TASK_PP(16'h1C49B,4);
TASK_PP(16'h1C49C,4);
TASK_PP(16'h1C49D,4);
TASK_PP(16'h1C49E,4);
TASK_PP(16'h1C49F,4);
TASK_PP(16'h1C4A0,4);
TASK_PP(16'h1C4A1,4);
TASK_PP(16'h1C4A2,4);
TASK_PP(16'h1C4A3,4);
TASK_PP(16'h1C4A4,4);
TASK_PP(16'h1C4A5,4);
TASK_PP(16'h1C4A6,4);
TASK_PP(16'h1C4A7,4);
TASK_PP(16'h1C4A8,4);
TASK_PP(16'h1C4A9,4);
TASK_PP(16'h1C4AA,4);
TASK_PP(16'h1C4AB,4);
TASK_PP(16'h1C4AC,4);
TASK_PP(16'h1C4AD,4);
TASK_PP(16'h1C4AE,4);
TASK_PP(16'h1C4AF,4);
TASK_PP(16'h1C4B0,4);
TASK_PP(16'h1C4B1,4);
TASK_PP(16'h1C4B2,4);
TASK_PP(16'h1C4B3,4);
TASK_PP(16'h1C4B4,4);
TASK_PP(16'h1C4B5,4);
TASK_PP(16'h1C4B6,4);
TASK_PP(16'h1C4B7,4);
TASK_PP(16'h1C4B8,4);
TASK_PP(16'h1C4B9,4);
TASK_PP(16'h1C4BA,4);
TASK_PP(16'h1C4BB,4);
TASK_PP(16'h1C4BC,4);
TASK_PP(16'h1C4BD,4);
TASK_PP(16'h1C4BE,4);
TASK_PP(16'h1C4BF,4);
TASK_PP(16'h1C4C0,4);
TASK_PP(16'h1C4C1,4);
TASK_PP(16'h1C4C2,4);
TASK_PP(16'h1C4C3,4);
TASK_PP(16'h1C4C4,4);
TASK_PP(16'h1C4C5,4);
TASK_PP(16'h1C4C6,4);
TASK_PP(16'h1C4C7,4);
TASK_PP(16'h1C4C8,4);
TASK_PP(16'h1C4C9,4);
TASK_PP(16'h1C4CA,4);
TASK_PP(16'h1C4CB,4);
TASK_PP(16'h1C4CC,4);
TASK_PP(16'h1C4CD,4);
TASK_PP(16'h1C4CE,4);
TASK_PP(16'h1C4CF,4);
TASK_PP(16'h1C4D0,4);
TASK_PP(16'h1C4D1,4);
TASK_PP(16'h1C4D2,4);
TASK_PP(16'h1C4D3,4);
TASK_PP(16'h1C4D4,4);
TASK_PP(16'h1C4D5,4);
TASK_PP(16'h1C4D6,4);
TASK_PP(16'h1C4D7,4);
TASK_PP(16'h1C4D8,4);
TASK_PP(16'h1C4D9,4);
TASK_PP(16'h1C4DA,4);
TASK_PP(16'h1C4DB,4);
TASK_PP(16'h1C4DC,4);
TASK_PP(16'h1C4DD,4);
TASK_PP(16'h1C4DE,4);
TASK_PP(16'h1C4DF,4);
TASK_PP(16'h1C4E0,4);
TASK_PP(16'h1C4E1,4);
TASK_PP(16'h1C4E2,4);
TASK_PP(16'h1C4E3,4);
TASK_PP(16'h1C4E4,4);
TASK_PP(16'h1C4E5,4);
TASK_PP(16'h1C4E6,4);
TASK_PP(16'h1C4E7,4);
TASK_PP(16'h1C4E8,4);
TASK_PP(16'h1C4E9,4);
TASK_PP(16'h1C4EA,4);
TASK_PP(16'h1C4EB,4);
TASK_PP(16'h1C4EC,4);
TASK_PP(16'h1C4ED,4);
TASK_PP(16'h1C4EE,4);
TASK_PP(16'h1C4EF,4);
TASK_PP(16'h1C4F0,4);
TASK_PP(16'h1C4F1,4);
TASK_PP(16'h1C4F2,4);
TASK_PP(16'h1C4F3,4);
TASK_PP(16'h1C4F4,4);
TASK_PP(16'h1C4F5,4);
TASK_PP(16'h1C4F6,4);
TASK_PP(16'h1C4F7,4);
TASK_PP(16'h1C4F8,4);
TASK_PP(16'h1C4F9,4);
TASK_PP(16'h1C4FA,4);
TASK_PP(16'h1C4FB,4);
TASK_PP(16'h1C4FC,4);
TASK_PP(16'h1C4FD,4);
TASK_PP(16'h1C4FE,4);
TASK_PP(16'h1C4FF,4);
TASK_PP(16'h1C500,4);
TASK_PP(16'h1C501,4);
TASK_PP(16'h1C502,4);
TASK_PP(16'h1C503,4);
TASK_PP(16'h1C504,4);
TASK_PP(16'h1C505,4);
TASK_PP(16'h1C506,4);
TASK_PP(16'h1C507,4);
TASK_PP(16'h1C508,4);
TASK_PP(16'h1C509,4);
TASK_PP(16'h1C50A,4);
TASK_PP(16'h1C50B,4);
TASK_PP(16'h1C50C,4);
TASK_PP(16'h1C50D,4);
TASK_PP(16'h1C50E,4);
TASK_PP(16'h1C50F,4);
TASK_PP(16'h1C510,4);
TASK_PP(16'h1C511,4);
TASK_PP(16'h1C512,4);
TASK_PP(16'h1C513,4);
TASK_PP(16'h1C514,4);
TASK_PP(16'h1C515,4);
TASK_PP(16'h1C516,4);
TASK_PP(16'h1C517,4);
TASK_PP(16'h1C518,4);
TASK_PP(16'h1C519,4);
TASK_PP(16'h1C51A,4);
TASK_PP(16'h1C51B,4);
TASK_PP(16'h1C51C,4);
TASK_PP(16'h1C51D,4);
TASK_PP(16'h1C51E,4);
TASK_PP(16'h1C51F,4);
TASK_PP(16'h1C520,4);
TASK_PP(16'h1C521,4);
TASK_PP(16'h1C522,4);
TASK_PP(16'h1C523,4);
TASK_PP(16'h1C524,4);
TASK_PP(16'h1C525,4);
TASK_PP(16'h1C526,4);
TASK_PP(16'h1C527,4);
TASK_PP(16'h1C528,4);
TASK_PP(16'h1C529,4);
TASK_PP(16'h1C52A,4);
TASK_PP(16'h1C52B,4);
TASK_PP(16'h1C52C,4);
TASK_PP(16'h1C52D,4);
TASK_PP(16'h1C52E,4);
TASK_PP(16'h1C52F,4);
TASK_PP(16'h1C530,4);
TASK_PP(16'h1C531,4);
TASK_PP(16'h1C532,4);
TASK_PP(16'h1C533,4);
TASK_PP(16'h1C534,4);
TASK_PP(16'h1C535,4);
TASK_PP(16'h1C536,4);
TASK_PP(16'h1C537,4);
TASK_PP(16'h1C538,4);
TASK_PP(16'h1C539,4);
TASK_PP(16'h1C53A,4);
TASK_PP(16'h1C53B,4);
TASK_PP(16'h1C53C,4);
TASK_PP(16'h1C53D,4);
TASK_PP(16'h1C53E,4);
TASK_PP(16'h1C53F,4);
TASK_PP(16'h1C540,4);
TASK_PP(16'h1C541,4);
TASK_PP(16'h1C542,4);
TASK_PP(16'h1C543,4);
TASK_PP(16'h1C544,4);
TASK_PP(16'h1C545,4);
TASK_PP(16'h1C546,4);
TASK_PP(16'h1C547,4);
TASK_PP(16'h1C548,4);
TASK_PP(16'h1C549,4);
TASK_PP(16'h1C54A,4);
TASK_PP(16'h1C54B,4);
TASK_PP(16'h1C54C,4);
TASK_PP(16'h1C54D,4);
TASK_PP(16'h1C54E,4);
TASK_PP(16'h1C54F,4);
TASK_PP(16'h1C550,4);
TASK_PP(16'h1C551,4);
TASK_PP(16'h1C552,4);
TASK_PP(16'h1C553,4);
TASK_PP(16'h1C554,4);
TASK_PP(16'h1C555,4);
TASK_PP(16'h1C556,4);
TASK_PP(16'h1C557,4);
TASK_PP(16'h1C558,4);
TASK_PP(16'h1C559,4);
TASK_PP(16'h1C55A,4);
TASK_PP(16'h1C55B,4);
TASK_PP(16'h1C55C,4);
TASK_PP(16'h1C55D,4);
TASK_PP(16'h1C55E,4);
TASK_PP(16'h1C55F,4);
TASK_PP(16'h1C560,4);
TASK_PP(16'h1C561,4);
TASK_PP(16'h1C562,4);
TASK_PP(16'h1C563,4);
TASK_PP(16'h1C564,4);
TASK_PP(16'h1C565,4);
TASK_PP(16'h1C566,4);
TASK_PP(16'h1C567,4);
TASK_PP(16'h1C568,4);
TASK_PP(16'h1C569,4);
TASK_PP(16'h1C56A,4);
TASK_PP(16'h1C56B,4);
TASK_PP(16'h1C56C,4);
TASK_PP(16'h1C56D,4);
TASK_PP(16'h1C56E,4);
TASK_PP(16'h1C56F,4);
TASK_PP(16'h1C570,4);
TASK_PP(16'h1C571,4);
TASK_PP(16'h1C572,4);
TASK_PP(16'h1C573,4);
TASK_PP(16'h1C574,4);
TASK_PP(16'h1C575,4);
TASK_PP(16'h1C576,4);
TASK_PP(16'h1C577,4);
TASK_PP(16'h1C578,4);
TASK_PP(16'h1C579,4);
TASK_PP(16'h1C57A,4);
TASK_PP(16'h1C57B,4);
TASK_PP(16'h1C57C,4);
TASK_PP(16'h1C57D,4);
TASK_PP(16'h1C57E,4);
TASK_PP(16'h1C57F,4);
TASK_PP(16'h1C580,4);
TASK_PP(16'h1C581,4);
TASK_PP(16'h1C582,4);
TASK_PP(16'h1C583,4);
TASK_PP(16'h1C584,4);
TASK_PP(16'h1C585,4);
TASK_PP(16'h1C586,4);
TASK_PP(16'h1C587,4);
TASK_PP(16'h1C588,4);
TASK_PP(16'h1C589,4);
TASK_PP(16'h1C58A,4);
TASK_PP(16'h1C58B,4);
TASK_PP(16'h1C58C,4);
TASK_PP(16'h1C58D,4);
TASK_PP(16'h1C58E,4);
TASK_PP(16'h1C58F,4);
TASK_PP(16'h1C590,4);
TASK_PP(16'h1C591,4);
TASK_PP(16'h1C592,4);
TASK_PP(16'h1C593,4);
TASK_PP(16'h1C594,4);
TASK_PP(16'h1C595,4);
TASK_PP(16'h1C596,4);
TASK_PP(16'h1C597,4);
TASK_PP(16'h1C598,4);
TASK_PP(16'h1C599,4);
TASK_PP(16'h1C59A,4);
TASK_PP(16'h1C59B,4);
TASK_PP(16'h1C59C,4);
TASK_PP(16'h1C59D,4);
TASK_PP(16'h1C59E,4);
TASK_PP(16'h1C59F,4);
TASK_PP(16'h1C5A0,4);
TASK_PP(16'h1C5A1,4);
TASK_PP(16'h1C5A2,4);
TASK_PP(16'h1C5A3,4);
TASK_PP(16'h1C5A4,4);
TASK_PP(16'h1C5A5,4);
TASK_PP(16'h1C5A6,4);
TASK_PP(16'h1C5A7,4);
TASK_PP(16'h1C5A8,4);
TASK_PP(16'h1C5A9,4);
TASK_PP(16'h1C5AA,4);
TASK_PP(16'h1C5AB,4);
TASK_PP(16'h1C5AC,4);
TASK_PP(16'h1C5AD,4);
TASK_PP(16'h1C5AE,4);
TASK_PP(16'h1C5AF,4);
TASK_PP(16'h1C5B0,4);
TASK_PP(16'h1C5B1,4);
TASK_PP(16'h1C5B2,4);
TASK_PP(16'h1C5B3,4);
TASK_PP(16'h1C5B4,4);
TASK_PP(16'h1C5B5,4);
TASK_PP(16'h1C5B6,4);
TASK_PP(16'h1C5B7,4);
TASK_PP(16'h1C5B8,4);
TASK_PP(16'h1C5B9,4);
TASK_PP(16'h1C5BA,4);
TASK_PP(16'h1C5BB,4);
TASK_PP(16'h1C5BC,4);
TASK_PP(16'h1C5BD,4);
TASK_PP(16'h1C5BE,4);
TASK_PP(16'h1C5BF,4);
TASK_PP(16'h1C5C0,4);
TASK_PP(16'h1C5C1,4);
TASK_PP(16'h1C5C2,4);
TASK_PP(16'h1C5C3,4);
TASK_PP(16'h1C5C4,4);
TASK_PP(16'h1C5C5,4);
TASK_PP(16'h1C5C6,4);
TASK_PP(16'h1C5C7,4);
TASK_PP(16'h1C5C8,4);
TASK_PP(16'h1C5C9,4);
TASK_PP(16'h1C5CA,4);
TASK_PP(16'h1C5CB,4);
TASK_PP(16'h1C5CC,4);
TASK_PP(16'h1C5CD,4);
TASK_PP(16'h1C5CE,4);
TASK_PP(16'h1C5CF,4);
TASK_PP(16'h1C5D0,4);
TASK_PP(16'h1C5D1,4);
TASK_PP(16'h1C5D2,4);
TASK_PP(16'h1C5D3,4);
TASK_PP(16'h1C5D4,4);
TASK_PP(16'h1C5D5,4);
TASK_PP(16'h1C5D6,4);
TASK_PP(16'h1C5D7,4);
TASK_PP(16'h1C5D8,4);
TASK_PP(16'h1C5D9,4);
TASK_PP(16'h1C5DA,4);
TASK_PP(16'h1C5DB,4);
TASK_PP(16'h1C5DC,4);
TASK_PP(16'h1C5DD,4);
TASK_PP(16'h1C5DE,4);
TASK_PP(16'h1C5DF,4);
TASK_PP(16'h1C5E0,4);
TASK_PP(16'h1C5E1,4);
TASK_PP(16'h1C5E2,4);
TASK_PP(16'h1C5E3,4);
TASK_PP(16'h1C5E4,4);
TASK_PP(16'h1C5E5,4);
TASK_PP(16'h1C5E6,4);
TASK_PP(16'h1C5E7,4);
TASK_PP(16'h1C5E8,4);
TASK_PP(16'h1C5E9,4);
TASK_PP(16'h1C5EA,4);
TASK_PP(16'h1C5EB,4);
TASK_PP(16'h1C5EC,4);
TASK_PP(16'h1C5ED,4);
TASK_PP(16'h1C5EE,4);
TASK_PP(16'h1C5EF,4);
TASK_PP(16'h1C5F0,4);
TASK_PP(16'h1C5F1,4);
TASK_PP(16'h1C5F2,4);
TASK_PP(16'h1C5F3,4);
TASK_PP(16'h1C5F4,4);
TASK_PP(16'h1C5F5,4);
TASK_PP(16'h1C5F6,4);
TASK_PP(16'h1C5F7,4);
TASK_PP(16'h1C5F8,4);
TASK_PP(16'h1C5F9,4);
TASK_PP(16'h1C5FA,4);
TASK_PP(16'h1C5FB,4);
TASK_PP(16'h1C5FC,4);
TASK_PP(16'h1C5FD,4);
TASK_PP(16'h1C5FE,4);
TASK_PP(16'h1C5FF,4);
TASK_PP(16'h1C600,4);
TASK_PP(16'h1C601,4);
TASK_PP(16'h1C602,4);
TASK_PP(16'h1C603,4);
TASK_PP(16'h1C604,4);
TASK_PP(16'h1C605,4);
TASK_PP(16'h1C606,4);
TASK_PP(16'h1C607,4);
TASK_PP(16'h1C608,4);
TASK_PP(16'h1C609,4);
TASK_PP(16'h1C60A,4);
TASK_PP(16'h1C60B,4);
TASK_PP(16'h1C60C,4);
TASK_PP(16'h1C60D,4);
TASK_PP(16'h1C60E,4);
TASK_PP(16'h1C60F,4);
TASK_PP(16'h1C610,4);
TASK_PP(16'h1C611,4);
TASK_PP(16'h1C612,4);
TASK_PP(16'h1C613,4);
TASK_PP(16'h1C614,4);
TASK_PP(16'h1C615,4);
TASK_PP(16'h1C616,4);
TASK_PP(16'h1C617,4);
TASK_PP(16'h1C618,4);
TASK_PP(16'h1C619,4);
TASK_PP(16'h1C61A,4);
TASK_PP(16'h1C61B,4);
TASK_PP(16'h1C61C,4);
TASK_PP(16'h1C61D,4);
TASK_PP(16'h1C61E,4);
TASK_PP(16'h1C61F,4);
TASK_PP(16'h1C620,4);
TASK_PP(16'h1C621,4);
TASK_PP(16'h1C622,4);
TASK_PP(16'h1C623,4);
TASK_PP(16'h1C624,4);
TASK_PP(16'h1C625,4);
TASK_PP(16'h1C626,4);
TASK_PP(16'h1C627,4);
TASK_PP(16'h1C628,4);
TASK_PP(16'h1C629,4);
TASK_PP(16'h1C62A,4);
TASK_PP(16'h1C62B,4);
TASK_PP(16'h1C62C,4);
TASK_PP(16'h1C62D,4);
TASK_PP(16'h1C62E,4);
TASK_PP(16'h1C62F,4);
TASK_PP(16'h1C630,4);
TASK_PP(16'h1C631,4);
TASK_PP(16'h1C632,4);
TASK_PP(16'h1C633,4);
TASK_PP(16'h1C634,4);
TASK_PP(16'h1C635,4);
TASK_PP(16'h1C636,4);
TASK_PP(16'h1C637,4);
TASK_PP(16'h1C638,4);
TASK_PP(16'h1C639,4);
TASK_PP(16'h1C63A,4);
TASK_PP(16'h1C63B,4);
TASK_PP(16'h1C63C,4);
TASK_PP(16'h1C63D,4);
TASK_PP(16'h1C63E,4);
TASK_PP(16'h1C63F,4);
TASK_PP(16'h1C640,4);
TASK_PP(16'h1C641,4);
TASK_PP(16'h1C642,4);
TASK_PP(16'h1C643,4);
TASK_PP(16'h1C644,4);
TASK_PP(16'h1C645,4);
TASK_PP(16'h1C646,4);
TASK_PP(16'h1C647,4);
TASK_PP(16'h1C648,4);
TASK_PP(16'h1C649,4);
TASK_PP(16'h1C64A,4);
TASK_PP(16'h1C64B,4);
TASK_PP(16'h1C64C,4);
TASK_PP(16'h1C64D,4);
TASK_PP(16'h1C64E,4);
TASK_PP(16'h1C64F,4);
TASK_PP(16'h1C650,4);
TASK_PP(16'h1C651,4);
TASK_PP(16'h1C652,4);
TASK_PP(16'h1C653,4);
TASK_PP(16'h1C654,4);
TASK_PP(16'h1C655,4);
TASK_PP(16'h1C656,4);
TASK_PP(16'h1C657,4);
TASK_PP(16'h1C658,4);
TASK_PP(16'h1C659,4);
TASK_PP(16'h1C65A,4);
TASK_PP(16'h1C65B,4);
TASK_PP(16'h1C65C,4);
TASK_PP(16'h1C65D,4);
TASK_PP(16'h1C65E,4);
TASK_PP(16'h1C65F,4);
TASK_PP(16'h1C660,4);
TASK_PP(16'h1C661,4);
TASK_PP(16'h1C662,4);
TASK_PP(16'h1C663,4);
TASK_PP(16'h1C664,4);
TASK_PP(16'h1C665,4);
TASK_PP(16'h1C666,4);
TASK_PP(16'h1C667,4);
TASK_PP(16'h1C668,4);
TASK_PP(16'h1C669,4);
TASK_PP(16'h1C66A,4);
TASK_PP(16'h1C66B,4);
TASK_PP(16'h1C66C,4);
TASK_PP(16'h1C66D,4);
TASK_PP(16'h1C66E,4);
TASK_PP(16'h1C66F,4);
TASK_PP(16'h1C670,4);
TASK_PP(16'h1C671,4);
TASK_PP(16'h1C672,4);
TASK_PP(16'h1C673,4);
TASK_PP(16'h1C674,4);
TASK_PP(16'h1C675,4);
TASK_PP(16'h1C676,4);
TASK_PP(16'h1C677,4);
TASK_PP(16'h1C678,4);
TASK_PP(16'h1C679,4);
TASK_PP(16'h1C67A,4);
TASK_PP(16'h1C67B,4);
TASK_PP(16'h1C67C,4);
TASK_PP(16'h1C67D,4);
TASK_PP(16'h1C67E,4);
TASK_PP(16'h1C67F,4);
TASK_PP(16'h1C680,4);
TASK_PP(16'h1C681,4);
TASK_PP(16'h1C682,4);
TASK_PP(16'h1C683,4);
TASK_PP(16'h1C684,4);
TASK_PP(16'h1C685,4);
TASK_PP(16'h1C686,4);
TASK_PP(16'h1C687,4);
TASK_PP(16'h1C688,4);
TASK_PP(16'h1C689,4);
TASK_PP(16'h1C68A,4);
TASK_PP(16'h1C68B,4);
TASK_PP(16'h1C68C,4);
TASK_PP(16'h1C68D,4);
TASK_PP(16'h1C68E,4);
TASK_PP(16'h1C68F,4);
TASK_PP(16'h1C690,4);
TASK_PP(16'h1C691,4);
TASK_PP(16'h1C692,4);
TASK_PP(16'h1C693,4);
TASK_PP(16'h1C694,4);
TASK_PP(16'h1C695,4);
TASK_PP(16'h1C696,4);
TASK_PP(16'h1C697,4);
TASK_PP(16'h1C698,4);
TASK_PP(16'h1C699,4);
TASK_PP(16'h1C69A,4);
TASK_PP(16'h1C69B,4);
TASK_PP(16'h1C69C,4);
TASK_PP(16'h1C69D,4);
TASK_PP(16'h1C69E,4);
TASK_PP(16'h1C69F,4);
TASK_PP(16'h1C6A0,4);
TASK_PP(16'h1C6A1,4);
TASK_PP(16'h1C6A2,4);
TASK_PP(16'h1C6A3,4);
TASK_PP(16'h1C6A4,4);
TASK_PP(16'h1C6A5,4);
TASK_PP(16'h1C6A6,4);
TASK_PP(16'h1C6A7,4);
TASK_PP(16'h1C6A8,4);
TASK_PP(16'h1C6A9,4);
TASK_PP(16'h1C6AA,4);
TASK_PP(16'h1C6AB,4);
TASK_PP(16'h1C6AC,4);
TASK_PP(16'h1C6AD,4);
TASK_PP(16'h1C6AE,4);
TASK_PP(16'h1C6AF,4);
TASK_PP(16'h1C6B0,4);
TASK_PP(16'h1C6B1,4);
TASK_PP(16'h1C6B2,4);
TASK_PP(16'h1C6B3,4);
TASK_PP(16'h1C6B4,4);
TASK_PP(16'h1C6B5,4);
TASK_PP(16'h1C6B6,4);
TASK_PP(16'h1C6B7,4);
TASK_PP(16'h1C6B8,4);
TASK_PP(16'h1C6B9,4);
TASK_PP(16'h1C6BA,4);
TASK_PP(16'h1C6BB,4);
TASK_PP(16'h1C6BC,4);
TASK_PP(16'h1C6BD,4);
TASK_PP(16'h1C6BE,4);
TASK_PP(16'h1C6BF,4);
TASK_PP(16'h1C6C0,4);
TASK_PP(16'h1C6C1,4);
TASK_PP(16'h1C6C2,4);
TASK_PP(16'h1C6C3,4);
TASK_PP(16'h1C6C4,4);
TASK_PP(16'h1C6C5,4);
TASK_PP(16'h1C6C6,4);
TASK_PP(16'h1C6C7,4);
TASK_PP(16'h1C6C8,4);
TASK_PP(16'h1C6C9,4);
TASK_PP(16'h1C6CA,4);
TASK_PP(16'h1C6CB,4);
TASK_PP(16'h1C6CC,4);
TASK_PP(16'h1C6CD,4);
TASK_PP(16'h1C6CE,4);
TASK_PP(16'h1C6CF,4);
TASK_PP(16'h1C6D0,4);
TASK_PP(16'h1C6D1,4);
TASK_PP(16'h1C6D2,4);
TASK_PP(16'h1C6D3,4);
TASK_PP(16'h1C6D4,4);
TASK_PP(16'h1C6D5,4);
TASK_PP(16'h1C6D6,4);
TASK_PP(16'h1C6D7,4);
TASK_PP(16'h1C6D8,4);
TASK_PP(16'h1C6D9,4);
TASK_PP(16'h1C6DA,4);
TASK_PP(16'h1C6DB,4);
TASK_PP(16'h1C6DC,4);
TASK_PP(16'h1C6DD,4);
TASK_PP(16'h1C6DE,4);
TASK_PP(16'h1C6DF,4);
TASK_PP(16'h1C6E0,4);
TASK_PP(16'h1C6E1,4);
TASK_PP(16'h1C6E2,4);
TASK_PP(16'h1C6E3,4);
TASK_PP(16'h1C6E4,4);
TASK_PP(16'h1C6E5,4);
TASK_PP(16'h1C6E6,4);
TASK_PP(16'h1C6E7,4);
TASK_PP(16'h1C6E8,4);
TASK_PP(16'h1C6E9,4);
TASK_PP(16'h1C6EA,4);
TASK_PP(16'h1C6EB,4);
TASK_PP(16'h1C6EC,4);
TASK_PP(16'h1C6ED,4);
TASK_PP(16'h1C6EE,4);
TASK_PP(16'h1C6EF,4);
TASK_PP(16'h1C6F0,4);
TASK_PP(16'h1C6F1,4);
TASK_PP(16'h1C6F2,4);
TASK_PP(16'h1C6F3,4);
TASK_PP(16'h1C6F4,4);
TASK_PP(16'h1C6F5,4);
TASK_PP(16'h1C6F6,4);
TASK_PP(16'h1C6F7,4);
TASK_PP(16'h1C6F8,4);
TASK_PP(16'h1C6F9,4);
TASK_PP(16'h1C6FA,4);
TASK_PP(16'h1C6FB,4);
TASK_PP(16'h1C6FC,4);
TASK_PP(16'h1C6FD,4);
TASK_PP(16'h1C6FE,4);
TASK_PP(16'h1C6FF,4);
TASK_PP(16'h1C700,4);
TASK_PP(16'h1C701,4);
TASK_PP(16'h1C702,4);
TASK_PP(16'h1C703,4);
TASK_PP(16'h1C704,4);
TASK_PP(16'h1C705,4);
TASK_PP(16'h1C706,4);
TASK_PP(16'h1C707,4);
TASK_PP(16'h1C708,4);
TASK_PP(16'h1C709,4);
TASK_PP(16'h1C70A,4);
TASK_PP(16'h1C70B,4);
TASK_PP(16'h1C70C,4);
TASK_PP(16'h1C70D,4);
TASK_PP(16'h1C70E,4);
TASK_PP(16'h1C70F,4);
TASK_PP(16'h1C710,4);
TASK_PP(16'h1C711,4);
TASK_PP(16'h1C712,4);
TASK_PP(16'h1C713,4);
TASK_PP(16'h1C714,4);
TASK_PP(16'h1C715,4);
TASK_PP(16'h1C716,4);
TASK_PP(16'h1C717,4);
TASK_PP(16'h1C718,4);
TASK_PP(16'h1C719,4);
TASK_PP(16'h1C71A,4);
TASK_PP(16'h1C71B,4);
TASK_PP(16'h1C71C,4);
TASK_PP(16'h1C71D,4);
TASK_PP(16'h1C71E,4);
TASK_PP(16'h1C71F,4);
TASK_PP(16'h1C720,4);
TASK_PP(16'h1C721,4);
TASK_PP(16'h1C722,4);
TASK_PP(16'h1C723,4);
TASK_PP(16'h1C724,4);
TASK_PP(16'h1C725,4);
TASK_PP(16'h1C726,4);
TASK_PP(16'h1C727,4);
TASK_PP(16'h1C728,4);
TASK_PP(16'h1C729,4);
TASK_PP(16'h1C72A,4);
TASK_PP(16'h1C72B,4);
TASK_PP(16'h1C72C,4);
TASK_PP(16'h1C72D,4);
TASK_PP(16'h1C72E,4);
TASK_PP(16'h1C72F,4);
TASK_PP(16'h1C730,4);
TASK_PP(16'h1C731,4);
TASK_PP(16'h1C732,4);
TASK_PP(16'h1C733,4);
TASK_PP(16'h1C734,4);
TASK_PP(16'h1C735,4);
TASK_PP(16'h1C736,4);
TASK_PP(16'h1C737,4);
TASK_PP(16'h1C738,4);
TASK_PP(16'h1C739,4);
TASK_PP(16'h1C73A,4);
TASK_PP(16'h1C73B,4);
TASK_PP(16'h1C73C,4);
TASK_PP(16'h1C73D,4);
TASK_PP(16'h1C73E,4);
TASK_PP(16'h1C73F,4);
TASK_PP(16'h1C740,4);
TASK_PP(16'h1C741,4);
TASK_PP(16'h1C742,4);
TASK_PP(16'h1C743,4);
TASK_PP(16'h1C744,4);
TASK_PP(16'h1C745,4);
TASK_PP(16'h1C746,4);
TASK_PP(16'h1C747,4);
TASK_PP(16'h1C748,4);
TASK_PP(16'h1C749,4);
TASK_PP(16'h1C74A,4);
TASK_PP(16'h1C74B,4);
TASK_PP(16'h1C74C,4);
TASK_PP(16'h1C74D,4);
TASK_PP(16'h1C74E,4);
TASK_PP(16'h1C74F,4);
TASK_PP(16'h1C750,4);
TASK_PP(16'h1C751,4);
TASK_PP(16'h1C752,4);
TASK_PP(16'h1C753,4);
TASK_PP(16'h1C754,4);
TASK_PP(16'h1C755,4);
TASK_PP(16'h1C756,4);
TASK_PP(16'h1C757,4);
TASK_PP(16'h1C758,4);
TASK_PP(16'h1C759,4);
TASK_PP(16'h1C75A,4);
TASK_PP(16'h1C75B,4);
TASK_PP(16'h1C75C,4);
TASK_PP(16'h1C75D,4);
TASK_PP(16'h1C75E,4);
TASK_PP(16'h1C75F,4);
TASK_PP(16'h1C760,4);
TASK_PP(16'h1C761,4);
TASK_PP(16'h1C762,4);
TASK_PP(16'h1C763,4);
TASK_PP(16'h1C764,4);
TASK_PP(16'h1C765,4);
TASK_PP(16'h1C766,4);
TASK_PP(16'h1C767,4);
TASK_PP(16'h1C768,4);
TASK_PP(16'h1C769,4);
TASK_PP(16'h1C76A,4);
TASK_PP(16'h1C76B,4);
TASK_PP(16'h1C76C,4);
TASK_PP(16'h1C76D,4);
TASK_PP(16'h1C76E,4);
TASK_PP(16'h1C76F,4);
TASK_PP(16'h1C770,4);
TASK_PP(16'h1C771,4);
TASK_PP(16'h1C772,4);
TASK_PP(16'h1C773,4);
TASK_PP(16'h1C774,4);
TASK_PP(16'h1C775,4);
TASK_PP(16'h1C776,4);
TASK_PP(16'h1C777,4);
TASK_PP(16'h1C778,4);
TASK_PP(16'h1C779,4);
TASK_PP(16'h1C77A,4);
TASK_PP(16'h1C77B,4);
TASK_PP(16'h1C77C,4);
TASK_PP(16'h1C77D,4);
TASK_PP(16'h1C77E,4);
TASK_PP(16'h1C77F,4);
TASK_PP(16'h1C780,4);
TASK_PP(16'h1C781,4);
TASK_PP(16'h1C782,4);
TASK_PP(16'h1C783,4);
TASK_PP(16'h1C784,4);
TASK_PP(16'h1C785,4);
TASK_PP(16'h1C786,4);
TASK_PP(16'h1C787,4);
TASK_PP(16'h1C788,4);
TASK_PP(16'h1C789,4);
TASK_PP(16'h1C78A,4);
TASK_PP(16'h1C78B,4);
TASK_PP(16'h1C78C,4);
TASK_PP(16'h1C78D,4);
TASK_PP(16'h1C78E,4);
TASK_PP(16'h1C78F,4);
TASK_PP(16'h1C790,4);
TASK_PP(16'h1C791,4);
TASK_PP(16'h1C792,4);
TASK_PP(16'h1C793,4);
TASK_PP(16'h1C794,4);
TASK_PP(16'h1C795,4);
TASK_PP(16'h1C796,4);
TASK_PP(16'h1C797,4);
TASK_PP(16'h1C798,4);
TASK_PP(16'h1C799,4);
TASK_PP(16'h1C79A,4);
TASK_PP(16'h1C79B,4);
TASK_PP(16'h1C79C,4);
TASK_PP(16'h1C79D,4);
TASK_PP(16'h1C79E,4);
TASK_PP(16'h1C79F,4);
TASK_PP(16'h1C7A0,4);
TASK_PP(16'h1C7A1,4);
TASK_PP(16'h1C7A2,4);
TASK_PP(16'h1C7A3,4);
TASK_PP(16'h1C7A4,4);
TASK_PP(16'h1C7A5,4);
TASK_PP(16'h1C7A6,4);
TASK_PP(16'h1C7A7,4);
TASK_PP(16'h1C7A8,4);
TASK_PP(16'h1C7A9,4);
TASK_PP(16'h1C7AA,4);
TASK_PP(16'h1C7AB,4);
TASK_PP(16'h1C7AC,4);
TASK_PP(16'h1C7AD,4);
TASK_PP(16'h1C7AE,4);
TASK_PP(16'h1C7AF,4);
TASK_PP(16'h1C7B0,4);
TASK_PP(16'h1C7B1,4);
TASK_PP(16'h1C7B2,4);
TASK_PP(16'h1C7B3,4);
TASK_PP(16'h1C7B4,4);
TASK_PP(16'h1C7B5,4);
TASK_PP(16'h1C7B6,4);
TASK_PP(16'h1C7B7,4);
TASK_PP(16'h1C7B8,4);
TASK_PP(16'h1C7B9,4);
TASK_PP(16'h1C7BA,4);
TASK_PP(16'h1C7BB,4);
TASK_PP(16'h1C7BC,4);
TASK_PP(16'h1C7BD,4);
TASK_PP(16'h1C7BE,4);
TASK_PP(16'h1C7BF,4);
TASK_PP(16'h1C7C0,4);
TASK_PP(16'h1C7C1,4);
TASK_PP(16'h1C7C2,4);
TASK_PP(16'h1C7C3,4);
TASK_PP(16'h1C7C4,4);
TASK_PP(16'h1C7C5,4);
TASK_PP(16'h1C7C6,4);
TASK_PP(16'h1C7C7,4);
TASK_PP(16'h1C7C8,4);
TASK_PP(16'h1C7C9,4);
TASK_PP(16'h1C7CA,4);
TASK_PP(16'h1C7CB,4);
TASK_PP(16'h1C7CC,4);
TASK_PP(16'h1C7CD,4);
TASK_PP(16'h1C7CE,4);
TASK_PP(16'h1C7CF,4);
TASK_PP(16'h1C7D0,4);
TASK_PP(16'h1C7D1,4);
TASK_PP(16'h1C7D2,4);
TASK_PP(16'h1C7D3,4);
TASK_PP(16'h1C7D4,4);
TASK_PP(16'h1C7D5,4);
TASK_PP(16'h1C7D6,4);
TASK_PP(16'h1C7D7,4);
TASK_PP(16'h1C7D8,4);
TASK_PP(16'h1C7D9,4);
TASK_PP(16'h1C7DA,4);
TASK_PP(16'h1C7DB,4);
TASK_PP(16'h1C7DC,4);
TASK_PP(16'h1C7DD,4);
TASK_PP(16'h1C7DE,4);
TASK_PP(16'h1C7DF,4);
TASK_PP(16'h1C7E0,4);
TASK_PP(16'h1C7E1,4);
TASK_PP(16'h1C7E2,4);
TASK_PP(16'h1C7E3,4);
TASK_PP(16'h1C7E4,4);
TASK_PP(16'h1C7E5,4);
TASK_PP(16'h1C7E6,4);
TASK_PP(16'h1C7E7,4);
TASK_PP(16'h1C7E8,4);
TASK_PP(16'h1C7E9,4);
TASK_PP(16'h1C7EA,4);
TASK_PP(16'h1C7EB,4);
TASK_PP(16'h1C7EC,4);
TASK_PP(16'h1C7ED,4);
TASK_PP(16'h1C7EE,4);
TASK_PP(16'h1C7EF,4);
TASK_PP(16'h1C7F0,4);
TASK_PP(16'h1C7F1,4);
TASK_PP(16'h1C7F2,4);
TASK_PP(16'h1C7F3,4);
TASK_PP(16'h1C7F4,4);
TASK_PP(16'h1C7F5,4);
TASK_PP(16'h1C7F6,4);
TASK_PP(16'h1C7F7,4);
TASK_PP(16'h1C7F8,4);
TASK_PP(16'h1C7F9,4);
TASK_PP(16'h1C7FA,4);
TASK_PP(16'h1C7FB,4);
TASK_PP(16'h1C7FC,4);
TASK_PP(16'h1C7FD,4);
TASK_PP(16'h1C7FE,4);
TASK_PP(16'h1C7FF,4);
TASK_PP(16'h1C800,4);
TASK_PP(16'h1C801,4);
TASK_PP(16'h1C802,4);
TASK_PP(16'h1C803,4);
TASK_PP(16'h1C804,4);
TASK_PP(16'h1C805,4);
TASK_PP(16'h1C806,4);
TASK_PP(16'h1C807,4);
TASK_PP(16'h1C808,4);
TASK_PP(16'h1C809,4);
TASK_PP(16'h1C80A,4);
TASK_PP(16'h1C80B,4);
TASK_PP(16'h1C80C,4);
TASK_PP(16'h1C80D,4);
TASK_PP(16'h1C80E,4);
TASK_PP(16'h1C80F,4);
TASK_PP(16'h1C810,4);
TASK_PP(16'h1C811,4);
TASK_PP(16'h1C812,4);
TASK_PP(16'h1C813,4);
TASK_PP(16'h1C814,4);
TASK_PP(16'h1C815,4);
TASK_PP(16'h1C816,4);
TASK_PP(16'h1C817,4);
TASK_PP(16'h1C818,4);
TASK_PP(16'h1C819,4);
TASK_PP(16'h1C81A,4);
TASK_PP(16'h1C81B,4);
TASK_PP(16'h1C81C,4);
TASK_PP(16'h1C81D,4);
TASK_PP(16'h1C81E,4);
TASK_PP(16'h1C81F,4);
TASK_PP(16'h1C820,4);
TASK_PP(16'h1C821,4);
TASK_PP(16'h1C822,4);
TASK_PP(16'h1C823,4);
TASK_PP(16'h1C824,4);
TASK_PP(16'h1C825,4);
TASK_PP(16'h1C826,4);
TASK_PP(16'h1C827,4);
TASK_PP(16'h1C828,4);
TASK_PP(16'h1C829,4);
TASK_PP(16'h1C82A,4);
TASK_PP(16'h1C82B,4);
TASK_PP(16'h1C82C,4);
TASK_PP(16'h1C82D,4);
TASK_PP(16'h1C82E,4);
TASK_PP(16'h1C82F,4);
TASK_PP(16'h1C830,4);
TASK_PP(16'h1C831,4);
TASK_PP(16'h1C832,4);
TASK_PP(16'h1C833,4);
TASK_PP(16'h1C834,4);
TASK_PP(16'h1C835,4);
TASK_PP(16'h1C836,4);
TASK_PP(16'h1C837,4);
TASK_PP(16'h1C838,4);
TASK_PP(16'h1C839,4);
TASK_PP(16'h1C83A,4);
TASK_PP(16'h1C83B,4);
TASK_PP(16'h1C83C,4);
TASK_PP(16'h1C83D,4);
TASK_PP(16'h1C83E,4);
TASK_PP(16'h1C83F,4);
TASK_PP(16'h1C840,4);
TASK_PP(16'h1C841,4);
TASK_PP(16'h1C842,4);
TASK_PP(16'h1C843,4);
TASK_PP(16'h1C844,4);
TASK_PP(16'h1C845,4);
TASK_PP(16'h1C846,4);
TASK_PP(16'h1C847,4);
TASK_PP(16'h1C848,4);
TASK_PP(16'h1C849,4);
TASK_PP(16'h1C84A,4);
TASK_PP(16'h1C84B,4);
TASK_PP(16'h1C84C,4);
TASK_PP(16'h1C84D,4);
TASK_PP(16'h1C84E,4);
TASK_PP(16'h1C84F,4);
TASK_PP(16'h1C850,4);
TASK_PP(16'h1C851,4);
TASK_PP(16'h1C852,4);
TASK_PP(16'h1C853,4);
TASK_PP(16'h1C854,4);
TASK_PP(16'h1C855,4);
TASK_PP(16'h1C856,4);
TASK_PP(16'h1C857,4);
TASK_PP(16'h1C858,4);
TASK_PP(16'h1C859,4);
TASK_PP(16'h1C85A,4);
TASK_PP(16'h1C85B,4);
TASK_PP(16'h1C85C,4);
TASK_PP(16'h1C85D,4);
TASK_PP(16'h1C85E,4);
TASK_PP(16'h1C85F,4);
TASK_PP(16'h1C860,4);
TASK_PP(16'h1C861,4);
TASK_PP(16'h1C862,4);
TASK_PP(16'h1C863,4);
TASK_PP(16'h1C864,4);
TASK_PP(16'h1C865,4);
TASK_PP(16'h1C866,4);
TASK_PP(16'h1C867,4);
TASK_PP(16'h1C868,4);
TASK_PP(16'h1C869,4);
TASK_PP(16'h1C86A,4);
TASK_PP(16'h1C86B,4);
TASK_PP(16'h1C86C,4);
TASK_PP(16'h1C86D,4);
TASK_PP(16'h1C86E,4);
TASK_PP(16'h1C86F,4);
TASK_PP(16'h1C870,4);
TASK_PP(16'h1C871,4);
TASK_PP(16'h1C872,4);
TASK_PP(16'h1C873,4);
TASK_PP(16'h1C874,4);
TASK_PP(16'h1C875,4);
TASK_PP(16'h1C876,4);
TASK_PP(16'h1C877,4);
TASK_PP(16'h1C878,4);
TASK_PP(16'h1C879,4);
TASK_PP(16'h1C87A,4);
TASK_PP(16'h1C87B,4);
TASK_PP(16'h1C87C,4);
TASK_PP(16'h1C87D,4);
TASK_PP(16'h1C87E,4);
TASK_PP(16'h1C87F,4);
TASK_PP(16'h1C880,4);
TASK_PP(16'h1C881,4);
TASK_PP(16'h1C882,4);
TASK_PP(16'h1C883,4);
TASK_PP(16'h1C884,4);
TASK_PP(16'h1C885,4);
TASK_PP(16'h1C886,4);
TASK_PP(16'h1C887,4);
TASK_PP(16'h1C888,4);
TASK_PP(16'h1C889,4);
TASK_PP(16'h1C88A,4);
TASK_PP(16'h1C88B,4);
TASK_PP(16'h1C88C,4);
TASK_PP(16'h1C88D,4);
TASK_PP(16'h1C88E,4);
TASK_PP(16'h1C88F,4);
TASK_PP(16'h1C890,4);
TASK_PP(16'h1C891,4);
TASK_PP(16'h1C892,4);
TASK_PP(16'h1C893,4);
TASK_PP(16'h1C894,4);
TASK_PP(16'h1C895,4);
TASK_PP(16'h1C896,4);
TASK_PP(16'h1C897,4);
TASK_PP(16'h1C898,4);
TASK_PP(16'h1C899,4);
TASK_PP(16'h1C89A,4);
TASK_PP(16'h1C89B,4);
TASK_PP(16'h1C89C,4);
TASK_PP(16'h1C89D,4);
TASK_PP(16'h1C89E,4);
TASK_PP(16'h1C89F,4);
TASK_PP(16'h1C8A0,4);
TASK_PP(16'h1C8A1,4);
TASK_PP(16'h1C8A2,4);
TASK_PP(16'h1C8A3,4);
TASK_PP(16'h1C8A4,4);
TASK_PP(16'h1C8A5,4);
TASK_PP(16'h1C8A6,4);
TASK_PP(16'h1C8A7,4);
TASK_PP(16'h1C8A8,4);
TASK_PP(16'h1C8A9,4);
TASK_PP(16'h1C8AA,4);
TASK_PP(16'h1C8AB,4);
TASK_PP(16'h1C8AC,4);
TASK_PP(16'h1C8AD,4);
TASK_PP(16'h1C8AE,4);
TASK_PP(16'h1C8AF,4);
TASK_PP(16'h1C8B0,4);
TASK_PP(16'h1C8B1,4);
TASK_PP(16'h1C8B2,4);
TASK_PP(16'h1C8B3,4);
TASK_PP(16'h1C8B4,4);
TASK_PP(16'h1C8B5,4);
TASK_PP(16'h1C8B6,4);
TASK_PP(16'h1C8B7,4);
TASK_PP(16'h1C8B8,4);
TASK_PP(16'h1C8B9,4);
TASK_PP(16'h1C8BA,4);
TASK_PP(16'h1C8BB,4);
TASK_PP(16'h1C8BC,4);
TASK_PP(16'h1C8BD,4);
TASK_PP(16'h1C8BE,4);
TASK_PP(16'h1C8BF,4);
TASK_PP(16'h1C8C0,4);
TASK_PP(16'h1C8C1,4);
TASK_PP(16'h1C8C2,4);
TASK_PP(16'h1C8C3,4);
TASK_PP(16'h1C8C4,4);
TASK_PP(16'h1C8C5,4);
TASK_PP(16'h1C8C6,4);
TASK_PP(16'h1C8C7,4);
TASK_PP(16'h1C8C8,4);
TASK_PP(16'h1C8C9,4);
TASK_PP(16'h1C8CA,4);
TASK_PP(16'h1C8CB,4);
TASK_PP(16'h1C8CC,4);
TASK_PP(16'h1C8CD,4);
TASK_PP(16'h1C8CE,4);
TASK_PP(16'h1C8CF,4);
TASK_PP(16'h1C8D0,4);
TASK_PP(16'h1C8D1,4);
TASK_PP(16'h1C8D2,4);
TASK_PP(16'h1C8D3,4);
TASK_PP(16'h1C8D4,4);
TASK_PP(16'h1C8D5,4);
TASK_PP(16'h1C8D6,4);
TASK_PP(16'h1C8D7,4);
TASK_PP(16'h1C8D8,4);
TASK_PP(16'h1C8D9,4);
TASK_PP(16'h1C8DA,4);
TASK_PP(16'h1C8DB,4);
TASK_PP(16'h1C8DC,4);
TASK_PP(16'h1C8DD,4);
TASK_PP(16'h1C8DE,4);
TASK_PP(16'h1C8DF,4);
TASK_PP(16'h1C8E0,4);
TASK_PP(16'h1C8E1,4);
TASK_PP(16'h1C8E2,4);
TASK_PP(16'h1C8E3,4);
TASK_PP(16'h1C8E4,4);
TASK_PP(16'h1C8E5,4);
TASK_PP(16'h1C8E6,4);
TASK_PP(16'h1C8E7,4);
TASK_PP(16'h1C8E8,4);
TASK_PP(16'h1C8E9,4);
TASK_PP(16'h1C8EA,4);
TASK_PP(16'h1C8EB,4);
TASK_PP(16'h1C8EC,4);
TASK_PP(16'h1C8ED,4);
TASK_PP(16'h1C8EE,4);
TASK_PP(16'h1C8EF,4);
TASK_PP(16'h1C8F0,4);
TASK_PP(16'h1C8F1,4);
TASK_PP(16'h1C8F2,4);
TASK_PP(16'h1C8F3,4);
TASK_PP(16'h1C8F4,4);
TASK_PP(16'h1C8F5,4);
TASK_PP(16'h1C8F6,4);
TASK_PP(16'h1C8F7,4);
TASK_PP(16'h1C8F8,4);
TASK_PP(16'h1C8F9,4);
TASK_PP(16'h1C8FA,4);
TASK_PP(16'h1C8FB,4);
TASK_PP(16'h1C8FC,4);
TASK_PP(16'h1C8FD,4);
TASK_PP(16'h1C8FE,4);
TASK_PP(16'h1C8FF,4);
TASK_PP(16'h1C900,4);
TASK_PP(16'h1C901,4);
TASK_PP(16'h1C902,4);
TASK_PP(16'h1C903,4);
TASK_PP(16'h1C904,4);
TASK_PP(16'h1C905,4);
TASK_PP(16'h1C906,4);
TASK_PP(16'h1C907,4);
TASK_PP(16'h1C908,4);
TASK_PP(16'h1C909,4);
TASK_PP(16'h1C90A,4);
TASK_PP(16'h1C90B,4);
TASK_PP(16'h1C90C,4);
TASK_PP(16'h1C90D,4);
TASK_PP(16'h1C90E,4);
TASK_PP(16'h1C90F,4);
TASK_PP(16'h1C910,4);
TASK_PP(16'h1C911,4);
TASK_PP(16'h1C912,4);
TASK_PP(16'h1C913,4);
TASK_PP(16'h1C914,4);
TASK_PP(16'h1C915,4);
TASK_PP(16'h1C916,4);
TASK_PP(16'h1C917,4);
TASK_PP(16'h1C918,4);
TASK_PP(16'h1C919,4);
TASK_PP(16'h1C91A,4);
TASK_PP(16'h1C91B,4);
TASK_PP(16'h1C91C,4);
TASK_PP(16'h1C91D,4);
TASK_PP(16'h1C91E,4);
TASK_PP(16'h1C91F,4);
TASK_PP(16'h1C920,4);
TASK_PP(16'h1C921,4);
TASK_PP(16'h1C922,4);
TASK_PP(16'h1C923,4);
TASK_PP(16'h1C924,4);
TASK_PP(16'h1C925,4);
TASK_PP(16'h1C926,4);
TASK_PP(16'h1C927,4);
TASK_PP(16'h1C928,4);
TASK_PP(16'h1C929,4);
TASK_PP(16'h1C92A,4);
TASK_PP(16'h1C92B,4);
TASK_PP(16'h1C92C,4);
TASK_PP(16'h1C92D,4);
TASK_PP(16'h1C92E,4);
TASK_PP(16'h1C92F,4);
TASK_PP(16'h1C930,4);
TASK_PP(16'h1C931,4);
TASK_PP(16'h1C932,4);
TASK_PP(16'h1C933,4);
TASK_PP(16'h1C934,4);
TASK_PP(16'h1C935,4);
TASK_PP(16'h1C936,4);
TASK_PP(16'h1C937,4);
TASK_PP(16'h1C938,4);
TASK_PP(16'h1C939,4);
TASK_PP(16'h1C93A,4);
TASK_PP(16'h1C93B,4);
TASK_PP(16'h1C93C,4);
TASK_PP(16'h1C93D,4);
TASK_PP(16'h1C93E,4);
TASK_PP(16'h1C93F,4);
TASK_PP(16'h1C940,4);
TASK_PP(16'h1C941,4);
TASK_PP(16'h1C942,4);
TASK_PP(16'h1C943,4);
TASK_PP(16'h1C944,4);
TASK_PP(16'h1C945,4);
TASK_PP(16'h1C946,4);
TASK_PP(16'h1C947,4);
TASK_PP(16'h1C948,4);
TASK_PP(16'h1C949,4);
TASK_PP(16'h1C94A,4);
TASK_PP(16'h1C94B,4);
TASK_PP(16'h1C94C,4);
TASK_PP(16'h1C94D,4);
TASK_PP(16'h1C94E,4);
TASK_PP(16'h1C94F,4);
TASK_PP(16'h1C950,4);
TASK_PP(16'h1C951,4);
TASK_PP(16'h1C952,4);
TASK_PP(16'h1C953,4);
TASK_PP(16'h1C954,4);
TASK_PP(16'h1C955,4);
TASK_PP(16'h1C956,4);
TASK_PP(16'h1C957,4);
TASK_PP(16'h1C958,4);
TASK_PP(16'h1C959,4);
TASK_PP(16'h1C95A,4);
TASK_PP(16'h1C95B,4);
TASK_PP(16'h1C95C,4);
TASK_PP(16'h1C95D,4);
TASK_PP(16'h1C95E,4);
TASK_PP(16'h1C95F,4);
TASK_PP(16'h1C960,4);
TASK_PP(16'h1C961,4);
TASK_PP(16'h1C962,4);
TASK_PP(16'h1C963,4);
TASK_PP(16'h1C964,4);
TASK_PP(16'h1C965,4);
TASK_PP(16'h1C966,4);
TASK_PP(16'h1C967,4);
TASK_PP(16'h1C968,4);
TASK_PP(16'h1C969,4);
TASK_PP(16'h1C96A,4);
TASK_PP(16'h1C96B,4);
TASK_PP(16'h1C96C,4);
TASK_PP(16'h1C96D,4);
TASK_PP(16'h1C96E,4);
TASK_PP(16'h1C96F,4);
TASK_PP(16'h1C970,4);
TASK_PP(16'h1C971,4);
TASK_PP(16'h1C972,4);
TASK_PP(16'h1C973,4);
TASK_PP(16'h1C974,4);
TASK_PP(16'h1C975,4);
TASK_PP(16'h1C976,4);
TASK_PP(16'h1C977,4);
TASK_PP(16'h1C978,4);
TASK_PP(16'h1C979,4);
TASK_PP(16'h1C97A,4);
TASK_PP(16'h1C97B,4);
TASK_PP(16'h1C97C,4);
TASK_PP(16'h1C97D,4);
TASK_PP(16'h1C97E,4);
TASK_PP(16'h1C97F,4);
TASK_PP(16'h1C980,4);
TASK_PP(16'h1C981,4);
TASK_PP(16'h1C982,4);
TASK_PP(16'h1C983,4);
TASK_PP(16'h1C984,4);
TASK_PP(16'h1C985,4);
TASK_PP(16'h1C986,4);
TASK_PP(16'h1C987,4);
TASK_PP(16'h1C988,4);
TASK_PP(16'h1C989,4);
TASK_PP(16'h1C98A,4);
TASK_PP(16'h1C98B,4);
TASK_PP(16'h1C98C,4);
TASK_PP(16'h1C98D,4);
TASK_PP(16'h1C98E,4);
TASK_PP(16'h1C98F,4);
TASK_PP(16'h1C990,4);
TASK_PP(16'h1C991,4);
TASK_PP(16'h1C992,4);
TASK_PP(16'h1C993,4);
TASK_PP(16'h1C994,4);
TASK_PP(16'h1C995,4);
TASK_PP(16'h1C996,4);
TASK_PP(16'h1C997,4);
TASK_PP(16'h1C998,4);
TASK_PP(16'h1C999,4);
TASK_PP(16'h1C99A,4);
TASK_PP(16'h1C99B,4);
TASK_PP(16'h1C99C,4);
TASK_PP(16'h1C99D,4);
TASK_PP(16'h1C99E,4);
TASK_PP(16'h1C99F,4);
TASK_PP(16'h1C9A0,4);
TASK_PP(16'h1C9A1,4);
TASK_PP(16'h1C9A2,4);
TASK_PP(16'h1C9A3,4);
TASK_PP(16'h1C9A4,4);
TASK_PP(16'h1C9A5,4);
TASK_PP(16'h1C9A6,4);
TASK_PP(16'h1C9A7,4);
TASK_PP(16'h1C9A8,4);
TASK_PP(16'h1C9A9,4);
TASK_PP(16'h1C9AA,4);
TASK_PP(16'h1C9AB,4);
TASK_PP(16'h1C9AC,4);
TASK_PP(16'h1C9AD,4);
TASK_PP(16'h1C9AE,4);
TASK_PP(16'h1C9AF,4);
TASK_PP(16'h1C9B0,4);
TASK_PP(16'h1C9B1,4);
TASK_PP(16'h1C9B2,4);
TASK_PP(16'h1C9B3,4);
TASK_PP(16'h1C9B4,4);
TASK_PP(16'h1C9B5,4);
TASK_PP(16'h1C9B6,4);
TASK_PP(16'h1C9B7,4);
TASK_PP(16'h1C9B8,4);
TASK_PP(16'h1C9B9,4);
TASK_PP(16'h1C9BA,4);
TASK_PP(16'h1C9BB,4);
TASK_PP(16'h1C9BC,4);
TASK_PP(16'h1C9BD,4);
TASK_PP(16'h1C9BE,4);
TASK_PP(16'h1C9BF,4);
TASK_PP(16'h1C9C0,4);
TASK_PP(16'h1C9C1,4);
TASK_PP(16'h1C9C2,4);
TASK_PP(16'h1C9C3,4);
TASK_PP(16'h1C9C4,4);
TASK_PP(16'h1C9C5,4);
TASK_PP(16'h1C9C6,4);
TASK_PP(16'h1C9C7,4);
TASK_PP(16'h1C9C8,4);
TASK_PP(16'h1C9C9,4);
TASK_PP(16'h1C9CA,4);
TASK_PP(16'h1C9CB,4);
TASK_PP(16'h1C9CC,4);
TASK_PP(16'h1C9CD,4);
TASK_PP(16'h1C9CE,4);
TASK_PP(16'h1C9CF,4);
TASK_PP(16'h1C9D0,4);
TASK_PP(16'h1C9D1,4);
TASK_PP(16'h1C9D2,4);
TASK_PP(16'h1C9D3,4);
TASK_PP(16'h1C9D4,4);
TASK_PP(16'h1C9D5,4);
TASK_PP(16'h1C9D6,4);
TASK_PP(16'h1C9D7,4);
TASK_PP(16'h1C9D8,4);
TASK_PP(16'h1C9D9,4);
TASK_PP(16'h1C9DA,4);
TASK_PP(16'h1C9DB,4);
TASK_PP(16'h1C9DC,4);
TASK_PP(16'h1C9DD,4);
TASK_PP(16'h1C9DE,4);
TASK_PP(16'h1C9DF,4);
TASK_PP(16'h1C9E0,4);
TASK_PP(16'h1C9E1,4);
TASK_PP(16'h1C9E2,4);
TASK_PP(16'h1C9E3,4);
TASK_PP(16'h1C9E4,4);
TASK_PP(16'h1C9E5,4);
TASK_PP(16'h1C9E6,4);
TASK_PP(16'h1C9E7,4);
TASK_PP(16'h1C9E8,4);
TASK_PP(16'h1C9E9,4);
TASK_PP(16'h1C9EA,4);
TASK_PP(16'h1C9EB,4);
TASK_PP(16'h1C9EC,4);
TASK_PP(16'h1C9ED,4);
TASK_PP(16'h1C9EE,4);
TASK_PP(16'h1C9EF,4);
TASK_PP(16'h1C9F0,4);
TASK_PP(16'h1C9F1,4);
TASK_PP(16'h1C9F2,4);
TASK_PP(16'h1C9F3,4);
TASK_PP(16'h1C9F4,4);
TASK_PP(16'h1C9F5,4);
TASK_PP(16'h1C9F6,4);
TASK_PP(16'h1C9F7,4);
TASK_PP(16'h1C9F8,4);
TASK_PP(16'h1C9F9,4);
TASK_PP(16'h1C9FA,4);
TASK_PP(16'h1C9FB,4);
TASK_PP(16'h1C9FC,4);
TASK_PP(16'h1C9FD,4);
TASK_PP(16'h1C9FE,4);
TASK_PP(16'h1C9FF,4);
TASK_PP(16'h1CA00,4);
TASK_PP(16'h1CA01,4);
TASK_PP(16'h1CA02,4);
TASK_PP(16'h1CA03,4);
TASK_PP(16'h1CA04,4);
TASK_PP(16'h1CA05,4);
TASK_PP(16'h1CA06,4);
TASK_PP(16'h1CA07,4);
TASK_PP(16'h1CA08,4);
TASK_PP(16'h1CA09,4);
TASK_PP(16'h1CA0A,4);
TASK_PP(16'h1CA0B,4);
TASK_PP(16'h1CA0C,4);
TASK_PP(16'h1CA0D,4);
TASK_PP(16'h1CA0E,4);
TASK_PP(16'h1CA0F,4);
TASK_PP(16'h1CA10,4);
TASK_PP(16'h1CA11,4);
TASK_PP(16'h1CA12,4);
TASK_PP(16'h1CA13,4);
TASK_PP(16'h1CA14,4);
TASK_PP(16'h1CA15,4);
TASK_PP(16'h1CA16,4);
TASK_PP(16'h1CA17,4);
TASK_PP(16'h1CA18,4);
TASK_PP(16'h1CA19,4);
TASK_PP(16'h1CA1A,4);
TASK_PP(16'h1CA1B,4);
TASK_PP(16'h1CA1C,4);
TASK_PP(16'h1CA1D,4);
TASK_PP(16'h1CA1E,4);
TASK_PP(16'h1CA1F,4);
TASK_PP(16'h1CA20,4);
TASK_PP(16'h1CA21,4);
TASK_PP(16'h1CA22,4);
TASK_PP(16'h1CA23,4);
TASK_PP(16'h1CA24,4);
TASK_PP(16'h1CA25,4);
TASK_PP(16'h1CA26,4);
TASK_PP(16'h1CA27,4);
TASK_PP(16'h1CA28,4);
TASK_PP(16'h1CA29,4);
TASK_PP(16'h1CA2A,4);
TASK_PP(16'h1CA2B,4);
TASK_PP(16'h1CA2C,4);
TASK_PP(16'h1CA2D,4);
TASK_PP(16'h1CA2E,4);
TASK_PP(16'h1CA2F,4);
TASK_PP(16'h1CA30,4);
TASK_PP(16'h1CA31,4);
TASK_PP(16'h1CA32,4);
TASK_PP(16'h1CA33,4);
TASK_PP(16'h1CA34,4);
TASK_PP(16'h1CA35,4);
TASK_PP(16'h1CA36,4);
TASK_PP(16'h1CA37,4);
TASK_PP(16'h1CA38,4);
TASK_PP(16'h1CA39,4);
TASK_PP(16'h1CA3A,4);
TASK_PP(16'h1CA3B,4);
TASK_PP(16'h1CA3C,4);
TASK_PP(16'h1CA3D,4);
TASK_PP(16'h1CA3E,4);
TASK_PP(16'h1CA3F,4);
TASK_PP(16'h1CA40,4);
TASK_PP(16'h1CA41,4);
TASK_PP(16'h1CA42,4);
TASK_PP(16'h1CA43,4);
TASK_PP(16'h1CA44,4);
TASK_PP(16'h1CA45,4);
TASK_PP(16'h1CA46,4);
TASK_PP(16'h1CA47,4);
TASK_PP(16'h1CA48,4);
TASK_PP(16'h1CA49,4);
TASK_PP(16'h1CA4A,4);
TASK_PP(16'h1CA4B,4);
TASK_PP(16'h1CA4C,4);
TASK_PP(16'h1CA4D,4);
TASK_PP(16'h1CA4E,4);
TASK_PP(16'h1CA4F,4);
TASK_PP(16'h1CA50,4);
TASK_PP(16'h1CA51,4);
TASK_PP(16'h1CA52,4);
TASK_PP(16'h1CA53,4);
TASK_PP(16'h1CA54,4);
TASK_PP(16'h1CA55,4);
TASK_PP(16'h1CA56,4);
TASK_PP(16'h1CA57,4);
TASK_PP(16'h1CA58,4);
TASK_PP(16'h1CA59,4);
TASK_PP(16'h1CA5A,4);
TASK_PP(16'h1CA5B,4);
TASK_PP(16'h1CA5C,4);
TASK_PP(16'h1CA5D,4);
TASK_PP(16'h1CA5E,4);
TASK_PP(16'h1CA5F,4);
TASK_PP(16'h1CA60,4);
TASK_PP(16'h1CA61,4);
TASK_PP(16'h1CA62,4);
TASK_PP(16'h1CA63,4);
TASK_PP(16'h1CA64,4);
TASK_PP(16'h1CA65,4);
TASK_PP(16'h1CA66,4);
TASK_PP(16'h1CA67,4);
TASK_PP(16'h1CA68,4);
TASK_PP(16'h1CA69,4);
TASK_PP(16'h1CA6A,4);
TASK_PP(16'h1CA6B,4);
TASK_PP(16'h1CA6C,4);
TASK_PP(16'h1CA6D,4);
TASK_PP(16'h1CA6E,4);
TASK_PP(16'h1CA6F,4);
TASK_PP(16'h1CA70,4);
TASK_PP(16'h1CA71,4);
TASK_PP(16'h1CA72,4);
TASK_PP(16'h1CA73,4);
TASK_PP(16'h1CA74,4);
TASK_PP(16'h1CA75,4);
TASK_PP(16'h1CA76,4);
TASK_PP(16'h1CA77,4);
TASK_PP(16'h1CA78,4);
TASK_PP(16'h1CA79,4);
TASK_PP(16'h1CA7A,4);
TASK_PP(16'h1CA7B,4);
TASK_PP(16'h1CA7C,4);
TASK_PP(16'h1CA7D,4);
TASK_PP(16'h1CA7E,4);
TASK_PP(16'h1CA7F,4);
TASK_PP(16'h1CA80,4);
TASK_PP(16'h1CA81,4);
TASK_PP(16'h1CA82,4);
TASK_PP(16'h1CA83,4);
TASK_PP(16'h1CA84,4);
TASK_PP(16'h1CA85,4);
TASK_PP(16'h1CA86,4);
TASK_PP(16'h1CA87,4);
TASK_PP(16'h1CA88,4);
TASK_PP(16'h1CA89,4);
TASK_PP(16'h1CA8A,4);
TASK_PP(16'h1CA8B,4);
TASK_PP(16'h1CA8C,4);
TASK_PP(16'h1CA8D,4);
TASK_PP(16'h1CA8E,4);
TASK_PP(16'h1CA8F,4);
TASK_PP(16'h1CA90,4);
TASK_PP(16'h1CA91,4);
TASK_PP(16'h1CA92,4);
TASK_PP(16'h1CA93,4);
TASK_PP(16'h1CA94,4);
TASK_PP(16'h1CA95,4);
TASK_PP(16'h1CA96,4);
TASK_PP(16'h1CA97,4);
TASK_PP(16'h1CA98,4);
TASK_PP(16'h1CA99,4);
TASK_PP(16'h1CA9A,4);
TASK_PP(16'h1CA9B,4);
TASK_PP(16'h1CA9C,4);
TASK_PP(16'h1CA9D,4);
TASK_PP(16'h1CA9E,4);
TASK_PP(16'h1CA9F,4);
TASK_PP(16'h1CAA0,4);
TASK_PP(16'h1CAA1,4);
TASK_PP(16'h1CAA2,4);
TASK_PP(16'h1CAA3,4);
TASK_PP(16'h1CAA4,4);
TASK_PP(16'h1CAA5,4);
TASK_PP(16'h1CAA6,4);
TASK_PP(16'h1CAA7,4);
TASK_PP(16'h1CAA8,4);
TASK_PP(16'h1CAA9,4);
TASK_PP(16'h1CAAA,4);
TASK_PP(16'h1CAAB,4);
TASK_PP(16'h1CAAC,4);
TASK_PP(16'h1CAAD,4);
TASK_PP(16'h1CAAE,4);
TASK_PP(16'h1CAAF,4);
TASK_PP(16'h1CAB0,4);
TASK_PP(16'h1CAB1,4);
TASK_PP(16'h1CAB2,4);
TASK_PP(16'h1CAB3,4);
TASK_PP(16'h1CAB4,4);
TASK_PP(16'h1CAB5,4);
TASK_PP(16'h1CAB6,4);
TASK_PP(16'h1CAB7,4);
TASK_PP(16'h1CAB8,4);
TASK_PP(16'h1CAB9,4);
TASK_PP(16'h1CABA,4);
TASK_PP(16'h1CABB,4);
TASK_PP(16'h1CABC,4);
TASK_PP(16'h1CABD,4);
TASK_PP(16'h1CABE,4);
TASK_PP(16'h1CABF,4);
TASK_PP(16'h1CAC0,4);
TASK_PP(16'h1CAC1,4);
TASK_PP(16'h1CAC2,4);
TASK_PP(16'h1CAC3,4);
TASK_PP(16'h1CAC4,4);
TASK_PP(16'h1CAC5,4);
TASK_PP(16'h1CAC6,4);
TASK_PP(16'h1CAC7,4);
TASK_PP(16'h1CAC8,4);
TASK_PP(16'h1CAC9,4);
TASK_PP(16'h1CACA,4);
TASK_PP(16'h1CACB,4);
TASK_PP(16'h1CACC,4);
TASK_PP(16'h1CACD,4);
TASK_PP(16'h1CACE,4);
TASK_PP(16'h1CACF,4);
TASK_PP(16'h1CAD0,4);
TASK_PP(16'h1CAD1,4);
TASK_PP(16'h1CAD2,4);
TASK_PP(16'h1CAD3,4);
TASK_PP(16'h1CAD4,4);
TASK_PP(16'h1CAD5,4);
TASK_PP(16'h1CAD6,4);
TASK_PP(16'h1CAD7,4);
TASK_PP(16'h1CAD8,4);
TASK_PP(16'h1CAD9,4);
TASK_PP(16'h1CADA,4);
TASK_PP(16'h1CADB,4);
TASK_PP(16'h1CADC,4);
TASK_PP(16'h1CADD,4);
TASK_PP(16'h1CADE,4);
TASK_PP(16'h1CADF,4);
TASK_PP(16'h1CAE0,4);
TASK_PP(16'h1CAE1,4);
TASK_PP(16'h1CAE2,4);
TASK_PP(16'h1CAE3,4);
TASK_PP(16'h1CAE4,4);
TASK_PP(16'h1CAE5,4);
TASK_PP(16'h1CAE6,4);
TASK_PP(16'h1CAE7,4);
TASK_PP(16'h1CAE8,4);
TASK_PP(16'h1CAE9,4);
TASK_PP(16'h1CAEA,4);
TASK_PP(16'h1CAEB,4);
TASK_PP(16'h1CAEC,4);
TASK_PP(16'h1CAED,4);
TASK_PP(16'h1CAEE,4);
TASK_PP(16'h1CAEF,4);
TASK_PP(16'h1CAF0,4);
TASK_PP(16'h1CAF1,4);
TASK_PP(16'h1CAF2,4);
TASK_PP(16'h1CAF3,4);
TASK_PP(16'h1CAF4,4);
TASK_PP(16'h1CAF5,4);
TASK_PP(16'h1CAF6,4);
TASK_PP(16'h1CAF7,4);
TASK_PP(16'h1CAF8,4);
TASK_PP(16'h1CAF9,4);
TASK_PP(16'h1CAFA,4);
TASK_PP(16'h1CAFB,4);
TASK_PP(16'h1CAFC,4);
TASK_PP(16'h1CAFD,4);
TASK_PP(16'h1CAFE,4);
TASK_PP(16'h1CAFF,4);
TASK_PP(16'h1CB00,4);
TASK_PP(16'h1CB01,4);
TASK_PP(16'h1CB02,4);
TASK_PP(16'h1CB03,4);
TASK_PP(16'h1CB04,4);
TASK_PP(16'h1CB05,4);
TASK_PP(16'h1CB06,4);
TASK_PP(16'h1CB07,4);
TASK_PP(16'h1CB08,4);
TASK_PP(16'h1CB09,4);
TASK_PP(16'h1CB0A,4);
TASK_PP(16'h1CB0B,4);
TASK_PP(16'h1CB0C,4);
TASK_PP(16'h1CB0D,4);
TASK_PP(16'h1CB0E,4);
TASK_PP(16'h1CB0F,4);
TASK_PP(16'h1CB10,4);
TASK_PP(16'h1CB11,4);
TASK_PP(16'h1CB12,4);
TASK_PP(16'h1CB13,4);
TASK_PP(16'h1CB14,4);
TASK_PP(16'h1CB15,4);
TASK_PP(16'h1CB16,4);
TASK_PP(16'h1CB17,4);
TASK_PP(16'h1CB18,4);
TASK_PP(16'h1CB19,4);
TASK_PP(16'h1CB1A,4);
TASK_PP(16'h1CB1B,4);
TASK_PP(16'h1CB1C,4);
TASK_PP(16'h1CB1D,4);
TASK_PP(16'h1CB1E,4);
TASK_PP(16'h1CB1F,4);
TASK_PP(16'h1CB20,4);
TASK_PP(16'h1CB21,4);
TASK_PP(16'h1CB22,4);
TASK_PP(16'h1CB23,4);
TASK_PP(16'h1CB24,4);
TASK_PP(16'h1CB25,4);
TASK_PP(16'h1CB26,4);
TASK_PP(16'h1CB27,4);
TASK_PP(16'h1CB28,4);
TASK_PP(16'h1CB29,4);
TASK_PP(16'h1CB2A,4);
TASK_PP(16'h1CB2B,4);
TASK_PP(16'h1CB2C,4);
TASK_PP(16'h1CB2D,4);
TASK_PP(16'h1CB2E,4);
TASK_PP(16'h1CB2F,4);
TASK_PP(16'h1CB30,4);
TASK_PP(16'h1CB31,4);
TASK_PP(16'h1CB32,4);
TASK_PP(16'h1CB33,4);
TASK_PP(16'h1CB34,4);
TASK_PP(16'h1CB35,4);
TASK_PP(16'h1CB36,4);
TASK_PP(16'h1CB37,4);
TASK_PP(16'h1CB38,4);
TASK_PP(16'h1CB39,4);
TASK_PP(16'h1CB3A,4);
TASK_PP(16'h1CB3B,4);
TASK_PP(16'h1CB3C,4);
TASK_PP(16'h1CB3D,4);
TASK_PP(16'h1CB3E,4);
TASK_PP(16'h1CB3F,4);
TASK_PP(16'h1CB40,4);
TASK_PP(16'h1CB41,4);
TASK_PP(16'h1CB42,4);
TASK_PP(16'h1CB43,4);
TASK_PP(16'h1CB44,4);
TASK_PP(16'h1CB45,4);
TASK_PP(16'h1CB46,4);
TASK_PP(16'h1CB47,4);
TASK_PP(16'h1CB48,4);
TASK_PP(16'h1CB49,4);
TASK_PP(16'h1CB4A,4);
TASK_PP(16'h1CB4B,4);
TASK_PP(16'h1CB4C,4);
TASK_PP(16'h1CB4D,4);
TASK_PP(16'h1CB4E,4);
TASK_PP(16'h1CB4F,4);
TASK_PP(16'h1CB50,4);
TASK_PP(16'h1CB51,4);
TASK_PP(16'h1CB52,4);
TASK_PP(16'h1CB53,4);
TASK_PP(16'h1CB54,4);
TASK_PP(16'h1CB55,4);
TASK_PP(16'h1CB56,4);
TASK_PP(16'h1CB57,4);
TASK_PP(16'h1CB58,4);
TASK_PP(16'h1CB59,4);
TASK_PP(16'h1CB5A,4);
TASK_PP(16'h1CB5B,4);
TASK_PP(16'h1CB5C,4);
TASK_PP(16'h1CB5D,4);
TASK_PP(16'h1CB5E,4);
TASK_PP(16'h1CB5F,4);
TASK_PP(16'h1CB60,4);
TASK_PP(16'h1CB61,4);
TASK_PP(16'h1CB62,4);
TASK_PP(16'h1CB63,4);
TASK_PP(16'h1CB64,4);
TASK_PP(16'h1CB65,4);
TASK_PP(16'h1CB66,4);
TASK_PP(16'h1CB67,4);
TASK_PP(16'h1CB68,4);
TASK_PP(16'h1CB69,4);
TASK_PP(16'h1CB6A,4);
TASK_PP(16'h1CB6B,4);
TASK_PP(16'h1CB6C,4);
TASK_PP(16'h1CB6D,4);
TASK_PP(16'h1CB6E,4);
TASK_PP(16'h1CB6F,4);
TASK_PP(16'h1CB70,4);
TASK_PP(16'h1CB71,4);
TASK_PP(16'h1CB72,4);
TASK_PP(16'h1CB73,4);
TASK_PP(16'h1CB74,4);
TASK_PP(16'h1CB75,4);
TASK_PP(16'h1CB76,4);
TASK_PP(16'h1CB77,4);
TASK_PP(16'h1CB78,4);
TASK_PP(16'h1CB79,4);
TASK_PP(16'h1CB7A,4);
TASK_PP(16'h1CB7B,4);
TASK_PP(16'h1CB7C,4);
TASK_PP(16'h1CB7D,4);
TASK_PP(16'h1CB7E,4);
TASK_PP(16'h1CB7F,4);
TASK_PP(16'h1CB80,4);
TASK_PP(16'h1CB81,4);
TASK_PP(16'h1CB82,4);
TASK_PP(16'h1CB83,4);
TASK_PP(16'h1CB84,4);
TASK_PP(16'h1CB85,4);
TASK_PP(16'h1CB86,4);
TASK_PP(16'h1CB87,4);
TASK_PP(16'h1CB88,4);
TASK_PP(16'h1CB89,4);
TASK_PP(16'h1CB8A,4);
TASK_PP(16'h1CB8B,4);
TASK_PP(16'h1CB8C,4);
TASK_PP(16'h1CB8D,4);
TASK_PP(16'h1CB8E,4);
TASK_PP(16'h1CB8F,4);
TASK_PP(16'h1CB90,4);
TASK_PP(16'h1CB91,4);
TASK_PP(16'h1CB92,4);
TASK_PP(16'h1CB93,4);
TASK_PP(16'h1CB94,4);
TASK_PP(16'h1CB95,4);
TASK_PP(16'h1CB96,4);
TASK_PP(16'h1CB97,4);
TASK_PP(16'h1CB98,4);
TASK_PP(16'h1CB99,4);
TASK_PP(16'h1CB9A,4);
TASK_PP(16'h1CB9B,4);
TASK_PP(16'h1CB9C,4);
TASK_PP(16'h1CB9D,4);
TASK_PP(16'h1CB9E,4);
TASK_PP(16'h1CB9F,4);
TASK_PP(16'h1CBA0,4);
TASK_PP(16'h1CBA1,4);
TASK_PP(16'h1CBA2,4);
TASK_PP(16'h1CBA3,4);
TASK_PP(16'h1CBA4,4);
TASK_PP(16'h1CBA5,4);
TASK_PP(16'h1CBA6,4);
TASK_PP(16'h1CBA7,4);
TASK_PP(16'h1CBA8,4);
TASK_PP(16'h1CBA9,4);
TASK_PP(16'h1CBAA,4);
TASK_PP(16'h1CBAB,4);
TASK_PP(16'h1CBAC,4);
TASK_PP(16'h1CBAD,4);
TASK_PP(16'h1CBAE,4);
TASK_PP(16'h1CBAF,4);
TASK_PP(16'h1CBB0,4);
TASK_PP(16'h1CBB1,4);
TASK_PP(16'h1CBB2,4);
TASK_PP(16'h1CBB3,4);
TASK_PP(16'h1CBB4,4);
TASK_PP(16'h1CBB5,4);
TASK_PP(16'h1CBB6,4);
TASK_PP(16'h1CBB7,4);
TASK_PP(16'h1CBB8,4);
TASK_PP(16'h1CBB9,4);
TASK_PP(16'h1CBBA,4);
TASK_PP(16'h1CBBB,4);
TASK_PP(16'h1CBBC,4);
TASK_PP(16'h1CBBD,4);
TASK_PP(16'h1CBBE,4);
TASK_PP(16'h1CBBF,4);
TASK_PP(16'h1CBC0,4);
TASK_PP(16'h1CBC1,4);
TASK_PP(16'h1CBC2,4);
TASK_PP(16'h1CBC3,4);
TASK_PP(16'h1CBC4,4);
TASK_PP(16'h1CBC5,4);
TASK_PP(16'h1CBC6,4);
TASK_PP(16'h1CBC7,4);
TASK_PP(16'h1CBC8,4);
TASK_PP(16'h1CBC9,4);
TASK_PP(16'h1CBCA,4);
TASK_PP(16'h1CBCB,4);
TASK_PP(16'h1CBCC,4);
TASK_PP(16'h1CBCD,4);
TASK_PP(16'h1CBCE,4);
TASK_PP(16'h1CBCF,4);
TASK_PP(16'h1CBD0,4);
TASK_PP(16'h1CBD1,4);
TASK_PP(16'h1CBD2,4);
TASK_PP(16'h1CBD3,4);
TASK_PP(16'h1CBD4,4);
TASK_PP(16'h1CBD5,4);
TASK_PP(16'h1CBD6,4);
TASK_PP(16'h1CBD7,4);
TASK_PP(16'h1CBD8,4);
TASK_PP(16'h1CBD9,4);
TASK_PP(16'h1CBDA,4);
TASK_PP(16'h1CBDB,4);
TASK_PP(16'h1CBDC,4);
TASK_PP(16'h1CBDD,4);
TASK_PP(16'h1CBDE,4);
TASK_PP(16'h1CBDF,4);
TASK_PP(16'h1CBE0,4);
TASK_PP(16'h1CBE1,4);
TASK_PP(16'h1CBE2,4);
TASK_PP(16'h1CBE3,4);
TASK_PP(16'h1CBE4,4);
TASK_PP(16'h1CBE5,4);
TASK_PP(16'h1CBE6,4);
TASK_PP(16'h1CBE7,4);
TASK_PP(16'h1CBE8,4);
TASK_PP(16'h1CBE9,4);
TASK_PP(16'h1CBEA,4);
TASK_PP(16'h1CBEB,4);
TASK_PP(16'h1CBEC,4);
TASK_PP(16'h1CBED,4);
TASK_PP(16'h1CBEE,4);
TASK_PP(16'h1CBEF,4);
TASK_PP(16'h1CBF0,4);
TASK_PP(16'h1CBF1,4);
TASK_PP(16'h1CBF2,4);
TASK_PP(16'h1CBF3,4);
TASK_PP(16'h1CBF4,4);
TASK_PP(16'h1CBF5,4);
TASK_PP(16'h1CBF6,4);
TASK_PP(16'h1CBF7,4);
TASK_PP(16'h1CBF8,4);
TASK_PP(16'h1CBF9,4);
TASK_PP(16'h1CBFA,4);
TASK_PP(16'h1CBFB,4);
TASK_PP(16'h1CBFC,4);
TASK_PP(16'h1CBFD,4);
TASK_PP(16'h1CBFE,4);
TASK_PP(16'h1CBFF,4);
TASK_PP(16'h1CC00,4);
TASK_PP(16'h1CC01,4);
TASK_PP(16'h1CC02,4);
TASK_PP(16'h1CC03,4);
TASK_PP(16'h1CC04,4);
TASK_PP(16'h1CC05,4);
TASK_PP(16'h1CC06,4);
TASK_PP(16'h1CC07,4);
TASK_PP(16'h1CC08,4);
TASK_PP(16'h1CC09,4);
TASK_PP(16'h1CC0A,4);
TASK_PP(16'h1CC0B,4);
TASK_PP(16'h1CC0C,4);
TASK_PP(16'h1CC0D,4);
TASK_PP(16'h1CC0E,4);
TASK_PP(16'h1CC0F,4);
TASK_PP(16'h1CC10,4);
TASK_PP(16'h1CC11,4);
TASK_PP(16'h1CC12,4);
TASK_PP(16'h1CC13,4);
TASK_PP(16'h1CC14,4);
TASK_PP(16'h1CC15,4);
TASK_PP(16'h1CC16,4);
TASK_PP(16'h1CC17,4);
TASK_PP(16'h1CC18,4);
TASK_PP(16'h1CC19,4);
TASK_PP(16'h1CC1A,4);
TASK_PP(16'h1CC1B,4);
TASK_PP(16'h1CC1C,4);
TASK_PP(16'h1CC1D,4);
TASK_PP(16'h1CC1E,4);
TASK_PP(16'h1CC1F,4);
TASK_PP(16'h1CC20,4);
TASK_PP(16'h1CC21,4);
TASK_PP(16'h1CC22,4);
TASK_PP(16'h1CC23,4);
TASK_PP(16'h1CC24,4);
TASK_PP(16'h1CC25,4);
TASK_PP(16'h1CC26,4);
TASK_PP(16'h1CC27,4);
TASK_PP(16'h1CC28,4);
TASK_PP(16'h1CC29,4);
TASK_PP(16'h1CC2A,4);
TASK_PP(16'h1CC2B,4);
TASK_PP(16'h1CC2C,4);
TASK_PP(16'h1CC2D,4);
TASK_PP(16'h1CC2E,4);
TASK_PP(16'h1CC2F,4);
TASK_PP(16'h1CC30,4);
TASK_PP(16'h1CC31,4);
TASK_PP(16'h1CC32,4);
TASK_PP(16'h1CC33,4);
TASK_PP(16'h1CC34,4);
TASK_PP(16'h1CC35,4);
TASK_PP(16'h1CC36,4);
TASK_PP(16'h1CC37,4);
TASK_PP(16'h1CC38,4);
TASK_PP(16'h1CC39,4);
TASK_PP(16'h1CC3A,4);
TASK_PP(16'h1CC3B,4);
TASK_PP(16'h1CC3C,4);
TASK_PP(16'h1CC3D,4);
TASK_PP(16'h1CC3E,4);
TASK_PP(16'h1CC3F,4);
TASK_PP(16'h1CC40,4);
TASK_PP(16'h1CC41,4);
TASK_PP(16'h1CC42,4);
TASK_PP(16'h1CC43,4);
TASK_PP(16'h1CC44,4);
TASK_PP(16'h1CC45,4);
TASK_PP(16'h1CC46,4);
TASK_PP(16'h1CC47,4);
TASK_PP(16'h1CC48,4);
TASK_PP(16'h1CC49,4);
TASK_PP(16'h1CC4A,4);
TASK_PP(16'h1CC4B,4);
TASK_PP(16'h1CC4C,4);
TASK_PP(16'h1CC4D,4);
TASK_PP(16'h1CC4E,4);
TASK_PP(16'h1CC4F,4);
TASK_PP(16'h1CC50,4);
TASK_PP(16'h1CC51,4);
TASK_PP(16'h1CC52,4);
TASK_PP(16'h1CC53,4);
TASK_PP(16'h1CC54,4);
TASK_PP(16'h1CC55,4);
TASK_PP(16'h1CC56,4);
TASK_PP(16'h1CC57,4);
TASK_PP(16'h1CC58,4);
TASK_PP(16'h1CC59,4);
TASK_PP(16'h1CC5A,4);
TASK_PP(16'h1CC5B,4);
TASK_PP(16'h1CC5C,4);
TASK_PP(16'h1CC5D,4);
TASK_PP(16'h1CC5E,4);
TASK_PP(16'h1CC5F,4);
TASK_PP(16'h1CC60,4);
TASK_PP(16'h1CC61,4);
TASK_PP(16'h1CC62,4);
TASK_PP(16'h1CC63,4);
TASK_PP(16'h1CC64,4);
TASK_PP(16'h1CC65,4);
TASK_PP(16'h1CC66,4);
TASK_PP(16'h1CC67,4);
TASK_PP(16'h1CC68,4);
TASK_PP(16'h1CC69,4);
TASK_PP(16'h1CC6A,4);
TASK_PP(16'h1CC6B,4);
TASK_PP(16'h1CC6C,4);
TASK_PP(16'h1CC6D,4);
TASK_PP(16'h1CC6E,4);
TASK_PP(16'h1CC6F,4);
TASK_PP(16'h1CC70,4);
TASK_PP(16'h1CC71,4);
TASK_PP(16'h1CC72,4);
TASK_PP(16'h1CC73,4);
TASK_PP(16'h1CC74,4);
TASK_PP(16'h1CC75,4);
TASK_PP(16'h1CC76,4);
TASK_PP(16'h1CC77,4);
TASK_PP(16'h1CC78,4);
TASK_PP(16'h1CC79,4);
TASK_PP(16'h1CC7A,4);
TASK_PP(16'h1CC7B,4);
TASK_PP(16'h1CC7C,4);
TASK_PP(16'h1CC7D,4);
TASK_PP(16'h1CC7E,4);
TASK_PP(16'h1CC7F,4);
TASK_PP(16'h1CC80,4);
TASK_PP(16'h1CC81,4);
TASK_PP(16'h1CC82,4);
TASK_PP(16'h1CC83,4);
TASK_PP(16'h1CC84,4);
TASK_PP(16'h1CC85,4);
TASK_PP(16'h1CC86,4);
TASK_PP(16'h1CC87,4);
TASK_PP(16'h1CC88,4);
TASK_PP(16'h1CC89,4);
TASK_PP(16'h1CC8A,4);
TASK_PP(16'h1CC8B,4);
TASK_PP(16'h1CC8C,4);
TASK_PP(16'h1CC8D,4);
TASK_PP(16'h1CC8E,4);
TASK_PP(16'h1CC8F,4);
TASK_PP(16'h1CC90,4);
TASK_PP(16'h1CC91,4);
TASK_PP(16'h1CC92,4);
TASK_PP(16'h1CC93,4);
TASK_PP(16'h1CC94,4);
TASK_PP(16'h1CC95,4);
TASK_PP(16'h1CC96,4);
TASK_PP(16'h1CC97,4);
TASK_PP(16'h1CC98,4);
TASK_PP(16'h1CC99,4);
TASK_PP(16'h1CC9A,4);
TASK_PP(16'h1CC9B,4);
TASK_PP(16'h1CC9C,4);
TASK_PP(16'h1CC9D,4);
TASK_PP(16'h1CC9E,4);
TASK_PP(16'h1CC9F,4);
TASK_PP(16'h1CCA0,4);
TASK_PP(16'h1CCA1,4);
TASK_PP(16'h1CCA2,4);
TASK_PP(16'h1CCA3,4);
TASK_PP(16'h1CCA4,4);
TASK_PP(16'h1CCA5,4);
TASK_PP(16'h1CCA6,4);
TASK_PP(16'h1CCA7,4);
TASK_PP(16'h1CCA8,4);
TASK_PP(16'h1CCA9,4);
TASK_PP(16'h1CCAA,4);
TASK_PP(16'h1CCAB,4);
TASK_PP(16'h1CCAC,4);
TASK_PP(16'h1CCAD,4);
TASK_PP(16'h1CCAE,4);
TASK_PP(16'h1CCAF,4);
TASK_PP(16'h1CCB0,4);
TASK_PP(16'h1CCB1,4);
TASK_PP(16'h1CCB2,4);
TASK_PP(16'h1CCB3,4);
TASK_PP(16'h1CCB4,4);
TASK_PP(16'h1CCB5,4);
TASK_PP(16'h1CCB6,4);
TASK_PP(16'h1CCB7,4);
TASK_PP(16'h1CCB8,4);
TASK_PP(16'h1CCB9,4);
TASK_PP(16'h1CCBA,4);
TASK_PP(16'h1CCBB,4);
TASK_PP(16'h1CCBC,4);
TASK_PP(16'h1CCBD,4);
TASK_PP(16'h1CCBE,4);
TASK_PP(16'h1CCBF,4);
TASK_PP(16'h1CCC0,4);
TASK_PP(16'h1CCC1,4);
TASK_PP(16'h1CCC2,4);
TASK_PP(16'h1CCC3,4);
TASK_PP(16'h1CCC4,4);
TASK_PP(16'h1CCC5,4);
TASK_PP(16'h1CCC6,4);
TASK_PP(16'h1CCC7,4);
TASK_PP(16'h1CCC8,4);
TASK_PP(16'h1CCC9,4);
TASK_PP(16'h1CCCA,4);
TASK_PP(16'h1CCCB,4);
TASK_PP(16'h1CCCC,4);
TASK_PP(16'h1CCCD,4);
TASK_PP(16'h1CCCE,4);
TASK_PP(16'h1CCCF,4);
TASK_PP(16'h1CCD0,4);
TASK_PP(16'h1CCD1,4);
TASK_PP(16'h1CCD2,4);
TASK_PP(16'h1CCD3,4);
TASK_PP(16'h1CCD4,4);
TASK_PP(16'h1CCD5,4);
TASK_PP(16'h1CCD6,4);
TASK_PP(16'h1CCD7,4);
TASK_PP(16'h1CCD8,4);
TASK_PP(16'h1CCD9,4);
TASK_PP(16'h1CCDA,4);
TASK_PP(16'h1CCDB,4);
TASK_PP(16'h1CCDC,4);
TASK_PP(16'h1CCDD,4);
TASK_PP(16'h1CCDE,4);
TASK_PP(16'h1CCDF,4);
TASK_PP(16'h1CCE0,4);
TASK_PP(16'h1CCE1,4);
TASK_PP(16'h1CCE2,4);
TASK_PP(16'h1CCE3,4);
TASK_PP(16'h1CCE4,4);
TASK_PP(16'h1CCE5,4);
TASK_PP(16'h1CCE6,4);
TASK_PP(16'h1CCE7,4);
TASK_PP(16'h1CCE8,4);
TASK_PP(16'h1CCE9,4);
TASK_PP(16'h1CCEA,4);
TASK_PP(16'h1CCEB,4);
TASK_PP(16'h1CCEC,4);
TASK_PP(16'h1CCED,4);
TASK_PP(16'h1CCEE,4);
TASK_PP(16'h1CCEF,4);
TASK_PP(16'h1CCF0,4);
TASK_PP(16'h1CCF1,4);
TASK_PP(16'h1CCF2,4);
TASK_PP(16'h1CCF3,4);
TASK_PP(16'h1CCF4,4);
TASK_PP(16'h1CCF5,4);
TASK_PP(16'h1CCF6,4);
TASK_PP(16'h1CCF7,4);
TASK_PP(16'h1CCF8,4);
TASK_PP(16'h1CCF9,4);
TASK_PP(16'h1CCFA,4);
TASK_PP(16'h1CCFB,4);
TASK_PP(16'h1CCFC,4);
TASK_PP(16'h1CCFD,4);
TASK_PP(16'h1CCFE,4);
TASK_PP(16'h1CCFF,4);
TASK_PP(16'h1CD00,4);
TASK_PP(16'h1CD01,4);
TASK_PP(16'h1CD02,4);
TASK_PP(16'h1CD03,4);
TASK_PP(16'h1CD04,4);
TASK_PP(16'h1CD05,4);
TASK_PP(16'h1CD06,4);
TASK_PP(16'h1CD07,4);
TASK_PP(16'h1CD08,4);
TASK_PP(16'h1CD09,4);
TASK_PP(16'h1CD0A,4);
TASK_PP(16'h1CD0B,4);
TASK_PP(16'h1CD0C,4);
TASK_PP(16'h1CD0D,4);
TASK_PP(16'h1CD0E,4);
TASK_PP(16'h1CD0F,4);
TASK_PP(16'h1CD10,4);
TASK_PP(16'h1CD11,4);
TASK_PP(16'h1CD12,4);
TASK_PP(16'h1CD13,4);
TASK_PP(16'h1CD14,4);
TASK_PP(16'h1CD15,4);
TASK_PP(16'h1CD16,4);
TASK_PP(16'h1CD17,4);
TASK_PP(16'h1CD18,4);
TASK_PP(16'h1CD19,4);
TASK_PP(16'h1CD1A,4);
TASK_PP(16'h1CD1B,4);
TASK_PP(16'h1CD1C,4);
TASK_PP(16'h1CD1D,4);
TASK_PP(16'h1CD1E,4);
TASK_PP(16'h1CD1F,4);
TASK_PP(16'h1CD20,4);
TASK_PP(16'h1CD21,4);
TASK_PP(16'h1CD22,4);
TASK_PP(16'h1CD23,4);
TASK_PP(16'h1CD24,4);
TASK_PP(16'h1CD25,4);
TASK_PP(16'h1CD26,4);
TASK_PP(16'h1CD27,4);
TASK_PP(16'h1CD28,4);
TASK_PP(16'h1CD29,4);
TASK_PP(16'h1CD2A,4);
TASK_PP(16'h1CD2B,4);
TASK_PP(16'h1CD2C,4);
TASK_PP(16'h1CD2D,4);
TASK_PP(16'h1CD2E,4);
TASK_PP(16'h1CD2F,4);
TASK_PP(16'h1CD30,4);
TASK_PP(16'h1CD31,4);
TASK_PP(16'h1CD32,4);
TASK_PP(16'h1CD33,4);
TASK_PP(16'h1CD34,4);
TASK_PP(16'h1CD35,4);
TASK_PP(16'h1CD36,4);
TASK_PP(16'h1CD37,4);
TASK_PP(16'h1CD38,4);
TASK_PP(16'h1CD39,4);
TASK_PP(16'h1CD3A,4);
TASK_PP(16'h1CD3B,4);
TASK_PP(16'h1CD3C,4);
TASK_PP(16'h1CD3D,4);
TASK_PP(16'h1CD3E,4);
TASK_PP(16'h1CD3F,4);
TASK_PP(16'h1CD40,4);
TASK_PP(16'h1CD41,4);
TASK_PP(16'h1CD42,4);
TASK_PP(16'h1CD43,4);
TASK_PP(16'h1CD44,4);
TASK_PP(16'h1CD45,4);
TASK_PP(16'h1CD46,4);
TASK_PP(16'h1CD47,4);
TASK_PP(16'h1CD48,4);
TASK_PP(16'h1CD49,4);
TASK_PP(16'h1CD4A,4);
TASK_PP(16'h1CD4B,4);
TASK_PP(16'h1CD4C,4);
TASK_PP(16'h1CD4D,4);
TASK_PP(16'h1CD4E,4);
TASK_PP(16'h1CD4F,4);
TASK_PP(16'h1CD50,4);
TASK_PP(16'h1CD51,4);
TASK_PP(16'h1CD52,4);
TASK_PP(16'h1CD53,4);
TASK_PP(16'h1CD54,4);
TASK_PP(16'h1CD55,4);
TASK_PP(16'h1CD56,4);
TASK_PP(16'h1CD57,4);
TASK_PP(16'h1CD58,4);
TASK_PP(16'h1CD59,4);
TASK_PP(16'h1CD5A,4);
TASK_PP(16'h1CD5B,4);
TASK_PP(16'h1CD5C,4);
TASK_PP(16'h1CD5D,4);
TASK_PP(16'h1CD5E,4);
TASK_PP(16'h1CD5F,4);
TASK_PP(16'h1CD60,4);
TASK_PP(16'h1CD61,4);
TASK_PP(16'h1CD62,4);
TASK_PP(16'h1CD63,4);
TASK_PP(16'h1CD64,4);
TASK_PP(16'h1CD65,4);
TASK_PP(16'h1CD66,4);
TASK_PP(16'h1CD67,4);
TASK_PP(16'h1CD68,4);
TASK_PP(16'h1CD69,4);
TASK_PP(16'h1CD6A,4);
TASK_PP(16'h1CD6B,4);
TASK_PP(16'h1CD6C,4);
TASK_PP(16'h1CD6D,4);
TASK_PP(16'h1CD6E,4);
TASK_PP(16'h1CD6F,4);
TASK_PP(16'h1CD70,4);
TASK_PP(16'h1CD71,4);
TASK_PP(16'h1CD72,4);
TASK_PP(16'h1CD73,4);
TASK_PP(16'h1CD74,4);
TASK_PP(16'h1CD75,4);
TASK_PP(16'h1CD76,4);
TASK_PP(16'h1CD77,4);
TASK_PP(16'h1CD78,4);
TASK_PP(16'h1CD79,4);
TASK_PP(16'h1CD7A,4);
TASK_PP(16'h1CD7B,4);
TASK_PP(16'h1CD7C,4);
TASK_PP(16'h1CD7D,4);
TASK_PP(16'h1CD7E,4);
TASK_PP(16'h1CD7F,4);
TASK_PP(16'h1CD80,4);
TASK_PP(16'h1CD81,4);
TASK_PP(16'h1CD82,4);
TASK_PP(16'h1CD83,4);
TASK_PP(16'h1CD84,4);
TASK_PP(16'h1CD85,4);
TASK_PP(16'h1CD86,4);
TASK_PP(16'h1CD87,4);
TASK_PP(16'h1CD88,4);
TASK_PP(16'h1CD89,4);
TASK_PP(16'h1CD8A,4);
TASK_PP(16'h1CD8B,4);
TASK_PP(16'h1CD8C,4);
TASK_PP(16'h1CD8D,4);
TASK_PP(16'h1CD8E,4);
TASK_PP(16'h1CD8F,4);
TASK_PP(16'h1CD90,4);
TASK_PP(16'h1CD91,4);
TASK_PP(16'h1CD92,4);
TASK_PP(16'h1CD93,4);
TASK_PP(16'h1CD94,4);
TASK_PP(16'h1CD95,4);
TASK_PP(16'h1CD96,4);
TASK_PP(16'h1CD97,4);
TASK_PP(16'h1CD98,4);
TASK_PP(16'h1CD99,4);
TASK_PP(16'h1CD9A,4);
TASK_PP(16'h1CD9B,4);
TASK_PP(16'h1CD9C,4);
TASK_PP(16'h1CD9D,4);
TASK_PP(16'h1CD9E,4);
TASK_PP(16'h1CD9F,4);
TASK_PP(16'h1CDA0,4);
TASK_PP(16'h1CDA1,4);
TASK_PP(16'h1CDA2,4);
TASK_PP(16'h1CDA3,4);
TASK_PP(16'h1CDA4,4);
TASK_PP(16'h1CDA5,4);
TASK_PP(16'h1CDA6,4);
TASK_PP(16'h1CDA7,4);
TASK_PP(16'h1CDA8,4);
TASK_PP(16'h1CDA9,4);
TASK_PP(16'h1CDAA,4);
TASK_PP(16'h1CDAB,4);
TASK_PP(16'h1CDAC,4);
TASK_PP(16'h1CDAD,4);
TASK_PP(16'h1CDAE,4);
TASK_PP(16'h1CDAF,4);
TASK_PP(16'h1CDB0,4);
TASK_PP(16'h1CDB1,4);
TASK_PP(16'h1CDB2,4);
TASK_PP(16'h1CDB3,4);
TASK_PP(16'h1CDB4,4);
TASK_PP(16'h1CDB5,4);
TASK_PP(16'h1CDB6,4);
TASK_PP(16'h1CDB7,4);
TASK_PP(16'h1CDB8,4);
TASK_PP(16'h1CDB9,4);
TASK_PP(16'h1CDBA,4);
TASK_PP(16'h1CDBB,4);
TASK_PP(16'h1CDBC,4);
TASK_PP(16'h1CDBD,4);
TASK_PP(16'h1CDBE,4);
TASK_PP(16'h1CDBF,4);
TASK_PP(16'h1CDC0,4);
TASK_PP(16'h1CDC1,4);
TASK_PP(16'h1CDC2,4);
TASK_PP(16'h1CDC3,4);
TASK_PP(16'h1CDC4,4);
TASK_PP(16'h1CDC5,4);
TASK_PP(16'h1CDC6,4);
TASK_PP(16'h1CDC7,4);
TASK_PP(16'h1CDC8,4);
TASK_PP(16'h1CDC9,4);
TASK_PP(16'h1CDCA,4);
TASK_PP(16'h1CDCB,4);
TASK_PP(16'h1CDCC,4);
TASK_PP(16'h1CDCD,4);
TASK_PP(16'h1CDCE,4);
TASK_PP(16'h1CDCF,4);
TASK_PP(16'h1CDD0,4);
TASK_PP(16'h1CDD1,4);
TASK_PP(16'h1CDD2,4);
TASK_PP(16'h1CDD3,4);
TASK_PP(16'h1CDD4,4);
TASK_PP(16'h1CDD5,4);
TASK_PP(16'h1CDD6,4);
TASK_PP(16'h1CDD7,4);
TASK_PP(16'h1CDD8,4);
TASK_PP(16'h1CDD9,4);
TASK_PP(16'h1CDDA,4);
TASK_PP(16'h1CDDB,4);
TASK_PP(16'h1CDDC,4);
TASK_PP(16'h1CDDD,4);
TASK_PP(16'h1CDDE,4);
TASK_PP(16'h1CDDF,4);
TASK_PP(16'h1CDE0,4);
TASK_PP(16'h1CDE1,4);
TASK_PP(16'h1CDE2,4);
TASK_PP(16'h1CDE3,4);
TASK_PP(16'h1CDE4,4);
TASK_PP(16'h1CDE5,4);
TASK_PP(16'h1CDE6,4);
TASK_PP(16'h1CDE7,4);
TASK_PP(16'h1CDE8,4);
TASK_PP(16'h1CDE9,4);
TASK_PP(16'h1CDEA,4);
TASK_PP(16'h1CDEB,4);
TASK_PP(16'h1CDEC,4);
TASK_PP(16'h1CDED,4);
TASK_PP(16'h1CDEE,4);
TASK_PP(16'h1CDEF,4);
TASK_PP(16'h1CDF0,4);
TASK_PP(16'h1CDF1,4);
TASK_PP(16'h1CDF2,4);
TASK_PP(16'h1CDF3,4);
TASK_PP(16'h1CDF4,4);
TASK_PP(16'h1CDF5,4);
TASK_PP(16'h1CDF6,4);
TASK_PP(16'h1CDF7,4);
TASK_PP(16'h1CDF8,4);
TASK_PP(16'h1CDF9,4);
TASK_PP(16'h1CDFA,4);
TASK_PP(16'h1CDFB,4);
TASK_PP(16'h1CDFC,4);
TASK_PP(16'h1CDFD,4);
TASK_PP(16'h1CDFE,4);
TASK_PP(16'h1CDFF,4);
TASK_PP(16'h1CE00,4);
TASK_PP(16'h1CE01,4);
TASK_PP(16'h1CE02,4);
TASK_PP(16'h1CE03,4);
TASK_PP(16'h1CE04,4);
TASK_PP(16'h1CE05,4);
TASK_PP(16'h1CE06,4);
TASK_PP(16'h1CE07,4);
TASK_PP(16'h1CE08,4);
TASK_PP(16'h1CE09,4);
TASK_PP(16'h1CE0A,4);
TASK_PP(16'h1CE0B,4);
TASK_PP(16'h1CE0C,4);
TASK_PP(16'h1CE0D,4);
TASK_PP(16'h1CE0E,4);
TASK_PP(16'h1CE0F,4);
TASK_PP(16'h1CE10,4);
TASK_PP(16'h1CE11,4);
TASK_PP(16'h1CE12,4);
TASK_PP(16'h1CE13,4);
TASK_PP(16'h1CE14,4);
TASK_PP(16'h1CE15,4);
TASK_PP(16'h1CE16,4);
TASK_PP(16'h1CE17,4);
TASK_PP(16'h1CE18,4);
TASK_PP(16'h1CE19,4);
TASK_PP(16'h1CE1A,4);
TASK_PP(16'h1CE1B,4);
TASK_PP(16'h1CE1C,4);
TASK_PP(16'h1CE1D,4);
TASK_PP(16'h1CE1E,4);
TASK_PP(16'h1CE1F,4);
TASK_PP(16'h1CE20,4);
TASK_PP(16'h1CE21,4);
TASK_PP(16'h1CE22,4);
TASK_PP(16'h1CE23,4);
TASK_PP(16'h1CE24,4);
TASK_PP(16'h1CE25,4);
TASK_PP(16'h1CE26,4);
TASK_PP(16'h1CE27,4);
TASK_PP(16'h1CE28,4);
TASK_PP(16'h1CE29,4);
TASK_PP(16'h1CE2A,4);
TASK_PP(16'h1CE2B,4);
TASK_PP(16'h1CE2C,4);
TASK_PP(16'h1CE2D,4);
TASK_PP(16'h1CE2E,4);
TASK_PP(16'h1CE2F,4);
TASK_PP(16'h1CE30,4);
TASK_PP(16'h1CE31,4);
TASK_PP(16'h1CE32,4);
TASK_PP(16'h1CE33,4);
TASK_PP(16'h1CE34,4);
TASK_PP(16'h1CE35,4);
TASK_PP(16'h1CE36,4);
TASK_PP(16'h1CE37,4);
TASK_PP(16'h1CE38,4);
TASK_PP(16'h1CE39,4);
TASK_PP(16'h1CE3A,4);
TASK_PP(16'h1CE3B,4);
TASK_PP(16'h1CE3C,4);
TASK_PP(16'h1CE3D,4);
TASK_PP(16'h1CE3E,4);
TASK_PP(16'h1CE3F,4);
TASK_PP(16'h1CE40,4);
TASK_PP(16'h1CE41,4);
TASK_PP(16'h1CE42,4);
TASK_PP(16'h1CE43,4);
TASK_PP(16'h1CE44,4);
TASK_PP(16'h1CE45,4);
TASK_PP(16'h1CE46,4);
TASK_PP(16'h1CE47,4);
TASK_PP(16'h1CE48,4);
TASK_PP(16'h1CE49,4);
TASK_PP(16'h1CE4A,4);
TASK_PP(16'h1CE4B,4);
TASK_PP(16'h1CE4C,4);
TASK_PP(16'h1CE4D,4);
TASK_PP(16'h1CE4E,4);
TASK_PP(16'h1CE4F,4);
TASK_PP(16'h1CE50,4);
TASK_PP(16'h1CE51,4);
TASK_PP(16'h1CE52,4);
TASK_PP(16'h1CE53,4);
TASK_PP(16'h1CE54,4);
TASK_PP(16'h1CE55,4);
TASK_PP(16'h1CE56,4);
TASK_PP(16'h1CE57,4);
TASK_PP(16'h1CE58,4);
TASK_PP(16'h1CE59,4);
TASK_PP(16'h1CE5A,4);
TASK_PP(16'h1CE5B,4);
TASK_PP(16'h1CE5C,4);
TASK_PP(16'h1CE5D,4);
TASK_PP(16'h1CE5E,4);
TASK_PP(16'h1CE5F,4);
TASK_PP(16'h1CE60,4);
TASK_PP(16'h1CE61,4);
TASK_PP(16'h1CE62,4);
TASK_PP(16'h1CE63,4);
TASK_PP(16'h1CE64,4);
TASK_PP(16'h1CE65,4);
TASK_PP(16'h1CE66,4);
TASK_PP(16'h1CE67,4);
TASK_PP(16'h1CE68,4);
TASK_PP(16'h1CE69,4);
TASK_PP(16'h1CE6A,4);
TASK_PP(16'h1CE6B,4);
TASK_PP(16'h1CE6C,4);
TASK_PP(16'h1CE6D,4);
TASK_PP(16'h1CE6E,4);
TASK_PP(16'h1CE6F,4);
TASK_PP(16'h1CE70,4);
TASK_PP(16'h1CE71,4);
TASK_PP(16'h1CE72,4);
TASK_PP(16'h1CE73,4);
TASK_PP(16'h1CE74,4);
TASK_PP(16'h1CE75,4);
TASK_PP(16'h1CE76,4);
TASK_PP(16'h1CE77,4);
TASK_PP(16'h1CE78,4);
TASK_PP(16'h1CE79,4);
TASK_PP(16'h1CE7A,4);
TASK_PP(16'h1CE7B,4);
TASK_PP(16'h1CE7C,4);
TASK_PP(16'h1CE7D,4);
TASK_PP(16'h1CE7E,4);
TASK_PP(16'h1CE7F,4);
TASK_PP(16'h1CE80,4);
TASK_PP(16'h1CE81,4);
TASK_PP(16'h1CE82,4);
TASK_PP(16'h1CE83,4);
TASK_PP(16'h1CE84,4);
TASK_PP(16'h1CE85,4);
TASK_PP(16'h1CE86,4);
TASK_PP(16'h1CE87,4);
TASK_PP(16'h1CE88,4);
TASK_PP(16'h1CE89,4);
TASK_PP(16'h1CE8A,4);
TASK_PP(16'h1CE8B,4);
TASK_PP(16'h1CE8C,4);
TASK_PP(16'h1CE8D,4);
TASK_PP(16'h1CE8E,4);
TASK_PP(16'h1CE8F,4);
TASK_PP(16'h1CE90,4);
TASK_PP(16'h1CE91,4);
TASK_PP(16'h1CE92,4);
TASK_PP(16'h1CE93,4);
TASK_PP(16'h1CE94,4);
TASK_PP(16'h1CE95,4);
TASK_PP(16'h1CE96,4);
TASK_PP(16'h1CE97,4);
TASK_PP(16'h1CE98,4);
TASK_PP(16'h1CE99,4);
TASK_PP(16'h1CE9A,4);
TASK_PP(16'h1CE9B,4);
TASK_PP(16'h1CE9C,4);
TASK_PP(16'h1CE9D,4);
TASK_PP(16'h1CE9E,4);
TASK_PP(16'h1CE9F,4);
TASK_PP(16'h1CEA0,4);
TASK_PP(16'h1CEA1,4);
TASK_PP(16'h1CEA2,4);
TASK_PP(16'h1CEA3,4);
TASK_PP(16'h1CEA4,4);
TASK_PP(16'h1CEA5,4);
TASK_PP(16'h1CEA6,4);
TASK_PP(16'h1CEA7,4);
TASK_PP(16'h1CEA8,4);
TASK_PP(16'h1CEA9,4);
TASK_PP(16'h1CEAA,4);
TASK_PP(16'h1CEAB,4);
TASK_PP(16'h1CEAC,4);
TASK_PP(16'h1CEAD,4);
TASK_PP(16'h1CEAE,4);
TASK_PP(16'h1CEAF,4);
TASK_PP(16'h1CEB0,4);
TASK_PP(16'h1CEB1,4);
TASK_PP(16'h1CEB2,4);
TASK_PP(16'h1CEB3,4);
TASK_PP(16'h1CEB4,4);
TASK_PP(16'h1CEB5,4);
TASK_PP(16'h1CEB6,4);
TASK_PP(16'h1CEB7,4);
TASK_PP(16'h1CEB8,4);
TASK_PP(16'h1CEB9,4);
TASK_PP(16'h1CEBA,4);
TASK_PP(16'h1CEBB,4);
TASK_PP(16'h1CEBC,4);
TASK_PP(16'h1CEBD,4);
TASK_PP(16'h1CEBE,4);
TASK_PP(16'h1CEBF,4);
TASK_PP(16'h1CEC0,4);
TASK_PP(16'h1CEC1,4);
TASK_PP(16'h1CEC2,4);
TASK_PP(16'h1CEC3,4);
TASK_PP(16'h1CEC4,4);
TASK_PP(16'h1CEC5,4);
TASK_PP(16'h1CEC6,4);
TASK_PP(16'h1CEC7,4);
TASK_PP(16'h1CEC8,4);
TASK_PP(16'h1CEC9,4);
TASK_PP(16'h1CECA,4);
TASK_PP(16'h1CECB,4);
TASK_PP(16'h1CECC,4);
TASK_PP(16'h1CECD,4);
TASK_PP(16'h1CECE,4);
TASK_PP(16'h1CECF,4);
TASK_PP(16'h1CED0,4);
TASK_PP(16'h1CED1,4);
TASK_PP(16'h1CED2,4);
TASK_PP(16'h1CED3,4);
TASK_PP(16'h1CED4,4);
TASK_PP(16'h1CED5,4);
TASK_PP(16'h1CED6,4);
TASK_PP(16'h1CED7,4);
TASK_PP(16'h1CED8,4);
TASK_PP(16'h1CED9,4);
TASK_PP(16'h1CEDA,4);
TASK_PP(16'h1CEDB,4);
TASK_PP(16'h1CEDC,4);
TASK_PP(16'h1CEDD,4);
TASK_PP(16'h1CEDE,4);
TASK_PP(16'h1CEDF,4);
TASK_PP(16'h1CEE0,4);
TASK_PP(16'h1CEE1,4);
TASK_PP(16'h1CEE2,4);
TASK_PP(16'h1CEE3,4);
TASK_PP(16'h1CEE4,4);
TASK_PP(16'h1CEE5,4);
TASK_PP(16'h1CEE6,4);
TASK_PP(16'h1CEE7,4);
TASK_PP(16'h1CEE8,4);
TASK_PP(16'h1CEE9,4);
TASK_PP(16'h1CEEA,4);
TASK_PP(16'h1CEEB,4);
TASK_PP(16'h1CEEC,4);
TASK_PP(16'h1CEED,4);
TASK_PP(16'h1CEEE,4);
TASK_PP(16'h1CEEF,4);
TASK_PP(16'h1CEF0,4);
TASK_PP(16'h1CEF1,4);
TASK_PP(16'h1CEF2,4);
TASK_PP(16'h1CEF3,4);
TASK_PP(16'h1CEF4,4);
TASK_PP(16'h1CEF5,4);
TASK_PP(16'h1CEF6,4);
TASK_PP(16'h1CEF7,4);
TASK_PP(16'h1CEF8,4);
TASK_PP(16'h1CEF9,4);
TASK_PP(16'h1CEFA,4);
TASK_PP(16'h1CEFB,4);
TASK_PP(16'h1CEFC,4);
TASK_PP(16'h1CEFD,4);
TASK_PP(16'h1CEFE,4);
TASK_PP(16'h1CEFF,4);
TASK_PP(16'h1CF00,4);
TASK_PP(16'h1CF01,4);
TASK_PP(16'h1CF02,4);
TASK_PP(16'h1CF03,4);
TASK_PP(16'h1CF04,4);
TASK_PP(16'h1CF05,4);
TASK_PP(16'h1CF06,4);
TASK_PP(16'h1CF07,4);
TASK_PP(16'h1CF08,4);
TASK_PP(16'h1CF09,4);
TASK_PP(16'h1CF0A,4);
TASK_PP(16'h1CF0B,4);
TASK_PP(16'h1CF0C,4);
TASK_PP(16'h1CF0D,4);
TASK_PP(16'h1CF0E,4);
TASK_PP(16'h1CF0F,4);
TASK_PP(16'h1CF10,4);
TASK_PP(16'h1CF11,4);
TASK_PP(16'h1CF12,4);
TASK_PP(16'h1CF13,4);
TASK_PP(16'h1CF14,4);
TASK_PP(16'h1CF15,4);
TASK_PP(16'h1CF16,4);
TASK_PP(16'h1CF17,4);
TASK_PP(16'h1CF18,4);
TASK_PP(16'h1CF19,4);
TASK_PP(16'h1CF1A,4);
TASK_PP(16'h1CF1B,4);
TASK_PP(16'h1CF1C,4);
TASK_PP(16'h1CF1D,4);
TASK_PP(16'h1CF1E,4);
TASK_PP(16'h1CF1F,4);
TASK_PP(16'h1CF20,4);
TASK_PP(16'h1CF21,4);
TASK_PP(16'h1CF22,4);
TASK_PP(16'h1CF23,4);
TASK_PP(16'h1CF24,4);
TASK_PP(16'h1CF25,4);
TASK_PP(16'h1CF26,4);
TASK_PP(16'h1CF27,4);
TASK_PP(16'h1CF28,4);
TASK_PP(16'h1CF29,4);
TASK_PP(16'h1CF2A,4);
TASK_PP(16'h1CF2B,4);
TASK_PP(16'h1CF2C,4);
TASK_PP(16'h1CF2D,4);
TASK_PP(16'h1CF2E,4);
TASK_PP(16'h1CF2F,4);
TASK_PP(16'h1CF30,4);
TASK_PP(16'h1CF31,4);
TASK_PP(16'h1CF32,4);
TASK_PP(16'h1CF33,4);
TASK_PP(16'h1CF34,4);
TASK_PP(16'h1CF35,4);
TASK_PP(16'h1CF36,4);
TASK_PP(16'h1CF37,4);
TASK_PP(16'h1CF38,4);
TASK_PP(16'h1CF39,4);
TASK_PP(16'h1CF3A,4);
TASK_PP(16'h1CF3B,4);
TASK_PP(16'h1CF3C,4);
TASK_PP(16'h1CF3D,4);
TASK_PP(16'h1CF3E,4);
TASK_PP(16'h1CF3F,4);
TASK_PP(16'h1CF40,4);
TASK_PP(16'h1CF41,4);
TASK_PP(16'h1CF42,4);
TASK_PP(16'h1CF43,4);
TASK_PP(16'h1CF44,4);
TASK_PP(16'h1CF45,4);
TASK_PP(16'h1CF46,4);
TASK_PP(16'h1CF47,4);
TASK_PP(16'h1CF48,4);
TASK_PP(16'h1CF49,4);
TASK_PP(16'h1CF4A,4);
TASK_PP(16'h1CF4B,4);
TASK_PP(16'h1CF4C,4);
TASK_PP(16'h1CF4D,4);
TASK_PP(16'h1CF4E,4);
TASK_PP(16'h1CF4F,4);
TASK_PP(16'h1CF50,4);
TASK_PP(16'h1CF51,4);
TASK_PP(16'h1CF52,4);
TASK_PP(16'h1CF53,4);
TASK_PP(16'h1CF54,4);
TASK_PP(16'h1CF55,4);
TASK_PP(16'h1CF56,4);
TASK_PP(16'h1CF57,4);
TASK_PP(16'h1CF58,4);
TASK_PP(16'h1CF59,4);
TASK_PP(16'h1CF5A,4);
TASK_PP(16'h1CF5B,4);
TASK_PP(16'h1CF5C,4);
TASK_PP(16'h1CF5D,4);
TASK_PP(16'h1CF5E,4);
TASK_PP(16'h1CF5F,4);
TASK_PP(16'h1CF60,4);
TASK_PP(16'h1CF61,4);
TASK_PP(16'h1CF62,4);
TASK_PP(16'h1CF63,4);
TASK_PP(16'h1CF64,4);
TASK_PP(16'h1CF65,4);
TASK_PP(16'h1CF66,4);
TASK_PP(16'h1CF67,4);
TASK_PP(16'h1CF68,4);
TASK_PP(16'h1CF69,4);
TASK_PP(16'h1CF6A,4);
TASK_PP(16'h1CF6B,4);
TASK_PP(16'h1CF6C,4);
TASK_PP(16'h1CF6D,4);
TASK_PP(16'h1CF6E,4);
TASK_PP(16'h1CF6F,4);
TASK_PP(16'h1CF70,4);
TASK_PP(16'h1CF71,4);
TASK_PP(16'h1CF72,4);
TASK_PP(16'h1CF73,4);
TASK_PP(16'h1CF74,4);
TASK_PP(16'h1CF75,4);
TASK_PP(16'h1CF76,4);
TASK_PP(16'h1CF77,4);
TASK_PP(16'h1CF78,4);
TASK_PP(16'h1CF79,4);
TASK_PP(16'h1CF7A,4);
TASK_PP(16'h1CF7B,4);
TASK_PP(16'h1CF7C,4);
TASK_PP(16'h1CF7D,4);
TASK_PP(16'h1CF7E,4);
TASK_PP(16'h1CF7F,4);
TASK_PP(16'h1CF80,4);
TASK_PP(16'h1CF81,4);
TASK_PP(16'h1CF82,4);
TASK_PP(16'h1CF83,4);
TASK_PP(16'h1CF84,4);
TASK_PP(16'h1CF85,4);
TASK_PP(16'h1CF86,4);
TASK_PP(16'h1CF87,4);
TASK_PP(16'h1CF88,4);
TASK_PP(16'h1CF89,4);
TASK_PP(16'h1CF8A,4);
TASK_PP(16'h1CF8B,4);
TASK_PP(16'h1CF8C,4);
TASK_PP(16'h1CF8D,4);
TASK_PP(16'h1CF8E,4);
TASK_PP(16'h1CF8F,4);
TASK_PP(16'h1CF90,4);
TASK_PP(16'h1CF91,4);
TASK_PP(16'h1CF92,4);
TASK_PP(16'h1CF93,4);
TASK_PP(16'h1CF94,4);
TASK_PP(16'h1CF95,4);
TASK_PP(16'h1CF96,4);
TASK_PP(16'h1CF97,4);
TASK_PP(16'h1CF98,4);
TASK_PP(16'h1CF99,4);
TASK_PP(16'h1CF9A,4);
TASK_PP(16'h1CF9B,4);
TASK_PP(16'h1CF9C,4);
TASK_PP(16'h1CF9D,4);
TASK_PP(16'h1CF9E,4);
TASK_PP(16'h1CF9F,4);
TASK_PP(16'h1CFA0,4);
TASK_PP(16'h1CFA1,4);
TASK_PP(16'h1CFA2,4);
TASK_PP(16'h1CFA3,4);
TASK_PP(16'h1CFA4,4);
TASK_PP(16'h1CFA5,4);
TASK_PP(16'h1CFA6,4);
TASK_PP(16'h1CFA7,4);
TASK_PP(16'h1CFA8,4);
TASK_PP(16'h1CFA9,4);
TASK_PP(16'h1CFAA,4);
TASK_PP(16'h1CFAB,4);
TASK_PP(16'h1CFAC,4);
TASK_PP(16'h1CFAD,4);
TASK_PP(16'h1CFAE,4);
TASK_PP(16'h1CFAF,4);
TASK_PP(16'h1CFB0,4);
TASK_PP(16'h1CFB1,4);
TASK_PP(16'h1CFB2,4);
TASK_PP(16'h1CFB3,4);
TASK_PP(16'h1CFB4,4);
TASK_PP(16'h1CFB5,4);
TASK_PP(16'h1CFB6,4);
TASK_PP(16'h1CFB7,4);
TASK_PP(16'h1CFB8,4);
TASK_PP(16'h1CFB9,4);
TASK_PP(16'h1CFBA,4);
TASK_PP(16'h1CFBB,4);
TASK_PP(16'h1CFBC,4);
TASK_PP(16'h1CFBD,4);
TASK_PP(16'h1CFBE,4);
TASK_PP(16'h1CFBF,4);
TASK_PP(16'h1CFC0,4);
TASK_PP(16'h1CFC1,4);
TASK_PP(16'h1CFC2,4);
TASK_PP(16'h1CFC3,4);
TASK_PP(16'h1CFC4,4);
TASK_PP(16'h1CFC5,4);
TASK_PP(16'h1CFC6,4);
TASK_PP(16'h1CFC7,4);
TASK_PP(16'h1CFC8,4);
TASK_PP(16'h1CFC9,4);
TASK_PP(16'h1CFCA,4);
TASK_PP(16'h1CFCB,4);
TASK_PP(16'h1CFCC,4);
TASK_PP(16'h1CFCD,4);
TASK_PP(16'h1CFCE,4);
TASK_PP(16'h1CFCF,4);
TASK_PP(16'h1CFD0,4);
TASK_PP(16'h1CFD1,4);
TASK_PP(16'h1CFD2,4);
TASK_PP(16'h1CFD3,4);
TASK_PP(16'h1CFD4,4);
TASK_PP(16'h1CFD5,4);
TASK_PP(16'h1CFD6,4);
TASK_PP(16'h1CFD7,4);
TASK_PP(16'h1CFD8,4);
TASK_PP(16'h1CFD9,4);
TASK_PP(16'h1CFDA,4);
TASK_PP(16'h1CFDB,4);
TASK_PP(16'h1CFDC,4);
TASK_PP(16'h1CFDD,4);
TASK_PP(16'h1CFDE,4);
TASK_PP(16'h1CFDF,4);
TASK_PP(16'h1CFE0,4);
TASK_PP(16'h1CFE1,4);
TASK_PP(16'h1CFE2,4);
TASK_PP(16'h1CFE3,4);
TASK_PP(16'h1CFE4,4);
TASK_PP(16'h1CFE5,4);
TASK_PP(16'h1CFE6,4);
TASK_PP(16'h1CFE7,4);
TASK_PP(16'h1CFE8,4);
TASK_PP(16'h1CFE9,4);
TASK_PP(16'h1CFEA,4);
TASK_PP(16'h1CFEB,4);
TASK_PP(16'h1CFEC,4);
TASK_PP(16'h1CFED,4);
TASK_PP(16'h1CFEE,4);
TASK_PP(16'h1CFEF,4);
TASK_PP(16'h1CFF0,4);
TASK_PP(16'h1CFF1,4);
TASK_PP(16'h1CFF2,4);
TASK_PP(16'h1CFF3,4);
TASK_PP(16'h1CFF4,4);
TASK_PP(16'h1CFF5,4);
TASK_PP(16'h1CFF6,4);
TASK_PP(16'h1CFF7,4);
TASK_PP(16'h1CFF8,4);
TASK_PP(16'h1CFF9,4);
TASK_PP(16'h1CFFA,4);
TASK_PP(16'h1CFFB,4);
TASK_PP(16'h1CFFC,4);
TASK_PP(16'h1CFFD,4);
TASK_PP(16'h1CFFE,4);
TASK_PP(16'h1CFFF,4);
TASK_PP(16'h1D000,4);
TASK_PP(16'h1D001,4);
TASK_PP(16'h1D002,4);
TASK_PP(16'h1D003,4);
TASK_PP(16'h1D004,4);
TASK_PP(16'h1D005,4);
TASK_PP(16'h1D006,4);
TASK_PP(16'h1D007,4);
TASK_PP(16'h1D008,4);
TASK_PP(16'h1D009,4);
TASK_PP(16'h1D00A,4);
TASK_PP(16'h1D00B,4);
TASK_PP(16'h1D00C,4);
TASK_PP(16'h1D00D,4);
TASK_PP(16'h1D00E,4);
TASK_PP(16'h1D00F,4);
TASK_PP(16'h1D010,4);
TASK_PP(16'h1D011,4);
TASK_PP(16'h1D012,4);
TASK_PP(16'h1D013,4);
TASK_PP(16'h1D014,4);
TASK_PP(16'h1D015,4);
TASK_PP(16'h1D016,4);
TASK_PP(16'h1D017,4);
TASK_PP(16'h1D018,4);
TASK_PP(16'h1D019,4);
TASK_PP(16'h1D01A,4);
TASK_PP(16'h1D01B,4);
TASK_PP(16'h1D01C,4);
TASK_PP(16'h1D01D,4);
TASK_PP(16'h1D01E,4);
TASK_PP(16'h1D01F,4);
TASK_PP(16'h1D020,4);
TASK_PP(16'h1D021,4);
TASK_PP(16'h1D022,4);
TASK_PP(16'h1D023,4);
TASK_PP(16'h1D024,4);
TASK_PP(16'h1D025,4);
TASK_PP(16'h1D026,4);
TASK_PP(16'h1D027,4);
TASK_PP(16'h1D028,4);
TASK_PP(16'h1D029,4);
TASK_PP(16'h1D02A,4);
TASK_PP(16'h1D02B,4);
TASK_PP(16'h1D02C,4);
TASK_PP(16'h1D02D,4);
TASK_PP(16'h1D02E,4);
TASK_PP(16'h1D02F,4);
TASK_PP(16'h1D030,4);
TASK_PP(16'h1D031,4);
TASK_PP(16'h1D032,4);
TASK_PP(16'h1D033,4);
TASK_PP(16'h1D034,4);
TASK_PP(16'h1D035,4);
TASK_PP(16'h1D036,4);
TASK_PP(16'h1D037,4);
TASK_PP(16'h1D038,4);
TASK_PP(16'h1D039,4);
TASK_PP(16'h1D03A,4);
TASK_PP(16'h1D03B,4);
TASK_PP(16'h1D03C,4);
TASK_PP(16'h1D03D,4);
TASK_PP(16'h1D03E,4);
TASK_PP(16'h1D03F,4);
TASK_PP(16'h1D040,4);
TASK_PP(16'h1D041,4);
TASK_PP(16'h1D042,4);
TASK_PP(16'h1D043,4);
TASK_PP(16'h1D044,4);
TASK_PP(16'h1D045,4);
TASK_PP(16'h1D046,4);
TASK_PP(16'h1D047,4);
TASK_PP(16'h1D048,4);
TASK_PP(16'h1D049,4);
TASK_PP(16'h1D04A,4);
TASK_PP(16'h1D04B,4);
TASK_PP(16'h1D04C,4);
TASK_PP(16'h1D04D,4);
TASK_PP(16'h1D04E,4);
TASK_PP(16'h1D04F,4);
TASK_PP(16'h1D050,4);
TASK_PP(16'h1D051,4);
TASK_PP(16'h1D052,4);
TASK_PP(16'h1D053,4);
TASK_PP(16'h1D054,4);
TASK_PP(16'h1D055,4);
TASK_PP(16'h1D056,4);
TASK_PP(16'h1D057,4);
TASK_PP(16'h1D058,4);
TASK_PP(16'h1D059,4);
TASK_PP(16'h1D05A,4);
TASK_PP(16'h1D05B,4);
TASK_PP(16'h1D05C,4);
TASK_PP(16'h1D05D,4);
TASK_PP(16'h1D05E,4);
TASK_PP(16'h1D05F,4);
TASK_PP(16'h1D060,4);
TASK_PP(16'h1D061,4);
TASK_PP(16'h1D062,4);
TASK_PP(16'h1D063,4);
TASK_PP(16'h1D064,4);
TASK_PP(16'h1D065,4);
TASK_PP(16'h1D066,4);
TASK_PP(16'h1D067,4);
TASK_PP(16'h1D068,4);
TASK_PP(16'h1D069,4);
TASK_PP(16'h1D06A,4);
TASK_PP(16'h1D06B,4);
TASK_PP(16'h1D06C,4);
TASK_PP(16'h1D06D,4);
TASK_PP(16'h1D06E,4);
TASK_PP(16'h1D06F,4);
TASK_PP(16'h1D070,4);
TASK_PP(16'h1D071,4);
TASK_PP(16'h1D072,4);
TASK_PP(16'h1D073,4);
TASK_PP(16'h1D074,4);
TASK_PP(16'h1D075,4);
TASK_PP(16'h1D076,4);
TASK_PP(16'h1D077,4);
TASK_PP(16'h1D078,4);
TASK_PP(16'h1D079,4);
TASK_PP(16'h1D07A,4);
TASK_PP(16'h1D07B,4);
TASK_PP(16'h1D07C,4);
TASK_PP(16'h1D07D,4);
TASK_PP(16'h1D07E,4);
TASK_PP(16'h1D07F,4);
TASK_PP(16'h1D080,4);
TASK_PP(16'h1D081,4);
TASK_PP(16'h1D082,4);
TASK_PP(16'h1D083,4);
TASK_PP(16'h1D084,4);
TASK_PP(16'h1D085,4);
TASK_PP(16'h1D086,4);
TASK_PP(16'h1D087,4);
TASK_PP(16'h1D088,4);
TASK_PP(16'h1D089,4);
TASK_PP(16'h1D08A,4);
TASK_PP(16'h1D08B,4);
TASK_PP(16'h1D08C,4);
TASK_PP(16'h1D08D,4);
TASK_PP(16'h1D08E,4);
TASK_PP(16'h1D08F,4);
TASK_PP(16'h1D090,4);
TASK_PP(16'h1D091,4);
TASK_PP(16'h1D092,4);
TASK_PP(16'h1D093,4);
TASK_PP(16'h1D094,4);
TASK_PP(16'h1D095,4);
TASK_PP(16'h1D096,4);
TASK_PP(16'h1D097,4);
TASK_PP(16'h1D098,4);
TASK_PP(16'h1D099,4);
TASK_PP(16'h1D09A,4);
TASK_PP(16'h1D09B,4);
TASK_PP(16'h1D09C,4);
TASK_PP(16'h1D09D,4);
TASK_PP(16'h1D09E,4);
TASK_PP(16'h1D09F,4);
TASK_PP(16'h1D0A0,4);
TASK_PP(16'h1D0A1,4);
TASK_PP(16'h1D0A2,4);
TASK_PP(16'h1D0A3,4);
TASK_PP(16'h1D0A4,4);
TASK_PP(16'h1D0A5,4);
TASK_PP(16'h1D0A6,4);
TASK_PP(16'h1D0A7,4);
TASK_PP(16'h1D0A8,4);
TASK_PP(16'h1D0A9,4);
TASK_PP(16'h1D0AA,4);
TASK_PP(16'h1D0AB,4);
TASK_PP(16'h1D0AC,4);
TASK_PP(16'h1D0AD,4);
TASK_PP(16'h1D0AE,4);
TASK_PP(16'h1D0AF,4);
TASK_PP(16'h1D0B0,4);
TASK_PP(16'h1D0B1,4);
TASK_PP(16'h1D0B2,4);
TASK_PP(16'h1D0B3,4);
TASK_PP(16'h1D0B4,4);
TASK_PP(16'h1D0B5,4);
TASK_PP(16'h1D0B6,4);
TASK_PP(16'h1D0B7,4);
TASK_PP(16'h1D0B8,4);
TASK_PP(16'h1D0B9,4);
TASK_PP(16'h1D0BA,4);
TASK_PP(16'h1D0BB,4);
TASK_PP(16'h1D0BC,4);
TASK_PP(16'h1D0BD,4);
TASK_PP(16'h1D0BE,4);
TASK_PP(16'h1D0BF,4);
TASK_PP(16'h1D0C0,4);
TASK_PP(16'h1D0C1,4);
TASK_PP(16'h1D0C2,4);
TASK_PP(16'h1D0C3,4);
TASK_PP(16'h1D0C4,4);
TASK_PP(16'h1D0C5,4);
TASK_PP(16'h1D0C6,4);
TASK_PP(16'h1D0C7,4);
TASK_PP(16'h1D0C8,4);
TASK_PP(16'h1D0C9,4);
TASK_PP(16'h1D0CA,4);
TASK_PP(16'h1D0CB,4);
TASK_PP(16'h1D0CC,4);
TASK_PP(16'h1D0CD,4);
TASK_PP(16'h1D0CE,4);
TASK_PP(16'h1D0CF,4);
TASK_PP(16'h1D0D0,4);
TASK_PP(16'h1D0D1,4);
TASK_PP(16'h1D0D2,4);
TASK_PP(16'h1D0D3,4);
TASK_PP(16'h1D0D4,4);
TASK_PP(16'h1D0D5,4);
TASK_PP(16'h1D0D6,4);
TASK_PP(16'h1D0D7,4);
TASK_PP(16'h1D0D8,4);
TASK_PP(16'h1D0D9,4);
TASK_PP(16'h1D0DA,4);
TASK_PP(16'h1D0DB,4);
TASK_PP(16'h1D0DC,4);
TASK_PP(16'h1D0DD,4);
TASK_PP(16'h1D0DE,4);
TASK_PP(16'h1D0DF,4);
TASK_PP(16'h1D0E0,4);
TASK_PP(16'h1D0E1,4);
TASK_PP(16'h1D0E2,4);
TASK_PP(16'h1D0E3,4);
TASK_PP(16'h1D0E4,4);
TASK_PP(16'h1D0E5,4);
TASK_PP(16'h1D0E6,4);
TASK_PP(16'h1D0E7,4);
TASK_PP(16'h1D0E8,4);
TASK_PP(16'h1D0E9,4);
TASK_PP(16'h1D0EA,4);
TASK_PP(16'h1D0EB,4);
TASK_PP(16'h1D0EC,4);
TASK_PP(16'h1D0ED,4);
TASK_PP(16'h1D0EE,4);
TASK_PP(16'h1D0EF,4);
TASK_PP(16'h1D0F0,4);
TASK_PP(16'h1D0F1,4);
TASK_PP(16'h1D0F2,4);
TASK_PP(16'h1D0F3,4);
TASK_PP(16'h1D0F4,4);
TASK_PP(16'h1D0F5,4);
TASK_PP(16'h1D0F6,4);
TASK_PP(16'h1D0F7,4);
TASK_PP(16'h1D0F8,4);
TASK_PP(16'h1D0F9,4);
TASK_PP(16'h1D0FA,4);
TASK_PP(16'h1D0FB,4);
TASK_PP(16'h1D0FC,4);
TASK_PP(16'h1D0FD,4);
TASK_PP(16'h1D0FE,4);
TASK_PP(16'h1D0FF,4);
TASK_PP(16'h1D100,4);
TASK_PP(16'h1D101,4);
TASK_PP(16'h1D102,4);
TASK_PP(16'h1D103,4);
TASK_PP(16'h1D104,4);
TASK_PP(16'h1D105,4);
TASK_PP(16'h1D106,4);
TASK_PP(16'h1D107,4);
TASK_PP(16'h1D108,4);
TASK_PP(16'h1D109,4);
TASK_PP(16'h1D10A,4);
TASK_PP(16'h1D10B,4);
TASK_PP(16'h1D10C,4);
TASK_PP(16'h1D10D,4);
TASK_PP(16'h1D10E,4);
TASK_PP(16'h1D10F,4);
TASK_PP(16'h1D110,4);
TASK_PP(16'h1D111,4);
TASK_PP(16'h1D112,4);
TASK_PP(16'h1D113,4);
TASK_PP(16'h1D114,4);
TASK_PP(16'h1D115,4);
TASK_PP(16'h1D116,4);
TASK_PP(16'h1D117,4);
TASK_PP(16'h1D118,4);
TASK_PP(16'h1D119,4);
TASK_PP(16'h1D11A,4);
TASK_PP(16'h1D11B,4);
TASK_PP(16'h1D11C,4);
TASK_PP(16'h1D11D,4);
TASK_PP(16'h1D11E,4);
TASK_PP(16'h1D11F,4);
TASK_PP(16'h1D120,4);
TASK_PP(16'h1D121,4);
TASK_PP(16'h1D122,4);
TASK_PP(16'h1D123,4);
TASK_PP(16'h1D124,4);
TASK_PP(16'h1D125,4);
TASK_PP(16'h1D126,4);
TASK_PP(16'h1D127,4);
TASK_PP(16'h1D128,4);
TASK_PP(16'h1D129,4);
TASK_PP(16'h1D12A,4);
TASK_PP(16'h1D12B,4);
TASK_PP(16'h1D12C,4);
TASK_PP(16'h1D12D,4);
TASK_PP(16'h1D12E,4);
TASK_PP(16'h1D12F,4);
TASK_PP(16'h1D130,4);
TASK_PP(16'h1D131,4);
TASK_PP(16'h1D132,4);
TASK_PP(16'h1D133,4);
TASK_PP(16'h1D134,4);
TASK_PP(16'h1D135,4);
TASK_PP(16'h1D136,4);
TASK_PP(16'h1D137,4);
TASK_PP(16'h1D138,4);
TASK_PP(16'h1D139,4);
TASK_PP(16'h1D13A,4);
TASK_PP(16'h1D13B,4);
TASK_PP(16'h1D13C,4);
TASK_PP(16'h1D13D,4);
TASK_PP(16'h1D13E,4);
TASK_PP(16'h1D13F,4);
TASK_PP(16'h1D140,4);
TASK_PP(16'h1D141,4);
TASK_PP(16'h1D142,4);
TASK_PP(16'h1D143,4);
TASK_PP(16'h1D144,4);
TASK_PP(16'h1D145,4);
TASK_PP(16'h1D146,4);
TASK_PP(16'h1D147,4);
TASK_PP(16'h1D148,4);
TASK_PP(16'h1D149,4);
TASK_PP(16'h1D14A,4);
TASK_PP(16'h1D14B,4);
TASK_PP(16'h1D14C,4);
TASK_PP(16'h1D14D,4);
TASK_PP(16'h1D14E,4);
TASK_PP(16'h1D14F,4);
TASK_PP(16'h1D150,4);
TASK_PP(16'h1D151,4);
TASK_PP(16'h1D152,4);
TASK_PP(16'h1D153,4);
TASK_PP(16'h1D154,4);
TASK_PP(16'h1D155,4);
TASK_PP(16'h1D156,4);
TASK_PP(16'h1D157,4);
TASK_PP(16'h1D158,4);
TASK_PP(16'h1D159,4);
TASK_PP(16'h1D15A,4);
TASK_PP(16'h1D15B,4);
TASK_PP(16'h1D15C,4);
TASK_PP(16'h1D15D,4);
TASK_PP(16'h1D15E,4);
TASK_PP(16'h1D15F,4);
TASK_PP(16'h1D160,4);
TASK_PP(16'h1D161,4);
TASK_PP(16'h1D162,4);
TASK_PP(16'h1D163,4);
TASK_PP(16'h1D164,4);
TASK_PP(16'h1D165,4);
TASK_PP(16'h1D166,4);
TASK_PP(16'h1D167,4);
TASK_PP(16'h1D168,4);
TASK_PP(16'h1D169,4);
TASK_PP(16'h1D16A,4);
TASK_PP(16'h1D16B,4);
TASK_PP(16'h1D16C,4);
TASK_PP(16'h1D16D,4);
TASK_PP(16'h1D16E,4);
TASK_PP(16'h1D16F,4);
TASK_PP(16'h1D170,4);
TASK_PP(16'h1D171,4);
TASK_PP(16'h1D172,4);
TASK_PP(16'h1D173,4);
TASK_PP(16'h1D174,4);
TASK_PP(16'h1D175,4);
TASK_PP(16'h1D176,4);
TASK_PP(16'h1D177,4);
TASK_PP(16'h1D178,4);
TASK_PP(16'h1D179,4);
TASK_PP(16'h1D17A,4);
TASK_PP(16'h1D17B,4);
TASK_PP(16'h1D17C,4);
TASK_PP(16'h1D17D,4);
TASK_PP(16'h1D17E,4);
TASK_PP(16'h1D17F,4);
TASK_PP(16'h1D180,4);
TASK_PP(16'h1D181,4);
TASK_PP(16'h1D182,4);
TASK_PP(16'h1D183,4);
TASK_PP(16'h1D184,4);
TASK_PP(16'h1D185,4);
TASK_PP(16'h1D186,4);
TASK_PP(16'h1D187,4);
TASK_PP(16'h1D188,4);
TASK_PP(16'h1D189,4);
TASK_PP(16'h1D18A,4);
TASK_PP(16'h1D18B,4);
TASK_PP(16'h1D18C,4);
TASK_PP(16'h1D18D,4);
TASK_PP(16'h1D18E,4);
TASK_PP(16'h1D18F,4);
TASK_PP(16'h1D190,4);
TASK_PP(16'h1D191,4);
TASK_PP(16'h1D192,4);
TASK_PP(16'h1D193,4);
TASK_PP(16'h1D194,4);
TASK_PP(16'h1D195,4);
TASK_PP(16'h1D196,4);
TASK_PP(16'h1D197,4);
TASK_PP(16'h1D198,4);
TASK_PP(16'h1D199,4);
TASK_PP(16'h1D19A,4);
TASK_PP(16'h1D19B,4);
TASK_PP(16'h1D19C,4);
TASK_PP(16'h1D19D,4);
TASK_PP(16'h1D19E,4);
TASK_PP(16'h1D19F,4);
TASK_PP(16'h1D1A0,4);
TASK_PP(16'h1D1A1,4);
TASK_PP(16'h1D1A2,4);
TASK_PP(16'h1D1A3,4);
TASK_PP(16'h1D1A4,4);
TASK_PP(16'h1D1A5,4);
TASK_PP(16'h1D1A6,4);
TASK_PP(16'h1D1A7,4);
TASK_PP(16'h1D1A8,4);
TASK_PP(16'h1D1A9,4);
TASK_PP(16'h1D1AA,4);
TASK_PP(16'h1D1AB,4);
TASK_PP(16'h1D1AC,4);
TASK_PP(16'h1D1AD,4);
TASK_PP(16'h1D1AE,4);
TASK_PP(16'h1D1AF,4);
TASK_PP(16'h1D1B0,4);
TASK_PP(16'h1D1B1,4);
TASK_PP(16'h1D1B2,4);
TASK_PP(16'h1D1B3,4);
TASK_PP(16'h1D1B4,4);
TASK_PP(16'h1D1B5,4);
TASK_PP(16'h1D1B6,4);
TASK_PP(16'h1D1B7,4);
TASK_PP(16'h1D1B8,4);
TASK_PP(16'h1D1B9,4);
TASK_PP(16'h1D1BA,4);
TASK_PP(16'h1D1BB,4);
TASK_PP(16'h1D1BC,4);
TASK_PP(16'h1D1BD,4);
TASK_PP(16'h1D1BE,4);
TASK_PP(16'h1D1BF,4);
TASK_PP(16'h1D1C0,4);
TASK_PP(16'h1D1C1,4);
TASK_PP(16'h1D1C2,4);
TASK_PP(16'h1D1C3,4);
TASK_PP(16'h1D1C4,4);
TASK_PP(16'h1D1C5,4);
TASK_PP(16'h1D1C6,4);
TASK_PP(16'h1D1C7,4);
TASK_PP(16'h1D1C8,4);
TASK_PP(16'h1D1C9,4);
TASK_PP(16'h1D1CA,4);
TASK_PP(16'h1D1CB,4);
TASK_PP(16'h1D1CC,4);
TASK_PP(16'h1D1CD,4);
TASK_PP(16'h1D1CE,4);
TASK_PP(16'h1D1CF,4);
TASK_PP(16'h1D1D0,4);
TASK_PP(16'h1D1D1,4);
TASK_PP(16'h1D1D2,4);
TASK_PP(16'h1D1D3,4);
TASK_PP(16'h1D1D4,4);
TASK_PP(16'h1D1D5,4);
TASK_PP(16'h1D1D6,4);
TASK_PP(16'h1D1D7,4);
TASK_PP(16'h1D1D8,4);
TASK_PP(16'h1D1D9,4);
TASK_PP(16'h1D1DA,4);
TASK_PP(16'h1D1DB,4);
TASK_PP(16'h1D1DC,4);
TASK_PP(16'h1D1DD,4);
TASK_PP(16'h1D1DE,4);
TASK_PP(16'h1D1DF,4);
TASK_PP(16'h1D1E0,4);
TASK_PP(16'h1D1E1,4);
TASK_PP(16'h1D1E2,4);
TASK_PP(16'h1D1E3,4);
TASK_PP(16'h1D1E4,4);
TASK_PP(16'h1D1E5,4);
TASK_PP(16'h1D1E6,4);
TASK_PP(16'h1D1E7,4);
TASK_PP(16'h1D1E8,4);
TASK_PP(16'h1D1E9,4);
TASK_PP(16'h1D1EA,4);
TASK_PP(16'h1D1EB,4);
TASK_PP(16'h1D1EC,4);
TASK_PP(16'h1D1ED,4);
TASK_PP(16'h1D1EE,4);
TASK_PP(16'h1D1EF,4);
TASK_PP(16'h1D1F0,4);
TASK_PP(16'h1D1F1,4);
TASK_PP(16'h1D1F2,4);
TASK_PP(16'h1D1F3,4);
TASK_PP(16'h1D1F4,4);
TASK_PP(16'h1D1F5,4);
TASK_PP(16'h1D1F6,4);
TASK_PP(16'h1D1F7,4);
TASK_PP(16'h1D1F8,4);
TASK_PP(16'h1D1F9,4);
TASK_PP(16'h1D1FA,4);
TASK_PP(16'h1D1FB,4);
TASK_PP(16'h1D1FC,4);
TASK_PP(16'h1D1FD,4);
TASK_PP(16'h1D1FE,4);
TASK_PP(16'h1D1FF,4);
TASK_PP(16'h1D200,4);
TASK_PP(16'h1D201,4);
TASK_PP(16'h1D202,4);
TASK_PP(16'h1D203,4);
TASK_PP(16'h1D204,4);
TASK_PP(16'h1D205,4);
TASK_PP(16'h1D206,4);
TASK_PP(16'h1D207,4);
TASK_PP(16'h1D208,4);
TASK_PP(16'h1D209,4);
TASK_PP(16'h1D20A,4);
TASK_PP(16'h1D20B,4);
TASK_PP(16'h1D20C,4);
TASK_PP(16'h1D20D,4);
TASK_PP(16'h1D20E,4);
TASK_PP(16'h1D20F,4);
TASK_PP(16'h1D210,4);
TASK_PP(16'h1D211,4);
TASK_PP(16'h1D212,4);
TASK_PP(16'h1D213,4);
TASK_PP(16'h1D214,4);
TASK_PP(16'h1D215,4);
TASK_PP(16'h1D216,4);
TASK_PP(16'h1D217,4);
TASK_PP(16'h1D218,4);
TASK_PP(16'h1D219,4);
TASK_PP(16'h1D21A,4);
TASK_PP(16'h1D21B,4);
TASK_PP(16'h1D21C,4);
TASK_PP(16'h1D21D,4);
TASK_PP(16'h1D21E,4);
TASK_PP(16'h1D21F,4);
TASK_PP(16'h1D220,4);
TASK_PP(16'h1D221,4);
TASK_PP(16'h1D222,4);
TASK_PP(16'h1D223,4);
TASK_PP(16'h1D224,4);
TASK_PP(16'h1D225,4);
TASK_PP(16'h1D226,4);
TASK_PP(16'h1D227,4);
TASK_PP(16'h1D228,4);
TASK_PP(16'h1D229,4);
TASK_PP(16'h1D22A,4);
TASK_PP(16'h1D22B,4);
TASK_PP(16'h1D22C,4);
TASK_PP(16'h1D22D,4);
TASK_PP(16'h1D22E,4);
TASK_PP(16'h1D22F,4);
TASK_PP(16'h1D230,4);
TASK_PP(16'h1D231,4);
TASK_PP(16'h1D232,4);
TASK_PP(16'h1D233,4);
TASK_PP(16'h1D234,4);
TASK_PP(16'h1D235,4);
TASK_PP(16'h1D236,4);
TASK_PP(16'h1D237,4);
TASK_PP(16'h1D238,4);
TASK_PP(16'h1D239,4);
TASK_PP(16'h1D23A,4);
TASK_PP(16'h1D23B,4);
TASK_PP(16'h1D23C,4);
TASK_PP(16'h1D23D,4);
TASK_PP(16'h1D23E,4);
TASK_PP(16'h1D23F,4);
TASK_PP(16'h1D240,4);
TASK_PP(16'h1D241,4);
TASK_PP(16'h1D242,4);
TASK_PP(16'h1D243,4);
TASK_PP(16'h1D244,4);
TASK_PP(16'h1D245,4);
TASK_PP(16'h1D246,4);
TASK_PP(16'h1D247,4);
TASK_PP(16'h1D248,4);
TASK_PP(16'h1D249,4);
TASK_PP(16'h1D24A,4);
TASK_PP(16'h1D24B,4);
TASK_PP(16'h1D24C,4);
TASK_PP(16'h1D24D,4);
TASK_PP(16'h1D24E,4);
TASK_PP(16'h1D24F,4);
TASK_PP(16'h1D250,4);
TASK_PP(16'h1D251,4);
TASK_PP(16'h1D252,4);
TASK_PP(16'h1D253,4);
TASK_PP(16'h1D254,4);
TASK_PP(16'h1D255,4);
TASK_PP(16'h1D256,4);
TASK_PP(16'h1D257,4);
TASK_PP(16'h1D258,4);
TASK_PP(16'h1D259,4);
TASK_PP(16'h1D25A,4);
TASK_PP(16'h1D25B,4);
TASK_PP(16'h1D25C,4);
TASK_PP(16'h1D25D,4);
TASK_PP(16'h1D25E,4);
TASK_PP(16'h1D25F,4);
TASK_PP(16'h1D260,4);
TASK_PP(16'h1D261,4);
TASK_PP(16'h1D262,4);
TASK_PP(16'h1D263,4);
TASK_PP(16'h1D264,4);
TASK_PP(16'h1D265,4);
TASK_PP(16'h1D266,4);
TASK_PP(16'h1D267,4);
TASK_PP(16'h1D268,4);
TASK_PP(16'h1D269,4);
TASK_PP(16'h1D26A,4);
TASK_PP(16'h1D26B,4);
TASK_PP(16'h1D26C,4);
TASK_PP(16'h1D26D,4);
TASK_PP(16'h1D26E,4);
TASK_PP(16'h1D26F,4);
TASK_PP(16'h1D270,4);
TASK_PP(16'h1D271,4);
TASK_PP(16'h1D272,4);
TASK_PP(16'h1D273,4);
TASK_PP(16'h1D274,4);
TASK_PP(16'h1D275,4);
TASK_PP(16'h1D276,4);
TASK_PP(16'h1D277,4);
TASK_PP(16'h1D278,4);
TASK_PP(16'h1D279,4);
TASK_PP(16'h1D27A,4);
TASK_PP(16'h1D27B,4);
TASK_PP(16'h1D27C,4);
TASK_PP(16'h1D27D,4);
TASK_PP(16'h1D27E,4);
TASK_PP(16'h1D27F,4);
TASK_PP(16'h1D280,4);
TASK_PP(16'h1D281,4);
TASK_PP(16'h1D282,4);
TASK_PP(16'h1D283,4);
TASK_PP(16'h1D284,4);
TASK_PP(16'h1D285,4);
TASK_PP(16'h1D286,4);
TASK_PP(16'h1D287,4);
TASK_PP(16'h1D288,4);
TASK_PP(16'h1D289,4);
TASK_PP(16'h1D28A,4);
TASK_PP(16'h1D28B,4);
TASK_PP(16'h1D28C,4);
TASK_PP(16'h1D28D,4);
TASK_PP(16'h1D28E,4);
TASK_PP(16'h1D28F,4);
TASK_PP(16'h1D290,4);
TASK_PP(16'h1D291,4);
TASK_PP(16'h1D292,4);
TASK_PP(16'h1D293,4);
TASK_PP(16'h1D294,4);
TASK_PP(16'h1D295,4);
TASK_PP(16'h1D296,4);
TASK_PP(16'h1D297,4);
TASK_PP(16'h1D298,4);
TASK_PP(16'h1D299,4);
TASK_PP(16'h1D29A,4);
TASK_PP(16'h1D29B,4);
TASK_PP(16'h1D29C,4);
TASK_PP(16'h1D29D,4);
TASK_PP(16'h1D29E,4);
TASK_PP(16'h1D29F,4);
TASK_PP(16'h1D2A0,4);
TASK_PP(16'h1D2A1,4);
TASK_PP(16'h1D2A2,4);
TASK_PP(16'h1D2A3,4);
