// ***************************************************************************************
// *
// * File Name: RUNP.vh
// * /RCS/ RUNL.vh Version: 1.00 12/06/2012
// *
// *******************************************************      
// *
// * Change_list 
// * Version Author Date Changes 
// * 1.0 G.Grise 05/18/11 initial coding 
// *
// *
// *_limitations : only works when BAMC chip is actually Macronix model clone  
// * 
// * 
// * Errors : 
// * 
// *
// **************************************************************************************** 
// * Description Run does:  
//   normal power-up and reset.  - part of spi_task_check_exps.vh
// 1) write to address 000000 should pass TASK_INIT_WRITE_PI TASK_PP2(16'h0000,256); 
// 2) WRITE INTO LAYER BUFFER;
// 3) READ LAYER BUFFER   
// 
// 	-	 -		-		-	    -		-		-	 -	 
// **************************************************************************************** 
	RUN_NUMBER = "P" ;
`include "./banners/+runP_start.vh"	        
`include "./banners/+test1.vh"
$display ("write to address 000000 should pass  ") ;

TASK_RSTEN;
TASK_RST;
//loadmem;

//TASK_SCE(0,160'h0111114325466878700,4'h1,8'h01,4'h1,16'h201,1,1,0,8'h11,64'h019219384010402,200'h1222645454554343435222227);

//TASK_SCEWAF(4096'b0000000000000000000000000000000000100110000000000000000000000000000100110000000000000000000000000011010010000000000000000000000000001001100000000000000000000000001011111000000000000000000000000001101001000000000000000000000000111101010000000000000000000000000001001100000000000000000000000010000111000000000000000000000000010111110000000000000000000000001100100010000000000000000000000000110100100000000000000000000000101000101000000000000000000000000111101010000000000000000000000011101110100000000000000000000000000010011000000000000000000000001001010110000000000000000000000001000011100000000000000000000000110110111000000000000000000000000010111110000000000000000000000010110000010000000000000000000000011001000100000000000000000000001111110001000000000000000000000000011010010000000000000000000000100011100100000000000000000000000101000101000000000000000000000011000101010000000000000000000000001111010100000000000000000000001010101101000000000000000000000001110111010000000000000000000000111000001100000000000000000000000000010011000000000000000000000010011100110000000000000000000000010010101100000000000000000000001101011011000000000000000000000000100001110000000000000000000000101110011100000000000000000000000110110111000000000000000000000011110011110000000000000000000000000101111100000000000000000000001000000000100000000000000000000001011000001000000000000000000000110011000010000000000000000000000011001000100000000000000000000010100110001000000000000000000000011111100010000000000000000000001110100100100000000000000000000000001101001000000000000000000000100100110010000000000000000000000100011100100000000000000000000011011111001000000000000000000000001010001010000000000000000000001011010010100000000000000000000001100010101000000000000000000000111110101010000000000000000000000001111010100000000000000000000010001001101000000000000000000000010101011010000000000000000000001100001110100000000000000000000000111011101000000000000000000000101011111010000000000000000000000111000001100000000000000000000011100100011000000000000000000000000000100110000000000000000000001001101001100000000000000000000001001110011000000000000000000000110100010110000000000000000000000010010101100000000000000000000010111101011000000000000000000000011010110110000000000000000000001111011101100000000000000000000000010000111000000000000000000000100001001110000000000000000000000101110011100000000000000000000011001010111000000000000000000000001101101110000000000000000000001010000111100000000000000000000001111001111000000000000000000000111011011110000000000000000000000000101111100000000000000000000010010111111000000000000000000000010000000001000000000000000000001101100000010000000000000000000000101100000100000000000000000000101100100001000000000000000000000110011000010000000000000000000011111110000100000000000000000000000110010001000000000000000000001000110100010000000000000000000001010011000100000000000000000000110001110001000000000000000000000011111100010000000000000000000010101000100100000000000000000000011101001001000000000000000000001110001010010000000000000000000000000110100100000000000000000000100111101001000000000000000000000100100110010000000000000000000011010101100100000000000000000000001000111001000000000000000000001011101110010000000000000000000001101111100100000000000000000000111100000101000000000000000000000001010001010000000000000000000010000010010100000000000000000000010110100101000000000000000000001100111001010000000000000000000000110001010100000000000000000000101001010101000000000000000000000111110101010000000000000000000011101011010100000000000000000000000011110101000000000000000000001001000011010000000000000000000001000100110100000000000000000000110111001101000000000000000000000010101011010000000000000000000010110110110100000000000000000000011000011101000000000000000000001111100111010000000000000000000000011101110100000000000000000000100010111101000000000000000000000101011111010000000000000000000011000000001100000000000000000000001110000011000000000000000000001010110000110000000000000000000001110010001100000000000000000000111001100011000000000000000000, 4096'b0000000001001100000000000000000000100110010011000000000000000000000100110100110000000000000000000011010011001100000000000000000000001001110011000000000000000000001011111100110000000000000000000001101000101100000000000000000000111101001011000000000000000000000001001010110000000000000000000010000110101100000000000000000000010111101011000000000000000000001100100110110000000000000000000000110101101100000000000000000000101000111011000000000000000000000111101110110000000000000000000011101111101100000000000000000000000010000111000000000000000000001001010001110000000000000000000001000010011100000000000000000000110110100111000000000000000000000010111001110000000000000000000010110001011100000000000000000000011001010111000000000000000000001111110101110000000000000000000000011011011100000000000000000000100011110111000000000000000000000101000011110000000000000000000011000100111100000000000000000000001111001111000000000000000000001010101011110000000000000000000001110110111100000000000000000000111000011111000000000000000000000000010111110000000000000000000010011101111100000000000000000000010010111111000000000000000000001101011111110000000000000000000000100000000010000000000000000000101110000000100000000000000000000110110000001000000000000000000011110010000010000000000000000000000101100000100000000000000000001000000100001000000000000000000001011001000010000000000000000000110011010000100000000000000000000011001100001000000000000000000010100111000010000000000000000000011111110000100000000000000000001110100010001000000000000000000000001100100010000000000000000000100100101000100000000000000000000100011010001000000000000000000011011110100010000000000000000000001010011000100000000000000000001011010110001000000000000000000001100011100010000000000000000000111110111000100000000000000000000001111110001000000000000000000010001000010010000000000000000000010101000100100000000000000000001100001001001000000000000000000000111010010010000000000000000000101011100100100000000000000000000111000101001000000000000000000011100101010010000000000000000000000000110100100000000000000000001001101101001000000000000000000001001111010010000000000000000000110100001100100000000000000000000010010011001000000000000000000010111100110010000000000000000000011010101100100000000000000000001111011011001000000000000000000000010001110010000000000000000000100001011100100000000000000000000101110111001000000000000000000011001011110010000000000000000000001101111100100000000000000000001010000000101000000000000000000001111000001010000000000000000000111011000010100000000000000000000000101000101000000000000000000010010110001010000000000000000000010000010010100000000000000000001101100100101000000000000000000000101101001010000000000000000000101100110010100000000000000000000110011100101000000000000000000011111111001010000000000000000000000110001010100000000000000000001000110010101000000000000000000001010010101010000000000000000000110001101010100000000000000000000011111010101000000000000000000010101001101010000000000000000000011101011010100000000000000000001110001110101000000000000000000000000111101010000000000000000000100111111010100000000000000000000100100001101000000000000000000011010100011010000000000000000000001000100110100000000000000000001011101001101000000000000000000001101110011010000000000000000000111100010110100000000000000000000001010101101000000000000000000010000011011010000000000000000000010110110110100000000000000000001100111101101000000000000000000000110000111010000000000000000000101001001110100000000000000000000111110011101000000000000000000011101010111010000000000000000000000011101110100000000000000000001001000111101000000000000000000001000101111010000000000000000000110111011110100000000000000000000010101111101000000000000000000010110111111010000000000000000000011000000001100000000000000000001111100000011000000000000000000000011100000110000000000000000000100010100001100000000000000000000101011000011000000000000000000011000001000110000000000000000000001110010001100000000000000000001010110100011000000000000000000001110011000110000000000000000000111001110001100000000000000000,160'hBFEDF72429B023D37D0D724D00A1248DB0FEAD3,4'h1,8'h22,4'h2,16'h2313,1,1,0,8'hAB,64'h2333333333321212,3828'h0111111111111111111111111111111111111111111111111111111111011111111111111111111111111111110101001010101010101010101010101010101010109F1,4096'h89, 573'h0);


TASK_EXPECT_PASS ;
$display ("============================================================") ;         


//TASK_NOP;

`include "./banners/+test1.vh"
$display ("write to address 000000 should pass  ") ;
TASK_INIT_WRITE_PI ;    
TASK_LBWR(16'h0001);
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;


`include "./banners/+test2.vh"
$display ("READ LAYER BUFFER") ;
TASK_RDLB(1);
TASK_EXPECT_PASS ;              
$display ("============================================================") ;

TASK_NOP;

`include "./banners/+test3.vh"
$display ("lock sector 0") ;    
//TASK_INIT_WRITE_PI;
TASK_INIT_WRITE_ONES;
TASK_PP(16'h0010,4);
// do expect checking
TASK_EXPECT_PASS ;              
$display ("============================================================") ;
    

`include "./banners/+test3.vh"
$display ("lock sector 0") ;    
TASK_INIT_WRITE_PI;
//TASK_INIT_WRITE_ONES;
TASK_PP(16'h0011,4);
// do expect checking
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;
      

`include "./banners/+test3.vh"
$display ("lock sector 0") ;    
TASK_INIT_WRITE_PI;
//TASK_INIT_WRITE_ONES;
TASK_PP(16'h0012,4);
// do expect checking
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;       


`include "./banners/+test3.vh"
$display ("lock sector 0") ;    
//TASK_INIT_WRITE_PI;
TASK_INIT_WRITE_ZEROS;
TASK_PP(16'h0013,4);
// do expect checking
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;
       

`include "./banners/+test4.vh"
$display ("lock sector 0") ;    
TASK_READ_READ(16'h0012,4);
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;


TASK_NOP;

`include "./banners/+test4.vh"
$display ("lock sector 0") ;    
TASK_READ_READ(16'h0013,4);
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;


TASK_NOP;

`include "./banners/+test4.vh"
$display ("lock sector 0") ;    
TASK_READ_READ(16'h0010,4);
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;


TASK_NOP;


`include "./banners/+test5.vh"
//TASK_INIT_WRITE_PI;
//TASK_INIT_WRITE_ONES;
TASK_MACCYC(0,32'h00100001);
//TASK_EXPECT_PASS ;              
//$display ("============================================================") ;


`include "./banners/+test6.vh"
TASK_INIT_WRITE_PI;
//TASK_INIT_WRITE_ONES;
TASK_BIASBUF(3,16'h0010);
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;


`include "./banners/+test6.vh"
//TASK_INIT_WRITE_PI;
//TASK_INIT_WRITE_ONES;
TASK_NEURONACT(32'h00100001);
//TASK_EXPECT_PASS ;              
$display ("============================================================") ;
        

`include "./banners/+runP_end.vh"	
