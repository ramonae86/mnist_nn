`include "./banners/+runP_start.vh"
`include "./banners/+test1.vh"
TASK_RSTEN;
TASK_RST;
