
// Verilog stimulus file.
`include "/proj/bingen/models/m31/M31GPSC900HL040PR_50N.v"
`include "/proj/bingen/models/m31/M31GPSC900HL040PH_50N_pwr.v"
`include "/home/don/workspace/bingen/M31GPSC900HL040PR_50N_pwr_del.v"
//`include "/proj/bingen/models/udp/M31GPSC900HL040PH_50N.v"
//`include "/proj/bingen/models/udp/M31GPSC900HL040PH_50N_pwr.v"
//`include "/proj/punk/20180206/HL40LPGP3VDIB03P1_DK/verilog/HL40LPGP2VDIB03.v"

// Default verilog stimulus. 

`timescale 1ns / 1ps


module testbench();

   
   parameter 
     por_cmd = 8'b11110000, 
     reset_mul_cmd = 8'b01100000,
     latch_acc_cmd = 8'b10100000,
     reset_acc_cmd = 8'b00100000,
     loadtm_cmd = 8'b11000000,
     write_cmd = 8'b01000000,
     read_cmd = 8'b10000000,
     nop_cmd = 8'b00000000,
     lbread_cmd = 8'b11100000,
     lbwrite_cmd = 8'b00010000,
     pd_act_cmd = 8'b01000000,
     latch_mul_cmd = 8'b01010000,
     bias_clk0_cmd = 8'b11010000,
     bias_clk1_cmd = 8'b00110000,
     bias_clk2_cmd = 8'b10110000,
     bias_clk3_cmd = 8'b01110000;
   
   wire VCC;
   wire VSS;
   
   
   //wire VDD;
   wire SO_P;
   wire SI_P;
   wire ACLK_P;
   wire BCLK_P;
   wire CCLK_P;
   wire CSn_P;
   wire DIGMON_P;
   wire MODE_SEL_P;
   
   
   assign VCC = 1;
   assign VSS = 0;
   //assign VDD = 1;
   
   
   ////////////////////
   //Registers to for IO wires
   /////////////////////////
   reg 	SI_R;
   reg 	ACLK_R;
   reg 	BCLK_R;
   reg 	CCLK_R;
   reg 	CSn_R;
   reg 	DIGMON_R;
   reg 	MODE_SEL_R;
   reg 	LB_BCLK_R;
   reg 	LB_ACLK_R;
   
   assign SI_P   = SI_R;
   assign ACLK_P = ACLK_R;
   assign BCLK_P = BCLK_R;
   assign CCLK_P = CCLK_R;
   assign CSn_P  = CSn_R;
   assign MODE_SEL_P = MODE_SEL_R;
   assign DIGMON_P = DIGMON_R;
   assign LB_ACLK_P = LB_ACLK_R;
   assign LB_BCLK_P = LB_BCLK_R;

     
   reg 	LB_SEL = 0;
   reg [7:0] LB_IN;
   
   reg [1023:0] COMMAND;
   
   integer 	i;
   integer      j;
   integer 	k;
   
   integer 	wr;

   reg 		BIAS_SEL;
   reg 		READ;
   reg 		WRITE;
   reg [9:0] 	WA;
   reg [5:0] 	BA;
   reg [3:0] 	SAAD;
   reg [7:0] 	CMD;
   reg [3:0] 	WHDATA;
   reg [2:0] 	NC;
   reg [4:0] 	DIGMON;
   
   // Test Modes from 64 to 0:
   reg          SCAN;
   reg 		MACBUS_EN;
   reg          PRGM_AF;
   reg          LB_INP_SEL;
   reg  	TM_SIGN_PRE_AF;
   reg  	TM_SIGN_POST_AF;
   reg [3:0] 	TM_SETTLE_DONE;
   reg [1:0] 	TM_MACSEL;
   reg 		LB_BUFSEL;
   reg [3:0] 	TM_WRHPW;
   reg [1:0] 	TM_WR2WR_DLY;
   reg 		TM_WLE;
   reg [4:0] 	TM_SET;
   reg [1:0] 	TM_MACMODE;   
   reg [3:0] 	TM_READ_DONE;
   reg [3:0] 	TM_FTOP;
   reg [4:0] 	TM_WRLC;
   reg [4:0] 	TM_WRHC;
   reg [6:0] 	TM_SATRIM;
   reg 		TM_PCHG_SF_BYP;
   reg [3:0] 	TM_PCHG_SF;
   reg 		TM_PCHG_RH_BYP;
   reg [3:0] 	TM_PCHG_RH;
   reg 		TM_DATATEST;
   reg 		LB_ACT;
   
   //  reg [63:0] TM;
   wire [63:0] 	TM;  
   assign TM = { MACBUS_EN, PRGM_AF, LB_INP_SEL, TM_MACSEL, LB_ACT, LB_BUFSEL, SCAN, 56'b0};

   //reg [8191:0] AF_data = 8192'b00000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000011000000000000000000000000000000001000000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000111000000000000000000000000000000001000000000000000000000000000010010000000000000000000000000000010100000000000000000000000000001101000000000000000000000000000000110000000000000000000000000000101100000000000000000000000000000111000000000000000000000000000011110000000000000000000000000000000010000000000000000000000000001000100000000000000000000000000001001000000000000000000000000000110010000000000000000000000000000000010000000000000000000000000000001100000000000000000000000000000000100000000000000000000000000000101000000000000000000000000000100110000000000000000000000000000000010000000000000000000000000001000100000000000000000000000000000011000000000000000000000000000000001000000000000000000000000010000010000000000000000000000000001000100000000000000000000000000000011000000000000000000000000000011110000000000000000000000000000000010000000000000000000000000010000100000000000000000000000000001001000000000000000000000000000000110000000000000000000000000000000010000000000000000000000000000010100000000000000000000000000000011000000000000000000000000000000001000000000000000000000000100000010000000000000000000000010000000100000000000000000000000010000001000000000000000000000000010000010000000000000000000000000001000100000000000000000000000000000011000000000000000000000000000111110000000000000000000000000000000010000000000000000000000010000000100000000000000000000000001000001000000000000000000000000000010010000000000000000000000001000000010000000000000000000000000010000100000000000000000000000000001001000000000000000000000000000011110000000000000000000000000000000010000000000000000000010000000000100000000000000000000000010000001000000000000000000000000000100010000000000000000000000000000010100000000000000000000000000000011000000000000000000000000000111110000000000000000000000000000000010000000000000000000100000000000100000000000000000000001000000001000000000000000000000001000000010000000000000000000000000010000100000000000000000000000000001001000000000000000000000000000001010000000000000000000000000011111100000000000000000000000000000000100000000000000000010000000000001000000000000000000000100000000010000000000000000000000100000000100000000000000000000000100000001000000000000000000000000010000010000000000000000000000000010000100000000000000000000000000010001000000000000000000000000000010010000000000000000000000000000111100000000000000000000000000000000100000000000000000010000000000001000000000000000000010000000000010000000000000000000010000000000100000000000000000000010000000001000000000000000000000010000000010000000000000000000000010000000100000000000000000000000010000001000000000000000000000000001000010000000000000000000000000000010100000000000000000000000000001111000000000000000000011111111111110000000000000000000000000000000010000000000000000100000000000000100000000000000000010000000000001000000000000000000110000000000010000000000000000000011000000000100000000000000000000000010000001000000000000000000000000001000010000000000000000000000000000100100000000000000000000000000000101000000000000000000000000001111110000000000000000000000000000000010000000000000010000000000000000100000000000000010000000000000001000000000000000010000000000000010000000000000000010000000000000100000000000000000010000000000001000000000000000000010000000000010000000000000000000001000000000100000000000000000000001000000001000000000000000000000001000000010000000000000000000000000100000100000000000000000000000000010001000000000000000000000000000010010000000000000000000000000000011100000000000000000000000000000000100000000000001000000000000000001000000000000001000000000000000010000000000000001000000000000000100000000000000001000000000000001000000000000000001000000000000010000000000000000001000000000000100000000000000000001000000000001000000000000000000001000000000010000000000000000000001000000000100000000000000000000001000000001000000000000000000000001000000010000000000000000000000001000000100000000000000000000000001000001000000000000000000000000001000010000000000000000000000000001000100000000000000000000000000001001000000000000000000000000000001010000000000000000000000000001110100000000000000100000000000000011000000000001001000000000000000110000000000001110000000000000001100000000000110110000000000000011000000000000011010000000000000110000000000010110010000000000001100000000000011100010000000000011000000000001111000010000000000110000000000000001000000000000011100000000000100010000000000001111000000000000100100000000000111110000000000011001000000000111111000000000000111111111111111111110000000000000000000000000000000010000000000000100000000000000000100000000000000010000000000000001000000000000000010000000000000010000000000000000001000000000000100000000000000000001000000000001000000000000000000001000000000010000000000000000000001000000000100000000000000000000001000000001000000000000000000000001000000010000000000000000000000001000000100000000000000000000000001000001000000000000000000000000001000010000000000000000000000000001000100000000000000000000000000001001000000000000000000000000000001010000000000000000000000000000001100000000000001000000000000000011000000000000000100000000000000110000000000000000100000000000001100000000000000000100000000000011000000000000000000100000000000110000000000000000000100000000001100000000000000000000100000000011000000000000000000000100000000110000000000000000000000001000001100000000000000000000000001000011000000000000000000000000001000110000000000000000000000000001001100000000000000000000000000000111000000000000100000000000000001110000000000000100000000000000011100000000000000100000000000000111000000000000000100000000000001110000000000000000100000000000011100000000000000000100000000000111000000000000000000100000000001110000000000000000000100000000011100000000000000000000100000000111000000000000000000000100000001110000000000000000000000100000011100000000000000000000000100000111000000000000000000000000100001110000000000000000000000000100011100000000000000000000000000100111000000000000000000000000000101110000000000000000000000000000111100000000000010000000000000001111000000000000001000000000000011110000000000000001000000000000111100000000000000001000000000001111000000000000000001000000000011110000000000000000001000000000111100000000000000000001000000001111000000000000000000001000000011110000000000000000000001000000111100000000000000000000001000001111000000000000000000000001000011110000000000000000000000000100111100000000000000000000000000101111000000000000000000000000000111110000000000001000000000000001111100000000000001000000000000011111000000000000001000000000000111110000000000000001000000000001111100000000000000001000000000011111000000000000000001000000000111110000000000000000001000000001111100000000000000000001000000011111000000000000000000001000000111110000000000000000000001000001111100000000000000000000001000011111000000000000000000000001000111110000000000000000000000001001111100000000000000000000000001011111000000000000000000000000001111110000000000001000000000000011111100000000000001000000000000111111000000000000001000000000001111110000000000000001000000000011111100000000000000001000000000111111000000000000000001000000001111110000000000000000001000000011111100000000000000000001000000111111000000000000000000001000001111110000000000000000000001000011111100000000000000000000001000111111000000000000000000000001001111110000000000000000000000001011111100000000000000000000000001111111000000000000100000000000011111110000000000000100000000000111111100000000000000100000000001111111000000000000000100000000011111110000000000000000100000000111111100000000000000000100000001111111000000000000000000100000011111110000000000000000000100000111111100000000000000000000100001111111000000000000000000000100011111110000000000000000000000100111111100000000000000000000000101111111000000000000000000000000111111110000000000000000000000011111111100000000000001000000000111111111000000000000000100000001111111110000000000000000010000011111111100000000000; //random reg values that are forced by task.v in the original scan chain sim

   reg [8191:0] AF_data = 8192'b00000000000000000000000000000000001001100000000000000000000000000001001100000000000000000000000000110100100000000000000000000000000010011000000000000000000000000010111110000000000000000000000000011010010000000000000000000000001111010100000000000000000000000000010011000000000000000000000000100001110000000000000000000000000101111100000000000000000000000011001000100000000000000000000000001101001000000000000000000000001010001010000000000000000000000001111010100000000000000000000000111011101000000000000000000000000000100110000000000000000000000010010101100000000000000000000000010000111000000000000000000000001101101110000000000000000000000000101111100000000000000000000000101100000100000000000000000000000110010001000000000000000000000011111100010000000000000000000000000110100100000000000000000000001000111001000000000000000000000001010001010000000000000000000000110001010100000000000000000000000011110101000000000000000000000010101011010000000000000000000000011101110100000000000000000000001110000011000000000000000000000000000100110000000000000000000000100111001100000000000000000000000100101011000000000000000000000011010110110000000000000000000000001000011100000000000000000000001011100111000000000000000000000001101101110000000000000000000000111100111100000000000000000000000001011111000000000000000000000010000000001000000000000000000000010110000010000000000000000000001100110000100000000000000000000000110010001000000000000000000000101001100010000000000000000000000111111000100000000000000000000011101001001000000000000000000000000011010010000000000000000000001001001100100000000000000000000001000111001000000000000000000000110111110010000000000000000000000010100010100000000000000000000010110100101000000000000000000000011000101010000000000000000000001111101010100000000000000000000000011110101000000000000000000000100010011010000000000000000000000101010110100000000000000000000011000011101000000000000000000000001110111010000000000000000000001010111110100000000000000000000001110000011000000000000000000000111001000110000000000000000000000000001001100000000000000000000010011010011000000000000000000000010011100110000000000000000000001101000101100000000000000000000000100101011000000000000000000000101111010110000000000000000000000110101101100000000000000000000011110111011000000000000000000000000100001110000000000000000000001000010011100000000000000000000001011100111000000000000000000000110010101110000000000000000000000011011011100000000000000000000010100001111000000000000000000000011110011110000000000000000000001110110111100000000000000000000000001011111000000000000000000000100101111110000000000000000000000100000000010000000000000000000011011000000100000000000000000000001011000001000000000000000000001011001000010000000000000000000001100110000100000000000000000000111111100001000000000000000000000001100100010000000000000000000010001101000100000000000000000000010100110001000000000000000000001100011100010000000000000000000000111111000100000000000000000000101010001001000000000000000000000111010010010000000000000000000011100010100100000000000000000000000001101001000000000000000000001001111010010000000000000000000001001001100100000000000000000000110101011001000000000000000000000010001110010000000000000000000010111011100100000000000000000000011011111001000000000000000000001111000001010000000000000000000000010100010100000000000000000000100000100101000000000000000000000101101001010000000000000000000011001110010100000000000000000000001100010101000000000000000000001010010101010000000000000000000001111101010100000000000000000000111010110101000000000000000000000000111101010000000000000000000010010000110100000000000000000000010001001101000000000000000000001101110011010000000000000000000000101010110100000000000000000000101101101101000000000000000000000110000111010000000000000000000011111001110100000000000000000000000111011101000000000000000000001000101111010000000000000000000001010111110100000000000000000000110000000011000000000000000000000011100000110000000000000000000010101100001100000000000000000000011100100011000000000000000000001110011000110000000000000000000000000001001100000000000000000000100110010011000000000000000000000100110100110000000000000000000011010011001100000000000000000000001001110011000000000000000000001011111100110000000000000000000001101000101100000000000000000000111101001011000000000000000000000001001010110000000000000000000010000110101100000000000000000000010111101011000000000000000000001100100110110000000000000000000000110101101100000000000000000000101000111011000000000000000000000111101110110000000000000000000011101111101100000000000000000000000010000111000000000000000000001001010001110000000000000000000001000010011100000000000000000000110110100111000000000000000000000010111001110000000000000000000010110001011100000000000000000000011001010111000000000000000000001111110101110000000000000000000000011011011100000000000000000000100011110111000000000000000000000101000011110000000000000000000011000100111100000000000000000000001111001111000000000000000000001010101011110000000000000000000001110110111100000000000000000000111000011111000000000000000000000000010111110000000000000000000010011101111100000000000000000000010010111111000000000000000000001101011111110000000000000000000000100000000010000000000000000000101110000000100000000000000000000110110000001000000000000000000011110010000010000000000000000000000101100000100000000000000000001000000100001000000000000000000001011001000010000000000000000000110011010000100000000000000000000011001100001000000000000000000010100111000010000000000000000000011111110000100000000000000000001110100010001000000000000000000000001100100010000000000000000000100100101000100000000000000000000100011010001000000000000000000011011110100010000000000000000000001010011000100000000000000000001011010110001000000000000000000001100011100010000000000000000000111110111000100000000000000000000001111110001000000000000000000010001000010010000000000000000000010101000100100000000000000000001100001001001000000000000000000000111010010010000000000000000000101011100100100000000000000000000111000101001000000000000000000011100101010010000000000000000000000000110100100000000000000000001001101101001000000000000000000001001111010010000000000000000000110100001100100000000000000000000010010011001000000000000000000010111100110010000000000000000000011010101100100000000000000000001111011011001000000000000000000000010001110010000000000000000000100001011100100000000000000000000101110111001000000000000000000011001011110010000000000000000000001101111100100000000000000000001010000000101000000000000000000001111000001010000000000000000000111011000010100000000000000000000000101000101000000000000000000010010110001010000000000000000000010000010010100000000000000000001101100100101000000000000000000000101101001010000000000000000000101100110010100000000000000000000110011100101000000000000000000011111111001010000000000000000000000110001010100000000000000000001000110010101000000000000000000001010010101010000000000000000000110001101010100000000000000000000011111010101000000000000000000010101001101010000000000000000000011101011010100000000000000000001110001110101000000000000000000000000111101010000000000000000000100111111010100000000000000000000100100001101000000000000000000011010100011010000000000000000000001000100110100000000000000000001011101001101000000000000000000001101110011010000000000000000000111100010110100000000000000000000001010101101000000000000000000010000011011010000000000000000000010110110110100000000000000000001100111101101000000000000000000000110000111010000000000000000000101001001110100000000000000000000111110011101000000000000000000011101010111010000000000000000000000011101110100000000000000000001001000111101000000000000000000001000101111010000000000000000000110111011110100000000000000000000010101111101000000000000000000010110111111010000000000000000000011000000001100000000000000000001111100000011000000000000000000000011100000110000000000000000000100010100001100000000000000000000101011000011000000000000000000011000001000110000000000000000000001110010001100000000000000000001010110100011000000000000000000001110011000110000000000000000000111001110001100000000000000000;
   
   
   //////////////////////////////////////////////////
   // TB STIMULUS SECTION
   //////////////////////////////////////////////////      
   `include "/proj/bingen/sim/00_TR/verilog/taskRZ.v"
   initial
     begin
	loadscanbits;

	MODE_SEL_R = 1;
	CSn_R = 1;
	ACLK_R = 0;
	BCLK_R = 0;
	CCLK_R = 0;
	LB_ACLK_R = 0;
	LB_BCLK_R = 0;
	DIGMON_R = 0;
	
	SI_R = 0;
	BIAS_SEL = 0;
	READ = 0;
	WRITE = 0;
	WA = 10'b0000000001;
	BA = 6'b000000;
	SAAD = 4'b0000;
	WHDATA = 4'b1001;
	NC = 3'b000;
	DIGMON = 5'b00000;
	COMMAND = "START";
	//TMs
	SCAN = 0;
	MACBUS_EN = 0;
	PRGM_AF = 0;
	LB_INP_SEL = 1;
	TM_MACSEL = 2'b00;
	LB_ACT = 0;
	LB_BUFSEL = 0;

	///////////////////////////////////////////////////
	//power on reset
	///////////////////////////////////////////////////
	CMD = por_cmd;	
	load_sc();	  
	runcommand(1000); // set C-Clock high for 1000ns
	
	#100
	  CMD = reset_mul_cmd;	
	load_sc();	  
	runcommand(10); // set C-Clock high for 1000ns

	#100
	  CMD = reset_acc_cmd;	
	load_sc();	  
	runcommand(10); // set C-Clock high for 1000ns

	#100
	  CMD = loadtm_cmd;
	load_sc();
	runcommand(10);

//	///////////////////////////////////////////////////
//	//program AF
//	///////////////////////////////////////////////////
//	#100
//	  PRGM_AF = 1;
//	SCAN = 1;
//	CMD = loadtm_cmd;
//	load_sc();
//	runcommand(10);
//
//	#100
//          scanAF(AF_data);
//
//	#100
//	  PRGM_AF = 0;
//	SCAN = 0;
//	CMD = loadtm_cmd;
//	load_sc();
//	runcommand(10);

	///////////////////////////////////////////////////
	//write data into array
	///////////////////////////////////////////////////
	#100
	  WA = 10'b1000000000;
	CMD = pd_act_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
        //four weights
	#100
	  writepattern(32'b00011000001111000111111000001011);

	#100
	  WA = 10'b1100000000;
	SAAD = 4'b0000;
	CMD = pd_act_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
        //four weights
	#100
	  writepattern(32'b10000001110000111110011100001000);

	#100
	  WA = 10'b1110000000;
	SAAD = 4'b0000;
	CMD = pd_act_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
        //one bias
	#100
	  writepattern(32'b00001111111100000101010110101010);

	#100
	  WA = 10'b1111000000;
	SAAD = 4'b0000;
	CMD = pd_act_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
        //another bias
	#100
	  writepattern(32'b00000000000010100000010100001111);

	#100
	  WA = 10'b1111100000;
	SAAD = 4'b0000;
	CMD = pd_act_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
        //still another bias
	#100
	  writepattern(32'b00000000000000000000000000000000);

	#100
	  WA = 10'b1111110000;
	SAAD = 4'b0000;
	CMD = pd_act_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
        //and another bias
	#100
	  writepattern(32'b00000000000000000000000000000000);

	///////////////////////////////////////////////////
	//write data into layer buffer
	///////////////////////////////////////////////////
	#100
	  LB_ACT = 1;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);
	
	#100
	  WA = 10'b0000000001;
	LB_IN = 8'b11001000;
	READ = 0;
	WRITE = 1;
	CMD = lbwrite_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);
        
	#100
	  WA = 10'b0000000011;
	LB_IN = 8'b10010110;
	CMD = lbwrite_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  LB_ACT = 0;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);
	
	///////////////////////////////////////////////////
	//read weight from array
	///////////////////////////////////////////////////
	#100
	  WA = 10'b1000000000;
	CMD = pd_act_cmd;
	READ = 1;
	WRITE = 0;
	load_sc();
	SI_R = 0;
	runcommand(10);

	///////////////////////////////////////////////////
	//read neuron value from layer buffer and MAC
	///////////////////////////////////////////////////
	#100
	  LB_ACT = 1;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);
	
	#100
	  WA = 10'b0000000001;
        CMD = lbread_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  baClock(8);

	#100
	  CMD = latch_acc_cmd;	
	load_sc();
	runcommand(10);
	
	#100
	  CMD = reset_mul_cmd;	
	load_sc();	  
	runcommand(10);

	#100
	  LB_ACT = 0;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	///////////////////////////////////////////////////
	//read the second weight from array
	///////////////////////////////////////////////////
	#100
	  WA = 10'b1100000000;
	CMD = pd_act_cmd;
	READ = 1;
	WRITE = 0;
	load_sc();
	SI_R = 0;
	runcommand(10);

	///////////////////////////////////////////////////
	//read neuron value from layer buffer and MAC
	///////////////////////////////////////////////////
	#100
	  LB_ACT = 1;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);
	
	#100
	  WA = 10'b0000000011;
        CMD = lbread_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
        runcommand(10);
	
	#100
	  baClock(8);
        
	#100
	  CMD = latch_acc_cmd;	
	load_sc();
	runcommand(10);

	#100
	  CMD = reset_mul_cmd;	
	load_sc();	  
	runcommand(10);

	#100
	  LB_ACT = 0;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	///////////////////////////////////////////////////
	//read bias from array
	///////////////////////////////////////////////////
	#100
	  BIAS_SEL = 1;
	WA = 10'b1110000000;
	CMD = pd_act_cmd;
	READ = 1;
	WRITE = 0;
	load_sc();
	SI_R = 0;
	runcommand(10);
	
	#100
	  CMD = bias_clk0_cmd;
	load_sc();
	runcommand(10);

	#100
	  WA = 10'b1111000000;
	CMD = pd_act_cmd;
	READ = 1;
	WRITE = 0;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = bias_clk1_cmd;
	load_sc();
	runcommand(10);

	#100
	  WA = 10'b1111100000;
	CMD = pd_act_cmd;
	READ = 1;
	WRITE = 0;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = bias_clk2_cmd;
	load_sc();
	runcommand(10);

	#100
	  WA = 10'b1111100000;
	CMD = pd_act_cmd;
	READ = 1;
	WRITE = 0;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = bias_clk3_cmd;
	load_sc();
	runcommand(10);

	///////////////////////////////////////////////////
	//accumulate bias
	///////////////////////////////////////////////////
	#100
	  CMD = latch_acc_cmd;	
	load_sc();
	runcommand(10);

	///////////////////////////////////////////////////
	//write AF output back to layer buffer
	///////////////////////////////////////////////////
	#100
	  CMD = loadtm_cmd;
	MACBUS_EN = 1;
        LB_INP_SEL = 0;
	load_sc();
	runcommand(10);
	$display("MAC BUS ENABLED");

	#100
	  LB_ACT = 1;
	CMD = loadtm_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  WA = 10'b1000000001;
	READ = 0;
	WRITE = 1;
	CMD = lbwrite_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = loadtm_cmd;
        TM_MACSEL = 2'b01;
	load_sc();
	runcommand(10);
	
	#100
	  WA = 10'b1000000011;
	READ = 0;
	WRITE = 1;
	CMD = lbwrite_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = loadtm_cmd;
        TM_MACSEL = 2'b10;
	load_sc();
	runcommand(10);
	
	#100
	  WA = 10'b1000000111;
	READ = 0;
	WRITE = 1;
	CMD = lbwrite_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = loadtm_cmd;
        TM_MACSEL = 2'b11;
	load_sc();
	runcommand(10);
	
	#100
	  WA = 10'b1000001111;
	READ = 0;
	WRITE = 1;
	CMD = lbwrite_cmd;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  CMD = loadtm_cmd;
        MACBUS_EN = 0;
	load_sc();
	runcommand(10);
	$display("MAC BUS DISABLED");

	#100
	  CMD = reset_acc_cmd;	
	load_sc();	  
	runcommand(10);

	///////////////////////////////////////////////////
	//move data inside layer buffer
	///////////////////////////////////////////////////
	#100
	  CMD = loadtm_cmd;
        LB_BUFSEL = 1;
	load_sc();
	runcommand(10);

	#100
	  WA = 10'b1000000001;
        CMD = lbread_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);

	#100
	  WA = 10'b0000000001;
        CMD = lbwrite_cmd;
	READ = 0;
	WRITE = 1;
	load_sc();
	SI_R = 0;
	runcommand(10);
	
	#10000
	  $finish;
     end
   
   //////////////////////////////////////////////////   
   // Instance Include
   //////////////////////////////////////////////////      
   //TR_MAIN_00_TR_schematic ICHIP( ACLK_P, BCLK_P, CCLK_P, CSn_P, SI_P,
   //     SO_P, VCC, VDD, VSS );
   TR_MAIN_00_TR_schematic ICHIP(    ACLK_P, BCLK_P, CCLK_P, CSn_P, DIGMON_P, LB_ACLK_P, 
				     LB_BCLK_P, MODE_SEL_P, SI_P, SO_P, VCC, VDD, VSS);
   
   
   //////////////////////////////////////////////////   
   // Dump Data
   //////////////////////////////////////////////////       
   initial
     begin
  	$dumpfile("RAWOUT/testbench.vcd");
  	$dumpvars(0);
  	$dumpon;
  	$dumpall;	
     end
   
   //////////////////////////////////////////////////
   //TASK runcommand
   //Loads Scan Chain
   //////////////////////////////////////////////////   
   task runcommand;
      input [255:0] command_time;
      
      begin

	 if( CMD == 8'b11110000) COMMAND = "POR";
	 if( CMD == 8'b01100000) COMMAND = "RESET_MULT";
	 if( CMD == 8'b10100000) COMMAND = "LATCH_ACC";
	 if( CMD == 8'b00100000) COMMAND = "RESET_ACC";
	 if( CMD == 8'b11000000) COMMAND = "LOAD_TM";
	 if( CMD == 8'b10000000) COMMAND = "READ";
	 if( CMD == 8'b00000000) COMMAND = "NOOP";
	 if( CMD == 8'b11100000) COMMAND = "LB_READ";
	 if( CMD == 8'b00010000) COMMAND = "LB_WRITE";
	 if( CMD == 8'b01000000) COMMAND = "PD_ACT";
	 if( CMD == 8'b01010000) COMMAND = "LATCH_MULT";
	 if( CMD == 8'b11010000) COMMAND = "BIAS_CLK0";
	 if( CMD == 8'b00110000) COMMAND = "BIAS_CLK1";
	 if( CMD == 8'b10110000) COMMAND = "BIAS_CLK2";
	 if( CMD == 8'b01110000) COMMAND = "BIAS_CLK3";
	 
	 CCLK_R = 1;
	 #(command_time)
	 CCLK_R = 0;

	 if (COMMAND == "PD_ACT") 
	   begin
	      if (WRITE == 1) $display("ARRAY WRITE DONE!");
	      if (READ == 1) $display("ARRAY READ DONE!");
	   end
	 else
	   begin
	      $display("%s DONE!", COMMAND);
	   end
	 
      end
   endtask; // runcommand
   //////////////////////////////////////////////////      

   

   //////////////////////////////////////////////////
   //TASK load_sc
   //Loads Scan Chain
   //////////////////////////////////////////////////   
   task load_sc;

      begin
	 #1
	   scanbits(TM,64);
	 scanbits(DIGMON, 5);
	 scanbits(NC, 3);
	 scanbits(CMD,8);
	 scanbits(BIAS_SEL,1);
	 scanbits(WRITE,1);
	 scanbits(READ,1);
	 scanbits(WA,10);
	 scanbits(BA,6);
	 scanbits(SAAD,4);
	 scanbits(LB_IN,8);
	 scanbits(WHDATA,4);
      end
   endtask; // load_sc
   //////////////////////////////////////////////////      


   
   //////////////////////////////////////////////////
   //TASK scanbits
   //Scans bits into SI and pulses ACLK / BCLK
   //////////////////////////////////////////////////   
   
   task scanbits;

      input [1023:0] sc_addr, numbits;

      begin

	 for(i=0; i< numbits; i = i+1) begin
	    
	    SI_R = sc_addr[i];
	    #10
	      ACLK_R = 1;
	    #10
	      ACLK_R = 0;
	    #10
	      BCLK_R = 1;
	    #10
	      BCLK_R = 0;
	    //#10
	      //BCLK_R = 0;
	 end
	 
      end
   endtask
   //////////////////////////////////////////////////   

   
   //////////////////////////////////////////////////
   //TASK writepattern0
   //////////////////////////////////////////////////   
   
   task writepattern;
      input [31:0] data;
      reg [1:0]    d1;
      reg [1:0]    d2;
      
      begin
	 for(k=0; k<16; k=k+1) begin
	    
	    if(data[k]==1)
	      d1 = 2'b10;
	    else
	      d1 = 2'b01;
	    
	    if(data[k+16]==1)
	      d2 = 2'b10;
	    else
	      d2 = 2'b01;

	    WHDATA = {d2, d1};
	    CMD = write_cmd;
	    load_sc();
	    SI_R=0;
	    runcommand(20000);

	    SAAD = SAAD +1;
	    
	 end	   
      end     
   endtask
   //////////////////////////////////////////////////

   
   
   //////////////////////////////////////////////////
   //TASK scan out 1 bit from LB
   //////////////////////////////////////////////////   
   task baClock;
      input [255:0] n;
      
      begin

	 for(j = 0; j < n; j = j+1) begin
	    #5
		 LB_BCLK_R = 1;
	    #5
	      LB_BCLK_R = 0;
	    
	    #10
	      CMD = latch_mul_cmd;	
	    load_sc();
	    runcommand(10);
	    
	    #5
	      LB_ACLK_R = 1;
	    #5
	      LB_ACLK_R = 0;
	 end
      end
   endtask // baClock

   //////////////////////////////////////////////////
   //TASK scan in 1 bit into AF
   //////////////////////////////////////////////////   
   task scanAF;
      input [8191:0] d;
      
      begin

	 for(i=0; i<8192; i=i+1) begin
	    $display("%dth AF bit scanned in.", i);
	    
	    #10
	      SI_R = d[8191-i];
	    ACLK_R = 1;

	    #10
	      ACLK_R = 0;

	    #10
	      BCLK_R = 1;

	    #10
	      BCLK_R = 0;
	 end // for (i=0; i<$bits(d); i++)
      end
   endtask //scanAF
   
endmodule 
